// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 08:12:19 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IWpfyuRTcyThCZXloRdPOZAk4P8IRdDci2RrqnawiaMHyZOh8Ol1uspkk3P6l0Tt
84jOUW7Ytk987M+ce6+1ZtVDrZMvLEDkp3YJcnpn4TcCJby8fVfyADzT3yrTeXhL
byZa8uCTm1/spDqwGk3X3ivJRpEyEM908QhnXaPkjsU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1310704)
78tTb1iDzn4fUDtIooyuUa2f1mDJDDl8uFFU6BK5EBe3eof+oijbl7hWwsLkDj4c
Ix6Pe5P5/kG8XNUrVkbC/22UXDuTgkb9BUDmu2Em8YhT81WLD9f2X/6GMK8onenw
gArIrnubzlQfCuC07pcbyaEansgJ78ZrawoHVpPReELubyhlJKheoQOSurGCjCQT
lW0dFkOC8xoudHcATskCLhLOJQR28SZlkWvzNzdB55koaooW9fOP/J1zsjzT354W
AGAUcDdM6vk3x7oLn+o7CUO5BTwyvNnHzMANT2bVqNSyy7Wuv3S+l4thaGdqPYFl
rxo7o0BSuss+1i+Rx6yOpDLshYex1cX75TlVVZm3TT1Zg59dZHZMVbYl05QvBzyd
nVrYCp2z8PbMzCVVP1i8Y2ZHPXL9Anv3x6wRm3a3yoJsXI+WXwWtmTEV9rf+WSNa
sR+JCoioTRQLTlOlV6gZzYB0MYuN4sNKfMxxI42a4hzpCepyEZDR21L0amcdgsBA
qOcADJhB4+khsKbiilsnYqh/ZtE5CjvOgpqAys7w9/NE4DZJJny3zGgUAcDaV84Q
g2Xq6RK8fNXixbHVVUqSbeYok5N7sMnqSG/TJYCnmcuLcOZ7h/rUnaes7LpvGJC2
5dEqVzfpieKi4kup25RbukEkvvEBNiP0wH0n8vGQMaBGoUDQ1jYfkg7JmRWXqIE0
v2R42arEUiaM108taroDdR97qvAAl7M4Tb3NMcjCMlIc4bUggw72xOxten7Sh7t/
cVLcLB+FkEAK/7ekSZ1f05qaz0eZt8drMHTdESJyB20KeDFJvzHZ+KY3epZjLBad
Ff3PY+NwATKgH8La0R3DA/jDMYMhCYlwjeR2V3CvhvqvlsmP8/ABAl7uJXTu7Qdy
tuvE/LrtKTCvPIJw/pwVUlS9aNgQ+dZI9lVQAJGanV0Pgp2CsAEXZnxsIXKFbaKZ
1O9ng3jUfELu9TL30gVcrX2hHgrJOdifwJ6ecaJ9fVLSCOFZrLk/hNGZSBIvEWrp
U05rli92J9Abx+K4e2dtsHT76zj6j+n2DUd2ScuS9frsMs29Vf5uzZ24u1I5BKgz
Yw/ZnnyJoPvSbm7mmp8bgp08pOSZ66dpruK85+ZTD+wlvlnVY82mENRe5l+LMqJ8
34eGIWo4ImOYdV+5CImstLbnNgAZD4UFb7j+c39C5a20BPBwOhR3BQYR/cGKsGLD
2vg7pcElHQ9c7zhTOpKgj0FyaI0WVP9U0R+4+e3Ul4ZbIeqk5bNKwf8Arv6EQlM+
NEeAqi/kAwFKEbXIyt4uNPWD6erQhRzoR8LgOFtQUzsAtuX8Hrl0WVDW5QIWDx7d
pp2IHoFmKolXwP0ykHNkoZD4b9jikHT5zlM8lC6XIcC67zVJl2mA++kS6XkO8nMk
8mwBHsx4GkiZN56ZfrADMcYYo+X5iskZOcvy6GPg0M+Q0jtmCNNw5gRDI5W8aHkp
1SXSFhAu8HkYopfgGzSq9oiRPAdRQLA6U2CukhV5WfS64aI8b7np+T9ylzABGKOK
AAzw0WvhMyF7p6YCPqM00xxT2oQKNYXajebdw7LDVA6XiNAQ0iz0HvXjsuRPEP+g
ZHsQF7DwDqSEVEEVeGiiswZ7kWDdqgMc6JDckA8Kqiu+9Oz7M/+nQfHOPG+WlVyC
BxFCSZPJsegvxkgnG4jKM+Ffkvx2gJlHWZN/AJZPavlCmjZnV3RUFfHbwqhAJW4e
vKqbxbWDEm+7o4lGKL8nFkRX428MXmvIZ4fWuMCKmivXqYxTZ1g+BIXW/oP6An+a
Vno51B5vzQhUR7GsxifE7Nri2+mAcVTDv7bTuuyk9wxMqj6RoFflnLG6ySDgUJdG
gtRKBXZaqpIhDXRyqHkaXwEWQfHE01XMC0RYjQOB0meU8Zn4GFjc0hcb+cefNce1
mQBiY7bpMyFBLVfmlpa/HYEi5adrmVIuRU8cB4GHiIvNrXqE8UNs9/c32nQs5ftQ
PTKUzMb/O5N6XfI+k8iuLQr6P2Jrilj6zWEbLQ2isYwyrTHrPo9BlHO18yBqxGkj
y7sVKrAfhFGr8lA0HXi5Rm+UV9AiqXwBZwLRDVYh3g93zkvosOF651aV8rrPmVvq
WhY4M+JcG5pHHwg8zCEdadAJikYWsm7sHElx33ipmcypjO581xaxm0uGJkeHwngw
fFaf0CzTG0ldX5uec/GljM3Zl2kZEsf6ZDDjOvJkvoPizBz9zp0EK0Gv/HClvuUa
RjtQKEd8C7pCbwADmUzE5J59fnH90p04+gaF+zUHbof/D/0CSZKjM1vk5GHr0VYy
6luqW95kjFiu4IaDULEHVVTH89VZtWEsSUdRbRsdSfxBHnjeV3IIF8cSOf8KC/zW
yVUvYkokUY151ZWNovw8DfrvkmWHunfuNzNMHe+oOIhwQsV7U84y/cza3G7zqqyw
7QFRYycu8dO9cUkWDPfrzs+1HnhUUECn5vDx9Vgd849/dtTbQ75t1gdVYkr2tkG6
x9dfstckNhRWMGr7gPZLob35IejohIJFXb6aZi48ThZskPbuoInr+A9z8CJA7MIP
jKbIG84YfuGQhfy4KMvOutKjeHNXG2KUIUDe4yaiApH+8j32V9w2kdfN2G+haJ3A
o7KlPp3BwhQjN75cE9UhQQbMAjc2lbNWgdgnal6lT2wAtNrT78P8RluM8hEeRzmN
+qqbBxWiasAIolj8gnVCwK0Gpt0yjTi73jNHZKL9v6oX4B2axAgf0bm7grrHcbk0
tAdjlE5gtHDrE/dGfJxhK7psqE4ci0u+E5grojc4+EF0SBcvUkSO+HLDSsQ0Z4RS
HLPJ3pAH2g10D+/aIz3GWFwtRgQ5EQ6uk9FrUNMiehczsCNGcTqds/0PLRJVopEL
fe5fsZ+7IrKWuT9Mw4C4z3QAWQ7/2WjFXbB+mtOW8WLhdKUUgzQj3BTRp1P1D7C1
q6UjodZnYy0ukOF0irk6DCdrcoK1evSm7Hj0JQrhPqjIel/JpxdHA5NwWnVu6ng1
fE8bt5DUBI2ARSnX+iJMXPB4RD5N5XzmKYF0xnm0iKco31riLFmDTpXQbMwICitB
+Ojf0GkcB23OFOc3S7eG3brTuH++WvmC1xuBOcBf6FZV96WGrQt0EYNoF9ToR1of
T/pNbCL8BMML9f4LrQwmFDBpEpJTCbRk/uS2rPdO6cYStGAXBW2nzyHrUsX+qyBx
1AQoDUGEJ6aVAkNyqX4ORfOvCZyiusgvov8DOhiLbOGDek/N3sIM2/J+4KJz7Bdy
D6Gh9K35188wOarzVyKbzkgQiie5l3yGeLQsOFgEwxR79cZ7L/HzugzR0rOw1r0i
araW1yr1htTvEB13yFK6PwNbzB0EL3Stp4n7DHteBjA4UY+maV8rsbXlrxYTXZiD
aQNZIi3VoDdkaIw5SyNd/dHfR/BNlRNIumgefEcfaoP0O1nVEl5ZzfKtT6qTuVin
0xPlw0fs4j8rZGRbxZoqrovQ6IlksaFJTNL5BAe2LzXGme5docV1MDQurSkdRCwD
9yY6CX4dTjsTYe+HshKtjqmrMP5uOzod3HdmMh44mlC2DCGeaFu+jyzNiOQ3OpyF
+pQScufBANiFUUQGbd1zhQ5qzwm4gsKltJC9qeAD/3pa4JqeCjNukQd92ld+40zA
yeK3+IiA3dOsTHBRh9rUaP9LwvZmYvKDam9Ix4DRdedQXVp4gtO6TEz+k+sqNU04
LXIuvnohdmtPy4HziqB/U7XLqGX6rjlUNlcHd8oGd0osvsDi2FHzbcFQPTNiuEfb
c/6tmvBSUYivf0b0ZJVMZoN7L8BuUD/XJOMxpR6gUX+TnP2U/y6SYJWeICPsfLyZ
Oz/cTp1TcbTw0Ubl968+Xl5oHgFpu/2kNOAwpOM7Xw7xH6sE2vzegE2gAsOluY8f
eTxWm0DnrRBJNXP3QKZB/4dH5t8BHblLXigto10xoHLdmgmsWqTiJk/xu2zn9NX4
6mN7eM1OqZ+5WR/108gCDgkswFdKVWdFfr7VFHk7B9vWR4iA5PgenKcGisS1CXoe
iboIfiVOY5Vx7INo4DlBXzqy28RnRZDY0RakodbA4XgWmDPtx8V5zMm83mVKmiJZ
obE2uQrrZWNXHmVaB7ypANk8EiRpmMSs68lYbdu+DBBlrTcUaTTk8e6DgDiDjHGG
O8I7F8uRGAfjkw9i+PRnfelpOLwkCjFlO4hGHVXfmHA7b6RencxBUGX/9vYldMRL
yMcYde5xx9CsUL4XyZCgm+Hv3OvGZpznVCPhfvtk+Y/BXiHsiwI/OFwZK2yTAc68
oTV3YqbytOlGfkrIWpnEKj3RtOVd8gzk1Eh6Vp2mZ3wYihjSEpvaEEU17cFLhYYT
yU0VOgThi4Q6aHtdQnkR39unxYCBOFE/A+8UaNnmg+/EGALRyZ0Nwvfn3IYxU5OP
xZU6sl+BeHk9iEgzbjdf8edCPR/773xZtdCn861U0jlCcVkngHnuAhvq5JuiRyCg
4xj7j6OvefVoAFYFBBRS+mPz+31YdnclQ+5NAKbZwTHZ/EU74SAyJ2a7KrPwiBgh
589vhVEk46szC/W4E7vsl9liULLBwMYE4sb6mbSScsKwsRxmHCH5FalMIzUhuZ+y
zqLlyajboDnup8NdLQqqjyJJAIkr9I0vvnUPN9Qb1hcvIZG0SzCU6wbBCNcos2hu
r6tIjJNtaJjplQ59Fr9EoVUji6lFdASG8StY6cepPo9ol0f2qYajOix1NgtMtabz
lk7j9ft+ssPi3LIsLpqesQOX7UoqfH9j7GEfSkqAyQNWNTMQ2hK+580txmkyV39H
zJoJNJKa5HrVz/5kInT20JUXSDx5E+0fb/sDbxADeCA8cUN6EqQyzeSRJKR1N9n5
N5Hkn/eUKQdQP/3Hl2gqTCpz5JJAbtA3ceRkiy/GS2pn6I/S4/w69QOTka93V71D
u5aWyJz76jeWl9Bpgj1YgBJAwQovcLZ9tJp5W2W6LWYv2vk/b3UosQsa8IJ7vuxh
Rdv6X8tHAy8BL00LdcFOwRmM16BiWrXo7w6lcMLleoyca7TJD4NQmpM+OxKH4Sy8
FZMzHrDogm5R4KbGjN8areqqhKrpF8GtYHj38QO7MOfXoVi1AJgLLK4XBuiiVL1H
oh2/1pkq0Xu6aVO3NjIlNxsXTSgNZms11nc2xt8THGGUk0mHG/8V79eDHnMoDExD
Ni4iK3a0EYXuLkmTIY8ZQztc9+ET2IPGeC+YfEwfMirjKodXAR5CLGpNwX7Zixut
k5YjFJiZ0kfHHDzYdLSyioeFipUPgIPWp/M0rgEl3Cdz2YSWVIs9UY5u7G60vRY2
HnWpQ6JsPrh37q3VQCD2heLdJk8z2jgG5H21nEi9PAbiib++pj4XXZ0geXEX2P6X
mg/YfcUJvg2v2Kj2GLV/Ff/jcsaYviyGFyuWb8SjDDjFblFVS5yr7h7Kcnd4vMmt
fZaEsvcHqPG5PLZvdNJyi1ZmdmWrPQvuxaCs4xT4LxzYn+golPAl+KJY86UZhKeD
kBflCVNgpuBneP6fNy3eauGlJxJvFrSOrtufgtGHrVZo5DQfTfBEAktZ3SBNKg/W
HBrnyKdh5R2ov4JR0M3Iz+LlAk+3zFHLIirOWIneogjmP7HNxLWKJED1CH7E30xz
kXqjqPmCmlUH8NfH9OiCanPEQuHXSKv/J5EePep6lv4wbXBdCiqap4WKYiMgFWtj
fdvBlw03ORkUDEPn3/yXJbwuT0GWsOFaK9yRzNvfNGjQrTc58N7gxkSI5cvTbhXr
XrX80P5TqwGcXyxORTrfHSak028bvJfJmjEK2ScmuTpDThxPMdWF6nnVnuI3AHqM
1XUTihDPJew+LkI05hqox1bR1pbhPLn1pMO8ha9p16iXinT0n7Kn9POLEjlYXSbs
U3Yt4xrD8HM1gmKkbHXIzwwSSyUqxLEXEWnqSkj1GVJXCMLG/bwjIdI1Dm3j0mR0
Fg1LxI3SeKXQMGv+sUCQNntBMzO0hHjGIOyE5lNKhx3CHug553Fhydz9TX7jCpon
mAd3mEilSe8E7yj24bf8ylDptEkDA3AZNc6z3cLwZRB0BxkeHQfNjzgM+pWIl7SY
mLNudtPPNvU+fP2cRAaYign1IbB2sdvdHzSi+7XKDn/1TqAdyHTBDZwcSYO099LH
aTpRZ9e7INFA9i8qhKPPIWyd5ZsJfxMCMBdzk0Gg7vJ5clnJ0lspnsJuj72kPpJ2
YwIIbVNAhKR2Y7jcaMaoaFIuqbRLPT1gI57MmAamxWA9h1pVxBEgaKgtgw/k18Ra
TP3Eey9tdCII1+3EmBDA/7i6Moa9K46c/nzmRgI0XGoFVnFYDBOyp9/AdeHooU1o
lx2BuvUnP27+uo0glrjcMRh+twEYl+6YRT2MfjxRveWCPfu8ZEK4LMhy7m8VPV21
b66Dh1dvDrtpXGgFPD65/TCNoOb3YtRb6HfJZWF22TATsVs32uP563OnmXnWLzhO
E6ML4bAF0SYdNdXou0dYhCM3y6zjBi7lOkEJiGf5RM7WR8gFGhQJj6+OaV83huvu
TQK5uzGiWV5IXogoIVUNTv8F4b3mVxnn+cjTzhvfMN+VWp2ygyGLmCLJF5OdBQ7w
dSNomWcY9CsZ0SsSuEbSKHp6NWj2M3Mhl7m2xV7v2S2ua1zzhRhkucfuytXZAF6N
HotGI2o7uvXRWJjOG21brOdt20T4hFsgU8ulems8UPlr0RvRTgkqxjRZoGzQWRhE
Q2exw65Qdw9bE12YtDJLBqsVkdgQY+zx67d+rygAwnexZab/V61W33BnWxdnly4L
C+a+JlnYE5xb4Nd+0lGwkX0QDaqYcgKYX+a/HCaSj6SB0QgmKBszGjzQ38c7SkUk
QWLr6/6vLg8S/FByB4we5D+Dgc5U1MujXSbm/YKQC8bNs7vlLTdszL15x7aNPEbb
ZewgxaQ6Ldww5kj0iAj+MxlOF4kQqvJf3dd+CizZh1za/2BNsndav4c85SBtB3iW
mHMoEaijf70hTZp5W0wrtRiIzd8vu7MtQtpM+os88Snd7PYtHEj6GEnSz630rKnA
GJYdpIVnRNn2AG0DFcf05F5/k0RARJq8Oq6ZSlxjWERT6ybCQzmQVn81TWHzVq28
2T0dO7VmVnXAnsTRRkHnUprrYe73RueCwmDQVKv4gQdc0laYFjObnhfgqwhXypN2
vQQUrm/5WTeQwO8GkRmqbOLVO1ebIWgu1zgGjN0zorK77j55cf9rls4iGM+l9cJi
TcZBGY9319HkE7gM7i2XQ8avLppr/DlVJnngI0Bf3nUYgywMXV8mXgIGKF2X9f21
nQAiaNdHK8X2krFE7e2enxTEp8da1PpDHb/tmzEM0zy7YSLtUEE7fcWSMdQmNGQV
r51mhqX0w3ZvAHEhmEZc/e0EWalAu+iMg0wN/MTmrQ/jvXRXwziRbjOCLnrHWCET
X7qBLN9iIfzxJUf7pmvQQoYLGV93W58Cx+Q2d7OD0lvUghZ/rpmcE89mEHM+5eKi
1nPlvAE7oh9qz5Es7iXFLq8vHRZe9rUvrAFHv7qekyWrWC0xOeS1crgbgdjMRD1P
zAZqIXVIDWqX9PB//2z9sS+IAJZT33UbH/QsJjSpRoZ+sqzg4Zqyo4B6h6+A8dnm
nN4CoL3egEEO4F4I9IOL/UeAr4VSQyg7eGZIkX6TWPbDy/ebyx7ZyvSs7U1m2X4b
ZbBv/WZOKQZFVhqo89hagXtC2groli8ELJNOB9svfKcvWrClwt+XXAPbYnMkt997
z9segehP4NrMJUxCHSyJ+1sZkoigyDTqN0usuBQPaeNWGoTBYYtTq7ekYQoLwT2X
Y5s7gVNVwMnaPmZuWdunXeQUyRsP+QRBqEYP2tQjqMMiXh98KBkZlGo72E9USgQx
7wj2e6FbW6aLlc0nEBlIwzKfXhu9QiEeigm5wGaoNgiZjVRMYjMvOSKtvuFfWHm+
xmrUsDR44NuoV0aMTjluFy2YwW0fJDrDG/qmRU5KUpgErHWFAWAjBz1RrVKKtvhN
xfDR98gPucJIUqOADrG2O4p6yyf0TqRM/tu1WT1WewhlVApTsmgHdRsVwQV0zB0f
4QOwgm12287Uk1kkayoNYxzCOnGK30R4JvMzTTXR3/oNepScWpOckKWMfm1ut1Xo
eFtF9ITT/Bub7inv+gppXxBij8vO/pyuSR//hodh0/mkrROXTcQolySgwFMaS/ka
OQvHdaxln2+j4vD2mahhIqnFzkTfVLEPh74TmlVb030+hoqkh7YSBvkVjxhSfq0i
0k8PNw1CAhOnJWXrF1yXsZfhArxauas5KDXdzxOxRZJInG54wA1zY2Tnqsosolki
QqkbL2IamRrlx3ci6VFFIWCGVz6E6AyzKvNSMx5YbaYvO4CsKTI5kM+UL1SfEy4C
nAKC8aJA3zw3hOCGT8j+aQMPCgVQ2NK4yfN77Wh+inUa9Hmg/w4uEfHwTl65NQ2S
RKaqgsi0zQFBnWnQ5dgUjbthSOev/FvY8a1muwuHuhhMXwa4DBXjk9mQZWyWizd4
qKrvyy27RavhvdYblGDrRH/kNy6p/JjMyQVatC+g1kxRph2VgujlFOZiIgkxNz9l
+PyUOTvZiZUQUo7c6FsgRjpuBwTXLH0JvD5TMZbUm8pMZnb6wvmjKtx0v018rP8C
7he3HRuvzVx5ORdYsj5VNQ157+q45Mm950CILbtHCPqOoyepm3jlmgupR6EYCPuN
8YPcd6PYuHewYd2j5nYTIBJlcIjyU1MzJWB3Mi4ZfW+7TDb6eVZV0m1qDEtNFaHq
1ATzndimRr6/A2689rGhf07gptqTbNKDgdBQoXxxR/gNOB5cKSL/ZAUKKMno8R7A
OudvxeVZ6TRNCy2kKF6Zm/bWRtT2ZfMgEuN20jYT6gBAS2TWdIZ3XRV3s1kKMrRq
e7rA2e1CvEpThN80xGKqyc/NQs1CY/44Z65StAuG1DkhQ+tmvkSOnzK1qsunxwCM
FXBCZvGHRrnCMswuzOUGr6+DuKz3VcoLOS+EIy6Q2mZb81f/B/5rRod7Rf9Ao9ad
f7Zzi6cYD7f/Iks7KwaYKaCdfjeOgvcuUcb3jxdqt4p9y7L6pDL0oViBvv5SxIem
J2lb+9YxoknLVitCHaME7G0oDyH2U7JCVvfe+OnvkDozSsF1OR4N4LRQ99Xv3mgK
3kUWgyNapV5ReFcImckBGJxQBng3/RDFGVwDhqtM/w1MDo0Zyk2Ami0m2QiWUOcI
fKfBheHrP3rqAMEowWz9XW8vuptqg5etP3PlOZ3BGeTSO7BNw//LLrvFCxEt71+B
xkvuSpetD5vUnHTM2be5jdjsOMpobLjBh+XOHi4/mPbUEkZp43JjXMMSuH/YuhEB
QJGv4iq8t5miuZjD+W9B2IistWL8gIq7XZ3fCPRZ40CtQQ2WStDk9Lf/iehlOSqU
AkxHSA4Z2Bb+MgCEsOkZNjKifX7IfA91a4MCRbgNDb7owW8QTVrFche+jkOWv9t4
sLrBH723w9NoMqVmnolJRlhPJbgkYarbPrHJdIHWYnTAaT3bEKbfHoHmArS++Jgy
nfi5qcvoNJZBBEmv7smOIpUG8SuB2T8xL6MWH8Nh4UEHSo8I0pa+hwq/k/ONbdvu
FYmPdFD0RmVCJO0eXdcWfQNYxu2IWF43dl3oOP+U7Eq2tYAqT2KLVAoGSYnEmcA+
dIyTWHijhtFVLqCa3BW/k8PA2pv9xzg9AN+pObhkilgF62R9/+pcdpmtUNGU+fnX
O52jUCRAIa8LX/LGsCbcYD14dI6BYICsgLq2k2aXduRUMXbLL5dEDrQvkMIRMgYW
rhtb1BEXwitRgAPyP8Cj2DBugat8Cgk/KBg7fWgbBox5ZMcCrPiDQR/HKP6gKAqQ
Ij9K+dGRMrjf4B5oCrOlhpBuW2+AkrXNcfPgzRIT9ywtuGXMyP2VZMvEkZU9RDd2
6hEyJnUk9MaWIciSW445+UT31QpTqQ3RPf1n55MkJwHjpWXnvAFlh4NGHqEhxIzt
Uu8Yc3W0JSy9ctTSSHm4YNGPEcz6jdoAP6WtvR2AnKrgsc0RJPXgIeBRtj9mIu4Y
S7DFwnw5bcLAI+BgUYcjm7tCZFpdfrPns5eXSbpyEK3P5EMDr2fW0S5a+aMrFh4W
ck20M7sOr6O5fSQR9t/Mgwe5UpOCrTQLqZQvJOd6I/xdIy4IcOh0D8kZxAZefE41
4ipr9KB4alqTrpYV8goPTXqIxP/Cs3i4FyimF3gwpdTwobaAYkJDyoiOr7rQjdSS
KOnQvsghlx7+M2rjSqP0g16Dnd8nVPCd9B05Q/3obVWwgXeNTcCZ4MqntY5wDn41
Yuz1BZep/5opnW3DZg2Q5QcDh5wHttuPgI7AgKHadrLJH4XMJdJgys2iW4KQMiko
IRGBYvxVmkM1mKp0yZluApWnvMChg/JK/u2TE+oLXfyLWbb9bp43r/Fs1QTFUszA
ZuUcXuKG+X647ugwcAcTPT4iOEkq/fNcG/pdqyyg9TdTmqz1JhX0CgHace5ioVY1
NU5zziuPD7THfkqswDqvCGpok9WCUfO3KOhmmfXb6lLIT34MVoE7HEgAyImBBdvy
8xcD7oYcQWP90X9eygByyVL/KZUT2EtEYPpiKIn1J/+QSCi/aEz+h7jxgrrVuz7O
DyYmh7N8pKR9URkTpaDnUiLnNH5Xw7sAt1QLAmcVL4GoAsoyNrmsOwuY/9vt63V4
WMi24zY5C64Mo9omaCGfsnDWWJSHx5fbkjQIiAkmmyW3/ibMBEhcAoqdo7N/rNHE
I66Fp8VWg6su/UfVrIybN7df00hGPUsGplhx+08lSuCaNGOoTe695fTZN3rMSI3W
x0eOVzfj661ba41Wf86sz8K/k5NoIwc0sY+Vx0WGL4phcH5UvkCc7SnF6dUYmS6+
0FV22MeVfv5dbjmeJ30XLRIQLX7sQ1l/uTUfki/Jb/TukXeT2i28l+59tvMqiHbY
k93BKA/L8Jf0CKtvRnKal+7lzvFXW+YlS1O/tQcucKstsO1lvZhLMmlewYSAVzMV
c68Rw2EIrvUYdsfCmZhFy/fBZhh8LpQWvrTlcqNIqaze9YslevdMwZR4LG7H3iKp
OeBNFHBPhec/lTFJCKqN6z5bIZDzCC/1Aqa2wGTPupMN+grBU+AvyJ+sdBr8CI/I
z9kUgqUibHfaN0ubFOKd4UoGt5gQoozsmB/f6Gs6eruEpdwJx68WXwTWeZswTRoB
mIrnEvl+lc/VxTCUGJaE8tG9VJXnuIC3CnrHvnxh2sHM302j6HCfJOh1psAKDS8a
sB90Ilqc/C2JAtkzjiA7UmwAvzf8IkgGMYU857gDkb7A6mFBbtA/c5F6N0axvvda
5t04U5LlU+8ODTOn87bJaZXd8zXQUm5HQPfzljQewWWMIjiyAXwVIt3JeECvbJJ6
MQ1v8+T+qbRbZkqCePSCaAZfDqgqF6ssuGmbC+0f/LIvFOxmq7eKPtYyj6hshC9O
8LM3SFaQbKEJPkJg1xLcSctS/21ccrRJ4DzGwbSXlYMYkq0V6oeSxA4w9yROWl7m
2vzKirp09nJAOfu0MyW1UwcY2mGrCqGODXlJf72PaPZcyPBWhQ/5j+aH2Za2W2tG
7oQi4WivQ9OEhI5GwAC1lDQv3G/4u2L4C9cy5X0Hd2ZCuC22C+eqGtszQIz9v2RQ
owZsckiHAM7JVF/KTsH/6ngaJCvvG4nGyuJL2TevqjdTG/tI8NQG3hGss1EtdSYu
7ITbpqQN9mdT9XrHOGrj0tiPecOnQNN2MyMHUmFGwX6wOKZJWA+/tfMC80sIVHcd
NdfHgaY1oINxa7p6gqlpz8ZrYE7KculNHxCazXfveTS2+l8dtQZRfUSZO00tsO29
MSIWVb68gSLvDIaYP7LHrxyfKr3y41HPdNAaGjRzNQDlB/1cyBCVFInAS1o7zHnC
O01v/NFpQjPynh6i+xfrrPkeJDnkCm/jNEgcpjZvVwDKqUbjWznAgz/oGBC1/acY
No8Sn+N+pMaeBGNXvQNnnJwyJtxX1x1J9idQGFnfUuBNse163SwLeQpvugghOYzd
bpAPsQPk3XEviZdrZoMMd+jzupBpZ8pRNob4mR4Pbf2qu0ViO2aDtU2hlPuLQ1vv
k/3/WtrbPg/1CygZ75Ww4MYgWcZEeuNSUVh+FXZHlpGS0IgoQHGc9ieDJ4AlwUOr
QxuMCRDOzKUqWFNiMPhEKZTZBPdQ4HrKlmKsLaHdgWGWtEK60CF+Cjwvgq1SkfDB
XFRoXh49x1v4PIrccb14pMMnIlzSVqJMua3CwyL6mwbMLYJ8m6qtjGkrWwW7vknc
fPgFXhJOhYiYP16E+M3OXZxR9Qu4PCYKFTkZcvOZeABuCuwf9BXRkapgK1UstRlh
yBOkV0gM0WPQa36r6hnme24mLm1YFlcw9Q0ePMmJtqFfScMxPQxFOi4vQtTzfw13
Nsk7rMvGY2pVd8QTBh6o24jOrK55fVo0uLtdzNWxeHV3lri49Uqde03uGu3dEkLy
kTxTSfw+JEtCNRDyupjn0R2/zuqVgEjqIapkjjMQEswWvlQVNXTJzFFGrX3utAkc
AbY6IMdpyLHObNr7pwGn3ygCK6Fr0uC+gSTKcsM94Iq7sCrtSXG+yh03VYmivNJa
V712YwfS7O0eyfpPVvm7LdbY+RTF1IMId60S315WgQZiPsaM3P2o7rGmzXBLjRfp
lQ90ExjPZFztiCffh0YN2QaSE6B7/SnKsf7pcvyWANuYPX5HG7IcGEZgZQNNaIkT
cvxMABRA5a/hy5IONS5MFJBNYdMKdVxMGAr2sio89gBOO2bhu7Wco+LFqsT6giWJ
+1q3euRuMo1fqm6HsaTGkIihe+Q0Lru+ZzohIPMiSzcrfiDJWh9IRsD0VCtC46o9
GTLdli0Sn+E6lL+3raakPa9tQQioYcw3tV2uFVXY6w7reN8b+eEfDSBeo/YzQSXT
htnElVZepDwICUFhJfRQ+V3b2uiIY7eI21uvAbGtfERYS5NrRjX295laSa3ZiA8c
5pmXtPvjMseHD0IExmMwt6zdTa/nr5X3TwtIwL8w1tJ62zFgenOC2FvPUY8XKoyD
TOP8trniNR+q1cV0//CAYRqKbElJCjaxfrZ/zZWfBcplgejEg/3/OOFJn/0vxOkw
JDqrsMQ2uJoaWsQQxqIeWtJMCOay9RpIzQqztJrssOzbXlpz8X9dAHJpwiFWMyQ7
R/fL284vV77/ue/5SBflBn8Wm3LsHxPjXMqPdveSvZ/kk2i3KzFs5U8BAqmrvEeQ
Yj9DRlDOteFBpQUeQQU4ovF1PoGwCEu4mv4qDvS749AJxGWskniwWLhqwGR1jJnp
LiCgueNtvPHX3GNeeTo5rtVarHI0f9txQqguJaFctOo+hI2QWrrB99ByAQ0cnmTJ
m2symjjxE3VkMDeBJAcF/TQ0SZiQDW2saTXgyKgB1NJ9JzJSqRv1Or11jLnt+UDC
TQp+MCeldI4U8pwlxCoVmZeKtsg0I5LESGjTYmuaCMxLLYTTgYFSGhu0GB+m1ZLZ
vlGE29rqA40WYo7mX1KJpYYpIO8q16favLs1kjh0c0MKLZzCqYqSEdPR9BkD7Ecl
GVXHS+CJMMfhPOP9NXTpknYIF3GUxjlFbYNgPZJkXoMQbs3THxGuMWxZK7MkwfkQ
fNLW8xrDlXZvx03m9nXHAWAOcDR4RPVQheIfWd3sedqmKQha/5AAgpII/7pJQ549
GeuWYzKuFFkRZt5OvZGGLIDHw4Z8fIe88LM/k4Z3y/Jz0nsR8mOrm/IMMvaMHihp
B+3wMB4eb+GEo+ev4reuimfLlYIVjz/th8YwOPrOWXWWCVkZNR8mlkUYtLIxFwMw
RetJnB6niQioel8pWjNokCGXOffRriyW6VJ+1Z9gI172uqwJMauPvQHZT2OZJ8Gz
1DYuIYaX0gkLGIw+WUB6YhCkGte346DGiqM2ytr2tfQ8FQq90XwnOpE3Nd1B8+5m
vnG8MgP9xTDi2dK6zFc83aTXii5n8dQa5J9BfG+8eAoFGuktyjYrj8/BgiMRxjRU
/t+rjWDOcSHOFZ4T3jaOvakMO1oOhqhmlq/Bm9p3vsxg+dgZ0TGp5Qp125J5NFaF
Srnx6jLfj0xxRM9Gym/WMelcquOgHQmuDl3OBkADdKauxE1IJZEONcvp8bXLrFV/
ceQXEoaeovpjfioCtpDoBlrsIMRisyzWjPAVagMUK8Qqg4mdvniMrTFMp2PrXBQR
bmhShCQzEtw580jMGB8VmIgjVYtbWjYhJBQjke6mMEpLHeKYNo65DWw9uzzfVqI9
pEqQH0MuBK6myxIA08FnbVtBeeoonn6UkXNLbiivbR8JeAxRvN28v99F7Fq7ex/J
8Ud8nabF7d0mO7PDMzIiIhoQxEEUg/z5yoAf9R22cdHgzPdGxSEoJF2EPv7Hb+z/
I+viUE1hYElodrrlBKqQmVowPtHe+3z0Oh58BHqOrwAHa8enErmgCq+ap10iTcR9
up66qA1snWL/E1wiXNoF1xs75kIg/RDH0sfTZ84/GneDvFsRzCdCj93PEYifYAon
v17Dg/9fBsiHqgwGXsuuMomRNMqUpQo4SuchN573h+nUzhx00Fj25QgzpAu9S0Wi
4TEnrV5BlazFcw2E8df9e/9aHpcPPvON2D1xjfUl2CVGkMbAo1IxRZE2/jRfuHwT
+BrFrog61udgfBHGPP8Q2nt8Y/eYjq9yDUoyfsbWjrDFEGlsRNAxydab9IVCPa0A
XLOKsdx/XEQsUza5BDt5bDGVHBqDMBLM24+i/c7IXupPARuBV/fPhvBhr6WIA/ZB
GHpKzUUEb/SC8hnswZ837ek5V2PlhVxVYsVLqeXJGvaWgmqCU6k3JX5JqwORNS5u
gv2HT6GQ40JP1cQrnDPLysWYFYalQm/TuvyJnd49tfFfR0XzLAFFK07+Uht1+CV6
lLfqq0h90vugz3A1piqjZYBQwMfPtJ6P7ctuKuq0HlvLNCBDOdT1XWM+rCpjFACr
4MIOBKa/AmCcH5TxlYA2BpYk+wy6x2zTUXBJCOMVWQ4gIwEwkseXOUPmsE2lUZZ5
WCoOYaZ6hY/8v1qZKovRYH3UAbyqv3btbv+WYvaCEMyn44aD+sHrtVm0aBWvvpy9
J11jHLc383EwSHWQJr1bTMlzqUnzm23GAnX9Uxsm+q1KAa7ARWZgEUY0cPgZoB19
h3KmadvwTzGRRPRKiClgUcyg08txQJwwzI7tesXSQuW2KpweQGlhIFkGSTzFwtnh
ZDQZpyA0gsVdA8SE/vygJx4Giz+S69RXuQTE9MCeFrGJegb1SUrrdE3CMzRRTM51
K2a9hGUz+XppnbSZgu59RPwPm23HuzUVfma2sMSU2n71a9VPskovbqbh2OVbY0Z1
HXc31NKozUMryHUkAI2AQYoimcLCem8R3DuG6WKdrC1Axc23ZJ81Uq4dJfT/Y4fS
RXNP4ZfLOOxL5FCzDHK8wxjkITXFvXEja0UpyINGG1SE3SOavRyTm1eRvF60WkGU
I337rshUm1VG3cfcX270V1HlmPG+o/xtx9gcAr6fM6d1ZvrmMu5FXTb1Kp6tvfnA
+6PsaAX3ks6stzWNhXVQ4W5vciL8I4knbxX60zwhrntSJDkugq68zs0kc45lKtT4
Wd+U4FQ/KllWBCnbEAExUarbg27OU+p4o9YodOJDw1fuWmi2vmpzc+v2k/vqw3ML
1qBlNp+YKqPZUg1MEFjiea4ybqU70B/7l+iKq3sCdRGtRhCNuRw3bv5g0hCiMWhy
UGof2mlx1NAe5Vpu1IEewD7VSvCHuLOxwukPDz0fM2HkAlHfW6w8pzbR5hUF92H8
hy+0SQV4GYO8gs7kgax5cH/zxi80pOfCBf6IYKqUEN13J0MoWq8yGW6B5891B4Qc
z1d2SdwPLbp7JxSnstqYW87kH5v4f/GECRtM2607AEZ4TIKuQQ4ZV/ssvf8KYR3h
920IUNY1OE2fpCi/AXuHzflrMquXrzgVZ9HHX4uBlFDaO7fAGNXuW7XfNnJT08bA
U3v2F+tothqL6NXoi2StHmLrXJtpDOqaGojBeBnixIgm+83zZHH3MUN559tZgogk
fApzfYhzkPKi3QPzH12FrBGfD936+BcpofKA6tJBie0jIlGpcfy54VzQZIrFFUFx
Xb7K1ILXD1NNqmt/TVSTigOvuVxMuFZ04UTTRTrKfp94h2m5rA/pCmOcam9iJi96
o5W5rYTlluBKma8JXa7U94WCrOR2762cW+3S8aCAdmMxMLTpoq3VGj2kDi4GdkyJ
+he9Xo2GbDNtUiuwA70r34lugmMBP/4GTahUmHSKweM4nutrB6Rb+my4wIrn0fL2
KkPPeNqwU+Pb41hRqy5qAqYCfms+AgQJwAmKrfsa1ZyKHbOT98a6r0NyLnsv7T6D
2talOUk3XmrRpkXDlZFmk3kCoMegfwAph5G/TJnO6rjgkTsC58D+qR2Wjv/4Gsfs
lxsXSnOj21+dBIyu2gvUpc/1AupvA6m6a9rWq3Afqp4fWl0iQKqMbDebsS8mfqAe
7SQ2IlWt8fP/06ZBxQ0fqWD2L7axvt8n/eKwzIWtU6m63ECRsupeNMlEg7y+Vkfh
uSU/eemQYtk0dljJ6u5vkLPqeY1qXNZIoLV5SfWYrKCV499/KhDa8UI1Yqpg3wJM
+Q7VbBr9esCctE2sZnNuvdkIzc53lHkSDA+isrnyj0CmJd3DYdbgMhKrjgXe8Tuz
jM2l5kEJda/ab2vnlB45aOHutH+02vR47EsrWtDPcS8ckeBcHfb197fh25nQ/HLX
ImjmXgZ8hizQNN8EVnTFFA11vImh0lE47iiwvZWSj4wn2ZkLVSfnBmZ071LyU6Ga
YsuGYtQPeEep1wYYkjaN4ozHuiv5JB3uHMXkbMjLvhMiOaTlhqFPzTB6uYEc8CPo
ej8NzFoc6C1g/OawOi7gmRLoauSHx8kbR0bIR9i1D7F9O83ANhOIFdcKUHF+7uTP
TPO7i1dzSPBoufceD3Z0ACBwc5UbOow0vm4uxE+NkaR1PlDv7HAy6R7SRMoU7nJ/
xCOfArRHNmUgXsZVJe0MtZh077u6rluoRZqdvmLz+/9Gm0P1ikm3D8aGUhuaWQGl
8o0AmxUCd00iN51o3k6CHUY1iuHsA6fLCeXjysZFMiMfz1Zm6bTIT4BhMsLJGXlX
xJrCYVYSf55v3+ZVCnH2HyRV3OdcK8xTCWtHuKlCtbgOyKci9z3gYkPcEH3XZdAC
2o+hOOWV6rqhYYsu9s+of7FQlKhxA8tegbtwxmUwPXSSJPITXH9IJKy2B1NMHM7n
jII6ieJT2X4ZNLIF1fnuAVAudADu5AnzxSOmk2rz38N8trraQ3e5XfeFKXyPrciB
yQ2Bqh5JSIqLmRdjPmmeRIkDzyUIKkIxIVHxNCTSaG+Zh2SepqD/d9xLr3WxZw74
363dcfRwb7it9oNzM7uvJNrczdk3hX1BAbP3r/VCn5PQq2Z5TUaEYXRxcv08di9m
LEiVlsM0TTnj9Rf1n+xv1PnLwtmO/4l48i65jAc5Mm8jLUvUwXb5BIcme8bf0Z/E
4e4oDRf3EVP0YKVg1D81tx+HC4ABf5MsTv4/CzK5cUvGoXg9l6Hy6iarn4hsVtgw
I66G92CAXvNFaIA5ukzzSqnuLaQQlHMPsXkIp/5KkuPu6GwGwSOb+WIfmjFqXiqn
QekVZogvw4OQLrWxXLMgTyURXgQQGwJFl1dmqGZvp97RnU56Xw4CvjZ/AHVvejHp
AzSmCRlauvtkETSkSYQ5dafaY/WBc5tWCk6Wr0d3wc/zTMcCZv9tZ+s0pnvmgSwz
bpvU+U0gAp3otaawrLEbPLTQw7Fp+k3VrgPdLRTyOVKZCwEAkEbubKMuLNgws5i5
A8dwVOTK6A4/j9fQeo4SlKYyem4PpHlqucfgqy2ztT/X0BRaRusP/OyNSO8Ii1YN
hMxuQ0Z43YBMrWlo8iyzN5gQsvbwaeJxSGvK/Cpl2k5kzxZ3Uwk2xMWdbJtai98q
2uM7nkxvBjDl/P5W/64fcRDL8UQnapMyrVlsgxA7mLjvXKyfdi+4o7tEHEd2dZ4v
nFYWY8uW1dqj0EEg1H20+oLPlIUbKLLzTIlM58Dfd1iwS78i7U/x/GDw9vcLJFgL
Zb7P8ZjKzIqp8Ig6SXUOBFcvekEYJ8fmUXrFekoaUVlir/qAJtrxPLDwmPYdWNhW
jgCTcdnMXy6pEXIervWEJMKi1fWMvR04sGp+1lvIFjnZCzj5jzaeCac3SGq8ty5Z
xeQOrWTMLJW8MVO3hPSDa68oVITWbV5vY1orxJv3W+7iOCApm/EOwzcQub9BON59
u/YFnHoR4xLJcQc3hj5Q3PZPSVmu0veQMCB2WHYlEI0f+nnqxZU6PefVHQdfdahG
BSAqbhKO7nrBdIpiHaWADm52vFYCTSMod2QVN0KLaTolRgJCDlAkoSbP+b6y2h21
LgMl252wzcH5hS9brqyYPhJgP2wKky5KYPHIrpdXrHiEfWVIVZm3iErGmMlqlVu4
Ym9Qcg9bsavk38oKIjL2DI5qNLAXhlCRebjG2xMXp6jmavP3u6bf3dsxlSqfXBDy
wPu4oZM9/9RiYr9ByRebzhgch1GcMjVO3+ArDnK/w93SW5VEGJE2BKa97Dj+hm/v
dXau5h5gOFOrEJAKZU/hpCO0Fojw4yac9xYZPDBDWlm1b5nB9xrdoaXwz9aN9Vit
eX7q5Enwb2SKCxoQZiPf3O2snZIBCFnsZYMa0sOXGUFOo30iptllRoNXO2b99pm7
a4nociIiSTGXbTP9cC6QBPkyQrsrMxK9q/ve64iMTvcZwzAMkfAf0w7lIepOApVv
pVC6Z7tub+KLwgPrOlnv0ydPZJkSkt9eZoObnlZu33ef6KR3nEWaiychh9J0/FBT
zzxVWxihgT+vOU/QwxUQCNvtnDP2tm+WlC7c/ex53ePZOJhKJNG1LSikPId41/lX
pZZIIiNRLXSjM83Is+/4KX5pTLAdX3p7KghgIrPed5U3zzCW/bzz9PKKC6OaU2vm
mOmEnodzQQ0VUxfpPhRDy6jPlx5PkbXj9EYBB5uyhzMjJzbWdW6ilCWrPe4764ar
8qCa/2exeWqusdHLD1hyMTy/cRO+gXLKGDMRrbmM9tqg1YYcV5F8PTFeoJEsj8HA
NFlD5JeNkKFbFSUccOShsJbVvRE20tZu+py6GgUQFJf+uIK+hHf5cg+ofDC68hA5
rC4WNGYbnb0JODopRcRygL8cosOl3t3WxPBLFJ/IZBGc0JZG2vDFEhjpRVdGI0sJ
0CQ61ikg7wMCToVuVx9XA43E292IoPZBHf5fbQsGQxScfdVzT8ErxvFjfOxd7v+/
iZmad6HD/AdQAx8DSawglYATQXo55vmgA3zIWBQsbQ/KUIQLM9WpQw6VWGB3hRrT
FxJ+c+PlG61K2l33qED0dJkrgRX/YX8D/BvsVa/Thn3wPjNOOaBu34A62RrD2r34
XQHrQYxNxE5s5PZWgmr58licIEN73Celo4UY6Gr1yNhCdmwTc2HVxlUD4KIE9Sj/
ixaQVc0ixbSTJuN+oqHBrNLQi3l6HMN4GFny8y0cMiC4sk3ihl+OyJ8QDV7QyvYR
/CZyer8lzvHQ2Y85n91vc07lXD3oAbH6DKGl3fnVr8AAMyJpiKagqJJY/wesQuXW
+bTBhq7EmS50H9NFwcueOqn1imFHCIa/o97wMZDxyQBatKhEmMw+SaDu3gvSTfCH
/WRXunP4z0X+STM9PrihK6u8BaGtLxobr7z6AjwJJqdTotBm/Vc1qvyvBQxKskub
3hAbe+0N3rnIgvW02V+GcgAu/C6E0l9IgS/4GP4R6XOM92jYGk4ZJf1T7qcjIgqP
ri2aMVyA8aR+tNTo2n1Al2yOmnmUOIUnXXCUErLxLmP/VosVNpqKBJCwGlRVKn9s
bVdJGHCk8K03Jgfz7TPSQKkdRHSj31TCt/bURSlxef52uNmpMOOv9KEgQKHZHliS
d1XaYVunpY3lNs0JljUNdTzpnVTrC279Nj1gSaRc+zVx8G5YmyS1qtP7p4I2OQ3/
28aGXtmAcOPRbVqnhyeHsXAfGGbn4NQkzoKSLhYuKdZaw7h/IaOgODmpxwX1Dopq
ncgmiSYPzH9y36nOV0YNnClZzxUR9jl6S78gMMN+FyJ9H62STKvfjZrspZHsRPXt
D/5GttSUWEp+G+jiobybgctyF8pkG4dvvYG4hEo1NirHr5Xdz5pNsQ9o5ZrhWNNE
Ds2Rg+SxepZD3f3sABepleS/45XC8VCQu6xBmLU6ic1+fz0n232DqEZk3oiFWNNb
AUkeOQI7jIFo0UrOpe1F9MTMj2udOw7K1kt/rLstSAMLhxVepsitna7Ud2GLEbB0
iv2mbpcm+CiVkWv0ixkCN2YAn1T/SBFpn/qVvt8n5yMR5XDFNE0i+cf/QnRI9XHe
u+fqdhWpW8o3vTqfQeTClWzkl8cLLELuA+Nf7eA6iYPcRq2sz+IJ7LzahUV+ojZm
U4YBDnVdBD66E9PUiUm9xtO9hrGv6SDGQYIl2eeAEe6/C3+iZGNFvWyg1WrqgbH+
Ozlh4ItO7yvycK2SeG6XG6fEGkdsMxj/anp7tL3sTofLxb5Nrf5DaiS52LVfShFw
ex0JvKEXx/ylA0SPuT3uUMV5BYGUUf5TLyPrlkMjwD01ufHJRxhXjyQbqioYMgDo
RzEw/QtA4N1bliQ1ICydzEels/ukGStgWT4+SjuQiudlsmovrfZUYFGkGg2pvIxI
atzq9xgOsD9MZ0UOT0O1A2iGuPLjfHuHjrcRogwaKUVg8eKs/6v8GZykVZwcINAt
wHtZnvI6QS3x4Ss82i8bsuhGAGMElMqE1cxhnrt26DZhsdHY6+Lfw2xbhZ9o/7TJ
ATmE8MIwK9wj/eFxX+utIWZHik2YuvV83TCM1+rZMM6fuwk8FosQINDEjOZ1HkDc
LkbjzzFI7QzNhDEk/uHgZn+V9OIavbOcwMDt0Fg5B9Urf1+g1izPSYPK5dcShjKt
DJMe7iSV73zR8L2GXy/untLCUBtlIiUCyWeov1gnKuWmSheGPDGc9jdZgLkwGePn
R+/syKpfuvACNdGypYVG1P3Q2ou7xsSFIp8ZFYDlWlVuy9M8eGRcH7taeYL/D+0j
VA9V66WpU2TUZlAubAcj3FHcu9K5rqITrxtlQEKmrfwUUITaWo8kTsPVn+TGpJJy
DzUpT+vmIa/+JbJYWslkdY4ZTzdwZuqS4IGeW6T6BuIMhfblaauT45ndhDeXAKxP
N0cUONgNeZoz6sY/UbibohzxNHaiMl4zwsJlvoZaLG9H/pYmlZePixnh9aLfwGjD
p5S0fl99sFaL1Me1Esgn2/G34ahM181AYqdjSSa2HQc9pG4lzsgWY1phismndYDO
+WcVVm4tXrAxHExCrHsg3GBLuk2LOvxakFivKTMNVPYGFjsU+LCFWm1rUezzjsR5
Lm/rOaTocTuUfWH4Hd5sqdJW0HyTf/XMS8hn7frH6MofqN4D2kUq/pzceM1/mFLW
TQSPDZAjTIPJK7kzwTSwx5WY5qsGb2YpRW1cDqq4i+QNp2BHaP9zUQ1Bf6l2QiIm
D9+26NIjTIK5nX3kFVGqhzEl2QTv36tpl+6GINUQph6RtdYkb/JBvS7jCW5KmkwC
Me9SGd1hIuvrWEC23z5vlKrS6FvkX3FWTthjVfHiWlQeGt330mDfEbeFoR0v0kAO
wbigmpJV1qOIqT25tpYowPWgZVFt0rSK8vx70SGLKeEqaAtrKcQpZ+HtZvaSA1v4
gbEsB7NCdn53TRmj5RQqFZDwEbq+KCClwq+A501gVyeD6zhhVqStrQtlkyu4ONpa
kFyl0zHeH6LPP0YsxEcr+BJ9JcGxky7OmAtS2fOPKxaI716MrTO46QRYHL/ylt4G
Sb5rWTJXqQf+XwTbI13vZZfRlVoa2tmazDTCxZiqe1IM/+l7ptjtyzrwr5FmY/hD
zOv0B2YTl7iQZLAq86PwM08GVAzCX2r1EoV1oXSiC2W4XJBsZW1/kupvurE882dJ
vXA5FJe1zYM1w+H7/V+XPSYU6ziXR9g9KueSVsEUG7XEZIBtYsfTArUqHoYXyKSo
PzbCQujqC5w/PLUoiO/q3InPwTcQ2B5o0ENw0sSyVGuyYg7THb7OOofwhGt6+yMW
mPR976EoStwljSv2DkiPgUiDo/Astw09UXFbRySveYAVUOHyMRSrjugdIAZG6MIF
3LCWgsMign45sR87vREZEkVUvHbYpgDYUJsK0e8osn93k+0Z9YahbLX4WK9ZFE0O
W8jLNbyzYa9iAp5XSI05I9lKTDKCTTvFku5wIvPsCpNbDQOF219n7ay3MjrBlmWG
avwRZ3boEpXwoI1BRye9FaXCZrsu3EBj6nW4alcveNgYmZsGRdVG1iANX1M71yyL
E2RWfjaPVXxsioS87itskxE+eAjMfjbipQi6iNWlhPwMTdfoKNaC5bZbYMratSJp
wzL0uNE19p6/adCqZFUJw25jZPQYmnCpRixvf+CwzUSmjfiAGVUfOkX8HkKkiC2/
n1uuBeHdfbzXbCjY+j/lv7m5A20QBnXAV2dn9eK7H1alQPVsRhGsZkWuvdyFKRax
3BvpsXTLy1289PQi8WSXo9UmvWDDnOPDmuvBGWKxsJWpZdgC0XI1Df9NCVgTWu8r
y2o7I3KbOQTU3wFKoWLe25DSkD4yRPmc3yVn99dT2WmMMl0H07YV/1Omiqc+3qqj
Z0kZdcvZJIBspoUrCEvqMcwnAzsfP2mFuFcymU/jQMV/pmToXqcCtJeWI7nYyqhe
fUYj5ybCX+JS6Rx8f3LDIgbo5S/186seXqUlF7ld0jnk8WpeBRIg3kD2cquLU8Zq
3wK5SNw/aPgMD5iZwGHPUH6JxgtKR+33tqc+E/YD4wd38umghyide19ned6G07uz
doqHh9xZed8MMQuS+so3J0s65Wuy3HMdLh8i4eXM0tAc45jXV2QyKuUEVZ4gGgT1
Hlf+MfnMrJXrRD2W/i6/jCWB4VZjziCpeo0itprCUBetBFPqnO1hFjB37E6g5ueO
ShMkdSbSQlxHahYNM1f6QXUK/zyNK4w6c29WbiqDtKC82HpeGMcHibgMJbCXDRdY
eWv8CF8e1y7TkIkWSFSzJR8uyMb3VrrafpbudKNPfxCzvnpF8Cb1cVCK98Ofj0Ku
vhWC0hXGiYrmXn+rQqQkTCeGXUbqXH7V95PtVuW4Yg1QmzL4BliN5whVMyxdxP2m
U8yasAW4nh4CrJHj50vcVR9mW6v5OggbM7Bej5tKj/WB+HptStRcPFJQRuo3g+jm
tU3ynMZb7pMOWNVcwjgdziQUVEFrhHDKiZM7Y3S1bIULZK7t47EcHtGjgayznJc+
6BQGv5cyE0/SYrLLbdoEDRhLU57cBam7oLs3DahIAnnYmC9WvLD+Ghd3WG9XqaXx
YrqPlwh1Ef2Uk2mcj3zoVCvjOiBiczsUWL3cMa42mR3tzFcVrUE89mZuzycuJ2oH
7Pl3KSirVk6p2vhdmvKMsPA5YdCtsQL4vrFDU5s9mgpk6DOO8lx0GA1N0nUaQS1G
4lid6db5L8hL82e5uy4AU1BhH2EO5DH9F/YzFmF8ud2IEEOULLcmNm+pP7/FGylw
Ox1Z2U+oEJE4TmnKvwiiomVZw39D86xqksfXFPL77/Pn1c3zfRrj0A4DqZQ1O7/s
/YdwKP1MoEBuM45MFTk7qtdwZrwRoHgteYQ7k2Xuf+FC4JSJnoToVtZECgM4Lkie
G5oVUjhNPQH76VGJhBOoSWe5CBs+inBp/EUKLfTpsptvKqcy5HeYMOSFJKWByZEG
ekldl2FNi7cT+XAPhsOxrDI9THmjk36WXuOh2/gqOOGym00fpRlIrfcH0dHyXwun
HOHRpGfGofwHUQj57ZNXlO7u8wuAuhoc+KCoTeQHgaHBvn6+X5NoiBtR2EVSzXnX
TaCbIO2bScdgUDnAkU0wI9zUOoIadKroNMpxKK/cNZ+45IoffF3b684ulQx4LV7V
2Jl7k2CXwEVvx0hd/Cgy+6v3PKddzm2GqfUCe5hFdxo95pbs3D0TTSO3Y627FjME
2OkhH7Gas3r2Q8U8vQjvBgHC8+bmNFGMH5YXqbVL0BkuAXq1MVaEKB0k0I1+7cT3
2xwhNHbJiPuwBwBmzONwKUOvTM4/HCRqYSJndLjn3Kxef3joUt5vIK2J3B/jwVhV
85otJHAfCfDvQhh0OcFguI5y85z5WJlucztFIvZkeZVMiyI+0sUbJnR7RXyZsk5D
RAOPH+jR332g6J3jVu647bZ7ISM1Fjbw5iylIJRNbnZAGZ3cRr5kx+SdF3I2iWj/
Vc463STTumyPRf3R0eSHxfQzVsZKqmYns+NOlePp257bbbi9iInHEP37pzQiu7mI
hIkhY8+QRTYJKmGA2BKAIF+KXmxGT9pquG3F1YBpDuH7X6w7LdQzQxHnsvstJAXH
kDKJxvajgWUWygxy1LGwGQB+yPjsnxPbuwBhN4tKi9zn0O32ieWlOg4GmRjaO+Qe
7v8xybVjrexYVap7TLJDEFLD3lzLIe3MEaP5Gm9TU1cGsixkMs0HGqM/4hNOEUPB
nDTjp44f9ZB7NxdHTludfKx1uanqMuAO+a33dwLMwBgKDBZPqyODrMJfbVTEcXmP
JdMNmbL8Km+6k/Ur7LC/DzPQTCCi0P7L6qv1BGgOgTlrRziP+Fv1+vRv36FiOVSq
r8ZeOYAULSiiTXIOwnGp0JI7vEz36KZNJvjJuWdhrJazRtPSUHyXiZX2FCWXgUyF
D1aVZiQGnVcIR+CXoukWE5l+/QqckNZZBnq2erCSl/L0KgDm5EyvtWRwhPGP7vWV
6MJrGqKxnqHPVLaYaHfwDXGN+Z1A0vflYxjIQJQXTjCzCPID1wVKoBPHqjDspPGm
rf/dOy+9p6PaJ8v0ixEOiTEPt9iP4Hi1dLbvYHdAO7ltA93FOLfWoMT+NjaJi8Xj
yq57WfgslTpLBiRpn2kN/xhJ4+2d8gm0YJL0gYNpB3/qDv9INfW+kb6uskWyGXvm
cof4vhHD3pgaLl1DlXltwUtM4dwZ4mOq1OCpUDZWFSjr77hH1SmFCzBWQa5ISfYc
hNFUCjMG5GYoyf1N+gnw7gO8zda5AV3q+dBysZLt73gPauHz0hhcqTXtE9ub6SDO
ozIsoQq46vuSNkgNQTa3Sv1N7YvrneQOmBWpiY5z33zZ4pwEX7j5r6hEXgYlQTFb
5c93315vAitVEb4CUUZsmWuRPR5fBC3ytLGvz19hdKXyhJaO6fzgaUC5VhcgmfAU
qUIgyAyt+vfF2CLqUA1AAB19HC77Ed53MBZwwpFf5d8N2SOEOVCSEp/6znWxDUrV
bzLo0ZK2rlk2h22Xi+9EgfsNWEf8DZN8Iq7NSwjKSR6fBE8Fny29HmPT+3M84Dew
ihZCmbcD1Ldjjvi/FjjDI0bT4IJijD3v0KJu254B+VcI2El72cymb7BTfIEAqOJQ
e1G9xqwhytsykjnKXd9kXHsKyvgZCaMTI2CfsCmq4sNfVHeMBoTTAb3EyMQ55I90
uGNgMk9mSxwmkVTJyZhdiWB9AqHgqykeFiCwb/410Y9d4hUljdmWh7bacn3zTGHg
aAcfh9jocoxEdBO7XLrrqJ8+2DJBjaofJHr10cqoEA9BHrWj+SDrk8ui0JTs/iO3
ie5cJSzjmUFoNG3VOEer+PQL19gQjMRRwUagTd/2tQ3cs2To81cJi1wk2zR4aI1S
JFz7nHg0w7KCj9Pih6fPElCGmyF3XGUSJCHHknUy7zcpm0TH2eqPndx9RfkX1NVf
B4RjWYkW2EG36rFJws547nyQNScFKOVw5BYoSquMyGNIz5L/x7yRnC8oX8f/SNvq
Ly4YPIpStehMHmJYuw0BIVZ2s8z79Ps/7g2Gaf0GdnwIUe1Jk5tsgdNJHeWvIqGc
t253fxKGHV2aHCUhHyW01IGSuF+iMjURYKOFZl9dsNagAfzHlSSX2EiVl5QYQV25
a45knUGwKc9Pc/tUS4xTnSUMmDztumz1wqtxUpXMdoRFOU5418trJfMoLaUiyboG
1qvXI1ZQzzCNY+qK7w9WVFpkiYzLHwmWVal+8WI2Q2DM3CelIZpNuXYtohGeGGCt
RfmHxFCIebvtSa99HdEfg1DyQ+1UT90PPSrdJgR7wyGWCpqP4PUW7cKtmHX0qCuj
rxsl63qza0U/+qYen3JcH+oxtJM//5EC+W3CvGOuxTjNceRFP4j5H2h3IZkoosQj
i3SNyusllbJRcVozMZ7LkF5l1AlEnLUs5/uGDhFAl33aPpKCT+RAzxdq3M3lZWhA
ApFTMJF8XmwmqjN0pLe5Amq76+jkUoHrLeGCYCIgu/TsV57TmfW6j8EDeT+R+7qd
cxnahK1CViMARRLnNVND7eNSy8TMUCRshhQ7sWdXeqWPI8O/eh0d6hfnxSNJf9Sj
t2VbECa13HZFwf/PxsFuBar7N8ZUGBDGhyyrKKCLq9PElKWfA3s+zS081N1EnvcR
0Ip2jbEcfY2lT2D3If7fN/r+ggzNxFjfQqKjYvejjpXX3w5+Z/AaIcjVt0+HJQGj
iY+BwGOPXULLViJFUjljqvx+RwxLL5b4OnHM2KQHg2rVQSNx33XFbD0BGuCiIB8C
NHHCpv4SSJB3pA52teAFB3DZHmyZVQGPSBlQiK9jVF4AhgPZ0UlyVjUzhdR/tjMW
TM/2fbDTv1z3WDGHuK9ziLCioxf+jiyW2FUfXDWgU/JAibA94i948WzOFga7mZAB
lsiI47VSIjLyLwrWykX2nkAh9OTYGn/M7X/qc5dBWJSqJ0lfVdi8w4ZuJkxC/XCJ
7+1Xb+4JDBJJo68B45TDr4xbtIjVE3e2mXoE5+WTNnG5pUwKDFi+2aSukdN79Gxc
c1IesCOAWo6d3SNb/v5QcaLySahbG4rX+qbp4L2MWsyeRfrv/A7CTpSP6eNVgbia
i+Mye5SDllHceNRE+PHb7Q8nbVd9Pzhsawc4PUh6TOdm8nuCNiOoftJX33SwkPLJ
pb1eDv5adxq7j7Bjf2KACPPMyTPaf8tnVOHteZDaGy6qn5tSYuSlfukTJmewmRE1
e+5/Aa4mTVhJc01ISvV6uFMODvHagE6vSH5/DMv0FI6R64MCBwvhUcKo8ArsOqms
r60QaASkwuGrxJI5fMsQH41HEtSS+ju/Cypx1gOMiOGJ8gPO5IswhfrKme1oK3RY
e7F9+CRoBADQCDqk2YIn3pwxkKEdpKWLplT6dARJQQ4fhhDRACAUyVmu4n8o/r7+
nfvjGAGJ8F+dacEpGiUKDl9czdy43QPQSPwsafcOcJBF4bSoqN5VBClbmA5pYHCB
OUpqLFyeoHcM3MDjGsC7816qltoa6KpDojxNS2d0InAY5/3HnQVpvYoEDxcX5o79
3GlQL94cW12PGVAPsXNaC6pkFlI/E4EXyUtCWc4p7XDfSb1aJ5dOVrGrGA4JQuwz
cJE3wFrt4FV7sDET6VT4ENyyiwtRWk0qGaF4RNQBLKmKgjub9tDBKOOh+yfeBrhp
MwKD0B+78tV4yzqRYrS/G/3fGAAmVwKgyRnS1+JuowpGxWImeiiAyYiAC+VufVlI
udH0sadRQ1leeGlg0NFwq+pDL26y/pRNgI78xGEi1Fd9aWn0WOHndjsrKVCeiKFj
AyL15eoj0EC2n6vm67Arq5lXbSvHx/ve4Kh2NosX9I++rEvK99rHsS/iJfLlwcml
dfJ0YIV75qNqC30bxfQ9bvvrJ8PANJ7I1qlDCj1CqYOi5P5MNha3XHPKRNWRfnbU
ZdK7kD57+FDByqG/kBHRmaoTLm838kLtL7ZZop1Z1LmeISdib/Mo+C+dk7JLRZyP
0BAcsTpbhjcOfBW3sjGoTRH4aUB1czTmi4bFnN97CtMjjcvMJV7M8iRUSFKWJfAy
THNLkcS63bQMGHu5xgDom7KAWDzNjOYBzGajWYTeINSDuihc9tlpVik9z2JmbYk4
P5YpMWYXwSXxBcL6/ibEyZINm1adXVjtYYn3PslGheP6TFpDPLsdxNy63qIGHeIi
y+xT8xMgwRLI5HXdcsTQcXCbGCe7VWD7vtghzZ00wrSKL35pNXdX6bH2M/yM+mek
F+JISvkVbh4ad8hTZLypQTnFq14NF6L6k63tKi52DSYna/VTJkZeXiIxMcaG6uJI
BpxlZBlNN19ANW1VnoIP3Flf42Uy9VAMHRX3usa3107mCx6DxPVu4fajpoMI+BTY
XShZ8O/X4yrY89wx0w/lFChDDh2hM4whk+Iul1624RfTOnWJkx2IUUNbRvFOoW1Q
NlaKbRw3LHHgrXWt+XQSwcZLtvkmJNYk4h1PGHa4O57qitYrm5abHltQ3jLRmOgF
mabYPoliIVt9sBq/7x/SHHDOnprrT2FI4KpcYndSN8iZPaI2sOaEd0+PnNWNZ01s
JB5hA32SJXuC9QV+XM2TYvizPzXdnc0P8jSWPo3AI3HmrVikNxobbPJKKrrP9gn3
fUQIVgLdX+eMHG1WFDj/GFkihYjKdhIjb6I0TWt0LKTfoSwA/nhjmtaUTUWjGnXG
D9/KR0e88PaznaMKz1Z8ENcsjKwY2MwrX3ySPS7BYDVyQg1QimxDlc9PqVsneqb8
BkONfLqNVqg+B54/T35Az6mdFD4Zw0V3Ou9W7GPDxqmvpuOKqsFWEmvCIM/2Z7y5
nLyCtfrAb9ZRTCmINLTzhvhKnzDrjW9XSM+0vg+NEpwnyzbzrdmk5K/iXXGCb8Ao
Pw2++gPoOOKtKAKPb7VZF2LwwAInUBqAcKk+TIFHDeZaZJsKGjWLfayc8POp4JZF
ksnOJwXKb6ptq/4Nsgg1oI7/5a6mqa1KXFVdIi2y9+KN6TbCLiNglIG2PyoS95Y9
LZol+teXzsmGiVPz98RTDatrl30SmGOTmT71ax0ofWqKgd7FpUqtLG2WZtYMCvFR
MHYoefYsPgIdOQrqjczRnswe80629F4GfOBifS67QrBMkBw1sMcb5Kb9p0jOf4hF
+55os455Cn6D2PFXY91thCZPQJTRRgFXR8oPW23MghNHBKWDTLDs3D90gToQcHqB
fsjqk+QubDosda0DKZZRsZ2EtxdLcpnEVHsXLj/ciIZW0MvB9T+1QkM0hGX5tnv9
BRY5b2rXgOrBzjENc5d6AjnY4UM99BlPDqj8YaIzfHLGvY9Gbx69nhMx5K/rYTmh
Nso1IjYF0+G7hTF7N35SxCO5BN5eJvOluNTvuWuRWbZYlxuJLZsUDDt0Roxj4RSC
DCeKGO2137XNkF3PrZm9D+y3LuIgzSutAsvGLpJEgPyOQEcPZwalJX9o7LBq2ikC
Fu+O9OuQv8Cart7Hf1tsATMX5LfApP9X6uMldFGlbWN+OqD9X2URJ8w30wx3D2iu
EGdLlUnIqW9TkwCW6RxctQ024FY8iPpivP0iyT7z0yYR/iOjvrOJ3TI7CBMoNJUN
PCcZnwhI1pi2vWuTBZdN7/Tpo4XDsH8/XDNxZB8tJIrxBHZedjDC22Zz+hn0tLOw
4nSVjAH2qDxVP+NEB882eVQySnOjsVcJnH6HIEAuyek10nIgYyb+o4CW1zuexx9/
TT2O0j/miaqohZRxmdThP4fjwYzmVVUPbFRmxB0TzBTcVuChC6BYN1L7fDK86eG6
hJUUv6J/QWY7QSHOJKcpCsQ17T8PTy0GVcAk9qYjDHSylPx11GSXOWWx6OG69x1y
TjPT3AIkw/1Wxt30nppej2zPRZ+H0pch0lnllp6Toh8uqZiqv9HvOeh3hEGE1ZKg
2HFydQ6sFRPosyGbN6XkyleTqV5P37cqqmveIGzNRhKIR231cALUBHrC0NAyzrSV
qxRVVPWq8TWGdpYgRdNBLyuSb5dC8Veu154a801T2bTnR3twNOq3pGqHNZOJkRSz
vcPgSBsZ5YAQN9UJL81otUu5gDTzI84XrsN3/TmkN61qAQQNhQ8gYlZ2NEzjWl8q
6922CB2/DnizKEoRZMXGdVW/+aSoltSUjqJfe54qoiLuguPWtDxFU5qEsEUf7okm
0gQMznd6wpW53M3VIBaEGU7wjeLnVq3SXJBWj5MHYi+t8ZLJy4kMare5C18xX+Zv
Zl2D1+J7JeUffFnWJFsQeCeKvKbx6snCVfPkp2jtN0UZjA/Jky41pMjEh7wJ+7S1
TNqIG+OGZ5wGW1+7b7dEPyBmX3Zl8SRSqo+wCxdKzWJYpBVfA9QYb79rEbJ6mB4E
Jnfn8PYgLzCLSa8jZT0Zd9HgqM2GTt43bQCqGHeIyuslpW6NnFs5MeHNaWIs0xaj
QSig4nFFbNYq946M1hjCKL9nDOGshkOxHBaST5DeuNnWnX+Q6rZphENyk6tTLLmD
FZc/vbvv659R7t+lf28WrE+pzYpzBciIxpSfRhTmWhoKY42H61VCfcLHWbnVvZrA
7smnO3H49aWQG/5vknvg306ThSE9y1amN+hUP1GuMujblmj0ko9uL1wnh37Gb/km
5zOIplcxdShNO+dC4Be+i0uDljx8zyYNN1aAEk/aEqhy9jd+7oTrSUafb2hDRCat
vAqxRmnb3F0AXgLb0TZYHQS4750rh6BFJjDJalKEffzKPVELeiyABU9UeoQXzItp
q2Zt8UAvLf/65aNzHpVTMtG7bAzPkP3WUU5XW0D6nkEzn7k42RVdeaGQQyenk0ZY
cu7qOd/XlQVQLg9feF9VPHlc0yvlWeJJbbd4i3HrguVnf/L/efq6t4uqvXePA6HO
ro5lKSunAJYRNkcRJmiGYJvekVvZ9zT/KzXLIc3e0pGmdl2uhJo35iLlZcRkOzv8
PXA+L0GlW543MIDVJhhOxfaJdYw/y5RdtD7561Qh4M4QsnfZ/MHzBAJqaosbHS1B
cOzjnnYWHIWjpiHRKhOdWf3UrjzFRpq/RCW2r4XPiyMi6aQ/R3uF02DEhRdCrOsh
k2vMcAbJ7ae5lQyRZDBkjyHR8BR0Ppcd56kOCBmRzpb4/YmxjYM6Ercscm93VeQA
3wwy1EYLNmNABGxwMBM+HcDhdSwlXAYsNzo/MCLgqQH39KAKNfw3cf+OXuAAYcPz
RZFkJ3qnUcUE8y0FGHNzfkNXo8x/XH3+NfupYOdDo86rPb7FWpzwMFAXDfpblZ79
Nc+hklHMONgQr/VNT1b0YxBpabMvDyNNcJWluVvds/wcqPkT720vUXY2SPh9mJo1
VxaZRujsuheFZWx9a/d9jExwJpMserBtglprrVCBx2V7rytvFVku0TDOQPkKilFX
mKX8nwFCuWq5AMqiKb2Wl0rhfc/xahuqPRRyl9QxTRU2BY6562m+WBRC0+qrRFh0
l6clc8zP7yuCnf4D51fdC39hbM16obEgtUZuKWTpYjv8JuhQhR87m4pjjN0z4XK8
249m8J7TsI3ECU01XPKmviWqyN/p88WBENPgJ34BXP3unuNvB4UCdaKg14prGvQH
pDIw2Y5Gc2+L4e8HF550j4Ra5C6w+vsOxjgD/vInEybOOqWr6csMpQgm3bghae1j
1UJmrtBXyQTCwlSxPjocWXGyHfK2iyYgW5YeSWDL7WneK09dx7j4ToiHObmFgciT
TSO3NBdBjac3iBmtso4F1nT6Fl8+oyE+iAdZKebM9uVJG/4saSXsmeFyPR3EHElx
EgBKidfTT7qr4aMTqaXTrvUMo4gRpaonOR4mkN2e6lj2FebFCnzSoj6ymlm2sFf4
CVOiuyZ0bV2oI8nYURXGQScMns9KopGEaFJdS62szqdl7We2lJCnGjjLgqdaSyyK
TThGw5TCHSdEMDPbjgU97BMh8RKIm5XcV2f3AIEP6s8zJ0qompjpdSKtK2GG24MB
tO6cB7JMHPHulOS5dmQpYQQiJM+Lx/Mg+Hw2Kar5LJ1y9FyW5xzv/tqBa3BKyDC8
188CWA5/NGgxRmLWOb1YUVwkgdcSaKFERL9DjPJBepvoIsEWe5h0OWuLANF/rZH6
Jsx3mnlTWBECQqTrKJjS8WdtZz1ma/W+U2T5s3e1/so8Ix0kSj5O6gsHXCTOEnLi
fiKxp5xlf8C/+Pr9xISPoAOTlk2R5V8Ils+KXshJn8QeF/T+uR7Ai/u6PJPtu+Rr
IUk/xzCNwRBKwZl5vLxkpiG6TGBn6rqtNVXsOiqOO5EfElgniUPyettyc/IzNAb6
rstCCSm/E6ohcGwdSTEDNyZbpq63nppt8BfldQ6vHRXumw+q/QYso0VqJBpQF+9u
gCfZTlCvYT+7cBVRTQFg57y6PW1YeUp/JwtD6dXFebMwyT0RaaTPw/H7++KyqLH4
aSl5bXddtBnZGkfXhBIl1ZpKam2/n2BiOy3GchUWwIImoJD6VqKHFommm6nsfyMT
waBB9tqxeyPDx2jh2oS+1/JSEnrVcz0SMaHxzQHS3dTbFSD9BpJbR8hKt3JD9fvP
7YdC+Yxi8+WEacYGW1+wf9nMc9/D0bxHF0aY5tbaaqLzeASp2OUcWeNuAGj9ansu
Ql472bONQNLmSdt1G2rs1ThpUgXtXh07uKbeHX3Jn6avLwHP1KxtvI2G7Q3wWr2L
S8vpMLwrcowDUgQUIGmL1g2kOKfzeUZ8y1mpGtPahr1Zd8h/Vxx8/mcZKQ8AHM5R
NdSxzxsmA6X3Z5IlFyxOE8GOsgNVa6vteA9AfrmOWBJWcXG/QT6FcMqjvt8FymPX
VSl9tTpLmKukfglgm+Pus/YVisyOoQssfdwvsLQnGURMLNQydFw+mVsITVuFRCb8
1KX3KZkL9AeOhuW5ZOcUsBWVyxXK8Zi2oL+aWglqxkYgLdPx3evHJm5Z0YBu6L4Y
OFS2MCo136BvScawPF9AkxAn7SpIHKMSmFenniyE6M1VCpnI0snoOf8diWJ8Njfe
JnN440KkjDngRzCiIDOWWpbqJHiZSGPUCxCwCKJbpf5Va2nFcxEDth0E7O0zk1W2
QryUPnGnhVQEijZf6HzpOdlZYTfZm0jNNgo3aFx4LG1/WfpkvNfcaKF6UjiSL2f1
MKnc46HZPxeHvHclcnrJC+VAlVI3lf4c9MAeVw60iaQcx778Jh6nI5l4w/BPD8Vz
Q7nzKo183Sc6WwjT1ufAOITGqo2Ve7GPAoABNaVDsvz3TulGsC7ipSADnFgFaxgE
q8KifhlxN6rkyGC0ediqmGZTDQf40n1s4GHS55HkcU2IeHIlq6I+qzQbtSsZs/Xe
weTAQz1X0UOp4H0imxpB6o6qJSkoDjOUZAL5tnSvd4hbwk0pUAvwpdNyM0Tkm2QN
PbWmhv0FBNnI/HC9ZSHvwcOjrEPLo9vhiy89Mtn92qxehZme3Qm2pvAK3c4GpR67
P5EdIYoJeNwnzHkcBEmXc7pKYKyI/EoJtX8O8J/+S/lp2m+5mKJtFsOaxLdWoN8a
M1rhEuT9IHeaIQ5oGjkHkwzWX/kG3Ef3iL3R6ao2XTXNGCJsxkaADMYPedBLzqPo
FVaPKAR2XmiAR9+euD4/QArSt83LcrgA/hvQnUkgL4o3m5+uX+Hvt5Nes/gQJEwk
EYmpPFzrqFr3rugNYnTxg7m5MART5sSZijn0NmHhxeltKJpGq5bNaR25wHtKdwlL
A+n6HZAkBTKAv8ogLOEBPNsUyhZNiHkyAnUcIKAnW0d6PAVUokekrAqybNzEDjBA
t4SLNPdy8PfBWCDDnowpnu0HGSm4d/B2UFKQxTzzHxisGqZR/Mn2DBiORq9yzYru
UwPRztkQoNL7gECaXukx+uBgjmTMjjDFFAWb8Cy9pZNsy17wuYLd9SKsP8iTy46H
WlPR6Nbo0Fp4FHsLykOc5Ot1nw2o1NNMB9EaqdkfmBiMTmt7iFFaGmIn+IsGlwxj
SGmqzO8342DclCgiAzKUW6aprl+hRDQLUQViD6rGKRf2UDz+ckiN9N20uVavP599
+tpzwD1lAegAcEnoYSTBvN79KA8KwVNuxW5i6dmXOFHLJPP1/1O74JFXirpSXHwG
NBt6o+B4kjk5bNt3iMcPUUFnaNgkh3NQLhsKrAE6Opau09EUj8R729Ac+7hYLv9t
k4XTOXjjj9KnrlQehAxSMn+7qk04wxB4EywHGjZCCG7yX06Skhh1FgCbTjL5oVxR
9dZAXnvLiCkdDx2RaL8vZjIY/Tdl1KTdy/FQ7xrvYCTklVlcEJOL3TAqtwMTimwk
xnKUoErHqa8H8QVLqpLz+AMNUtpPjplV0X8YldpnVXXohTA3CU6fiDJ7uY6whiMj
UPfDVnsn+l9z7aSpnB0iHFH0eS2+oKyU6RSPy+fyUfk05UK+nYTsBkDpEFAg3r7Q
+cbyT3cwmmo5KgShj2/9Vco61Pjz9tcZauZgU+LnxGlm66Af/z1lsS+Q8N9ShrMA
CVpZpZMB63rP5jVpT/kRYK8U/HRjcgb/+i+qCVwWrAWpDgLLCABNbqNds/to0JLv
PlfcKckcdNJ24gYxGlK7bKpJEFciM0z0xeZ74p4zJiinI5tzkwV2rDGQAMReO1dw
6XH/cp9e6VzPluwVkzL0hC/mdP+79rzA5lrvQD0hLPUhXOpFkgI4hvIDIK2Oc9AS
a1tpVzkynUXrz9F2izAcSrykKDbvkr08WGOBEmhB1KzsudiJpQfPv3jCC9+zRnNC
Zz77f4aVXkgYzmkjrJg0wENUBvHY4yjWRIi7HPdUaGTvb9WvbpzN7cof4Vnt/NGe
GRttK/BLJNdyZisTYPTjtqQZSUNQ72LyY9P8uBiJ5RVCNW3KjBWNZbdAmeBaH9Q0
WQVyolvZ2I23I/xUNZPnu9ViQGUYZfjen2xnlYRl3JVtwwWBWe1E1yvCK59o5vn8
yO07He0WxttHgyySzwpJZYaQ2FrlE4NbbiKom7sVqbl7RkTlPRwLqKyPFgoG8fGt
+wq822hyx6+ErvRVKnJydhbt2MYuVyihgPtPlRe3Jlyhe0h6r3I52svewc26EFrb
sEfsnkIFHDGqMVBm9w4iuYm3EHsc29oHOJ9n+ItpOkzBXS2grEwl2i1gD+Dcn+Rb
7tvpgjQk7L5umTLuxERm5zngC5g9wqdmyd+AFbMS4IouZwIj6NgoWkTrJJwYMuqb
H2/s9xdY7V3hl2PQJR3vWwRSORUTSA6aK/TsvMjLGL6hqDFcyPKhaOeB8Dr6W81X
Fot47DPSqpzpNEBrO/U66iz5HreDWM9abf8e7b+NXNY4eyDx5Q0hu7BLwCOStXER
AmZmOOYUAPQkURFIWxHHG8MihiocCXDmxh3oqhWLrGcLQDCcLJ69HikJzCZw4elF
od7CGzOcAW0B9k5Cr4/G41SA2INwFvmnxnZKA01XASaN5MLm/4aa2kpOWGXRNaWX
3+s9VzZ1a0np9CFcbzyB/Ph2Kzn6SCkaRGfaDBbiMW9ZoWIkUsDf5ptRd3k+9RL6
WzcYoehK1z+p7xFUH3TQ8+Op8utMmalx5cQ2c57RY43RdQcApqipTq1hPtqJMdLM
UzKlfHPRkNtGuUpVBmlbLJkmZpcQUNzRyW7gmmnk03Dtafk0+7mCbJ6Eoy7KZLNh
zrNEGBSyybZveQsyicHnyB1x1LpIGjGDNa9BbMBZpFpPVt/ux99MLWT6QFGW6D23
rOCyzHZ60iCPyPp4z8KENCztyCtWQORcnhjC32pZsWE+RXuKjpk3fWSIIUo9/P97
cgFBeBT/LofJC2Wz/RdWiV8gXeA48rl7VlUVhQlcFaSx9QXWmWOJ6s+jQPBw70GQ
R/PY6GVUJbV9lmyVP8213uLUOLKiFODqcsslYB9fKpYzsc2bzEy3GjzsWvaUlmSD
5Spgpk9rg6f1ied4ImGTU+npU4IeaI4nho3l34xQ9ogV7TjlGS4v2d+R4PWhOYBw
2bBWjW8/oXCbaj7w252j4BECLtngSGb2e9UocGLC4NkstiZyWmFRvLs+ariH/OjF
t5WKvFRKfKKVlJOtD4RRSR8v9e310wrkRK5wZCkbJg4LKx+PLOMvP0GiOw574Jxd
25ykO8ou2EtdLmK9e2UvJD4rPMcDfgS9KGcu8qTc+wtlvD7lS+EufQnxBEprVl2c
XmGYJmcRw8EvW2JsSrmKM0d64EGhJqcs52v9ahhhVAUN6pj85BRxM4u9Meu4ahOc
tlGSxdZTUHsG4P2mgmL0ZknWpXM2sujkdh2ySFy62hL3piQB/a76LAwupKIifrZh
Yfuyell7qTqtTsP/d3V0Yx1opovs9SgRqCugaEr4JAnRc4OXnd4SkB57yedSw3EK
5smWl5Brl+zKK4IkKfjTRVU+VSm0vPM7P3UNPRdgLxjKjSgfvS7iwuWw04QWMx8i
gqPkR3RNsFFzpk6CWRlwzSMnR0AP8PTld6zGCkwkmM07sG6fZ9zc85pyUDlocR8d
ieP/6QmOjqVPu8Sdy+89O3qGf04uGrzyYMNoQhu5omPWVZRbAk+C5h2wY0wjiOMt
XJmnG/C0uXqILForPtCNdEaBM2Wn4u2G60NUjkRBJTEAcCW+yD/Ma6F68FXfp/fS
3gY5IHg3UY3U1AOoWgO4aVhf6bU0t9jJwRDR+iCBjPGVbHXWzTebn60ZzETol9Aa
X4620GZ1VUOBbGJnE+sSLSzhtqUiHBSSkuqqQmOAVIp0sjEI9PrDRZBtqDPjyQs9
SbAJZiyhhfEsLODF+9t5JZdAXim517CGQF7Q7HhW9vMGWrjRqCJZ3ziiQClVZ/Jm
ggsKoa2Hg4Vci+eGRuuxvO2vJlTA8zMUUR/JRlHg84vvaz6kIIqNm28tYLdlNoz0
+7RORtEp0NHe3FlBepWpCzBZ1LvFSU6X7riaqs3bZBhjE/YR7ezWnHQqkicr4FD3
VuBHX9JZXzLPcIyW8/wJUyWfZHFNRYfmkAw9QSXKijTiW4qgErCTKAsEHIZu2FcC
n9ASP/+92oDVUapgvl/l1f3MEw3ivg/pB27nTIexa1aT2mJAd+FnGEcYjCwOwU45
DM4QzpqLPUmdWcOL5G/NK97qrVAi7ALxdKFdfSDZxQ0TmiCSjajCl46mJPjSnH76
093XnE7qATS/oK2XX7eiydq/YiYCeQjWS/m7eLcBo7Fr8zPiwE8HsvSPfcjbQVJh
vwzQVRFfyYb9WgYjcGMts5y3lSH8UCmtZij1az5y3Xb/+ZXMOmnAicM0epjf/K4A
Pa6gmsWPpDEbEZm/WVnpEbdb2MSre0GGXMeO9dZK+sdNiKZN+u4Mj3BLGwQDxKGR
n9CK8cIaDzpEntIzmRjeNIb1+O/FBamlfq5fYVHrcuDdLXuG9OO1RXVsiD57iLii
bRPrGPN5iL8R2+EtFLypYP9VVKMTrKzOsI+oVgO3L9RSMqlulGeIHtDohEPJAeXz
LBRzjzoUq5mEuXMceOsr1zlvpCbiYXyMedq+EVf23MAfsM78lQokX+tzMCqdjed0
2OboikOLd/9uN3583ycwa0aStfK5Jilhl5x9m+3UWQKY0BT0/5anFvb/n7Ud1e9x
uibjMj6BXns93joj8t3nl79CCE+bnR0qZ8L+A8NPolLmcOE+5xLAQZq2rflm89D3
2mj/YV0/sDi1AH9NnsK7t8qMI+7UBW4fKtJAAhlheWZ4RhWW+LVTHHmeM1zJKYRO
QLEnjZ+yCdPdVjVgcfwL0i/FmEG58tL8wNFglvfog0X1Vpy0lZ3NrXDYoCr+nsAT
3q6lOBfDezhmkH1wP8DMl1wDRZAUAahDCWhJpdiCUtJc91z1DEbz0HGN8hsXn1nN
FoGfta9ryIhBkIozIichCTbKx5M8YyqukgPJqQq4Dh8f4ahd+qD2Wc6cv3Hkku0w
CN1sK4x99etOgzp00bhDfylkt/6dXJz8e1WVmucBGZoc2acuno3+ZxvVpY5+2fTY
eWKPEt3X8lkXzAPlNfAsRQskJW4JI7j464VMziJaLSdBQdo6MqxJfqK7Wm7wbqk/
VN00bO/72YojOT9Hi0uVytYtK2qMwxJShrtHsMifQl6lFcf7T3lsby8Ts4dYIINC
UPjZdDMXVAL7eH1+J1nU6YfOs1GQGsGoUeJHdsDGQylLk90UxG/qupWqNazb91pS
J3uv+tSxd4SUvby9g1moX0B/IiRxK5TfoZhJzu/QIrFkSVQtAqN+OtD2fyfgi3vl
97wBUfwMzYMIAwah7ABob0SdYyTg2nSuMXmg6nFbvR4Isma3qC/zLomKrhqaFoac
sLjnQOaiDEnk9EtimopSPcH36Vv9o2GPgGhxgpFmo02jlgQl1oIH1569w2O1prCt
0IxzMCT9Ufo0zybEvp2mJfFs7aasvaDNy9zPao2XN3u55qyekz8+rrw4XYBVGVv4
XEoeyPC5ZLfRFsOmoSZCnUWuhw7h2l02oybbGaKoppizQmgbnSED8OfL4P+/CQR5
69IPUIHg4MtyfhzLi11QiJKgy9uJA/yP6dLbrcTKvwpcFYl1A0+jZ/4ALxbuPiA+
g+58pmvtPsXI9CVQQbc2Wk8+m82AaA32MnD9AuuWxoaVl6m76c9hfGDQs7hkm7Oq
dlgW5xRs2yak8CPkT5TapDisVgY3eQvhgxgcrPLXTLMD13hs3CGKq4eM1zxISoWG
ZAxZOOPXhVt+VQB1tT0WDE9QX1NDoxEJMfuHuJuDAygA/Y+PizRZ1bRSbc8nwI5U
SjddqMj91teQFWAovbskFl9Tyn0OP9e45n7suSOlEOiOYBIOfveAo4eWYTVhtka4
qk/3p9AsvEG3sMAYzm0VwJHY6uog1N+HWn0ZlHcW3Sat41ZLhJuVeJyCjxRzwrpY
pEYXrqg7dbmRFnCJ4XhPMP26NTsIT94O9t346RROaFl228QVy6TTInyyDqDLpCC5
QEEfXGl4ldx2ijWBvuTvAjiLH3wrxUToeqNtUKrmuF1XWjkPNdhogn1g2qUPxBcJ
01SzIvZUjpMbRo5oNrFkV9DPvB+4NRkW9o0qkzWkU0qtoxIvPCSemrDnYfkh36PU
Ku7M8tcPivPGVYc8M6t1OuwA4I6sAyBqAmREsFxs1mqKk7/UVeMsBkotQSnl0Lro
zu777WcxvrE6pkVyLLTupN7ae5/xp4sjP+1OkVPLmGKs8NrUBwu6MWiR8NAxfI+v
hKlnZgj0XEMV2hhidocoGq62lmNkykzbRikaG1WDjiO6pQxrv59fv4j+vUrQs0fK
gBxaWKJFr2d+Kshe/WZzbOmesjIxtVkJE39qrmQBjZDlvh4muC6yvlMh0EctZ5gw
SItwgLmG/3GW/7fPxpXvcpI/WzvG2v2SV4aci8gUaCyRwMSyDcnpjSt5vFMRHkAq
O4ZKqP1jJsO25xTLydoBL7k2PdLucJv99vWpvKDJv16DwFl1JteqgyKjd4r57Nik
vRUypysarp8qKeVwNtY+gaNcOSm3n8JeKKUkc4kr7PBEW574owS2n2ajDxqAABag
EgivoqZU4MPTRBjFcLO36IaJJn/dxKqy5saBKrq9OY4z9D4Vw1fak9uwgti472Rt
W/o8ksm3A/2/5t3ShGCpwAq3/SBh+5Hp77aRqcYg+f52ji+fkn9ya1itikuf9aKP
mDxaN5DFRySPV+cIc3d/ecl2wc8PdS3ZeaqKHgFFD0QKbIjoTj4fplaZnXxpSrmx
NMV0mXnhBo3XoEtlnxw8Dj9Jdm0d8uGDGcxr7IyNSM4PO9ptcrPOCt96ONhQ0qnU
W0RzCQciMUd9uOlaIEm/PS0eZyLbVXfu+vZjKh+Xfzf5A6+Y8I4IhX9nru75GosL
o6EgbBt2yu/H1Z3sjwySzMEpdZ/v0zJjbII0S0OQH/Zcr7/A0SeDM7bPYaun5CsC
Ck5v9ow+AsE0Cnzx+xg6iZNbnXZ7GGDzhLyLxlVvjQtvCFgYbcSVM0zPPptLjWCF
7NMvnEl+sbTX1r1ngPukVG7wk0VOkGykZMsM30c+5H7WpTK+KOczP7TR550h0k2B
uSkkxooJk+OEfLiPvBGf6fuX50ReGEwjfNN3jSSE4fRPBVvmaMl4DFzYkDPgtFhO
W8cNHgBgaqXBiK2Ws7SVUKL2BL/m5scSLFVtWLCoUkx3eBkV5o9KEpUVnb+qvecK
fbWUAzZrjAswn+QFR0tH/n4gw//NPWC1f4OH/Vl9uzQb8lEDgfrVLhQUlIKJ4W6/
Z1zmRSAkevuE0vL+PhIuRbpzBeWyteUWQ4pjSlVsHhycymKQwV6rKxl46tvZsvsz
e2eLxsBBLp2zAfUBC7i/xrcMKRu06ONtQbEiR4+w10mCCqlerByRaeNnXvudiVmX
KMDCpDRpz1+Papw/sOBS6EaW4QPVA1JuU3UO0/7MW2TrMzkRJ74cpYzavEHewi9a
v7pK518mAhhOq78qC4gyKSEjpPrOZUAskKJzCN4JoluHYepICbpDFQDz/BJdsMg8
Pl7vw9fHYErsR6M1Xy7KGUHRC+vfPH2n08Bm/1zxJdq3J576wGwqbMGnOnTzmtRl
esT8FDaykGwmwUMnBzvHGm8mm/db38IVBgqUFVC2YVqqmGTqYK1V8Ig6EpPBYv/8
8Q8O2FiSCutK2j7mLfn5+p1+XJ9W8JT2lNnpU4Uqpey5sMuHtpziYrXNqI219Nu+
nFppGPDK59irr73ENZKYlDBjF/oLdMTCJnkBkL+LZhhENOF/FNTh7P9z9ek6Emj1
TwFOIokdFRGi1H4nL4+8SiLd/e07bgyR7dSjhR5qsaxjPUXG3xTGhXKPskC4J9GH
fN+UuDFgBjufd4ZERIuJdIkRop2afsxiCIkAvymVztfv/Ahb8O3auECQ6O2RZCLV
BQWvn2M8wCmB/SRvzAWuofW3CNhdJCcm+YeTnc+TjKJukscS8fL8qWaqCuj2HrlB
GvLXO3D7bGWV3fGII676GJ69aNmZktJsc5E6wv7vbRMWBgH2ZcX0qnqgGy/ikdCU
EJuSxzcMY3cc4df4B/cPgNDYe0WNHE4chMQrXstHpKaOm4l+dFqfGkXUvvWWrn16
cdLPt82Wo1LzIdC0y23qYXfxGgMYqjBaU1gwm+VyPA0n3v2pJJvq5+Rm5yqPv6CB
TJ+lZQz6t7MwQ4Jl+fb/KpWYkH9O/QxBgifuQbHEoD9U1TVxM234Opwa9DLgRrBK
ZVQHeZs4PgSjA+q8Z4KQEVaegM8JEWWJyUHptiSaBuuyfqCgQrhjZwDYFN6S95cg
LnvU+Q/CcThEFG4yHyc1EDvfuk1ERpqRbv8+o+we+HgnVluYTidZFFbgZN4DLfgE
RgxyH5QvLegAL4tinMyeoVvCPVzSZTTSnPUFTNeac9PRSu9TehVjGfK0hwSEBnMN
9gcTGyk5Tq2HtgdIfTgj/g9nAXy3Czj3xwbCcNLhUv01FQPBKGvSqJIwXtpt/JaB
EWmUfr4kjOWvlh8s5hSQxWAcZh9/uN0i/mjXL4+Lx4gCqiB1AAQQuKZmnceEo2Wu
TiUPLC85MOSrjeuXqZiD8Xplm+oe0W5YUGKZqN+xqSpGhbwgQr2n/sTb4IlgsmLf
PQ1sIi+CWvaKViBNU5uX3e2qqMemUoBgDz4mImaCdzdoAoeToya3ftz15ZIR8yLk
QYw+egcMGOouZdAF2EanmF7Y+3jIW/cfwO6qKtLndm2hzqQx7Dwv1iP6wKOxxiZB
IQNR+oYWS8Al5KFajRNbhW1JXQn4Brs7MSjAdJv1rABRRGkJqAduKEx8mc7iYrvK
VPmmsW5YqNya+9kGFHIXA51adTPnhw9UxAOEBfoqRrihNUPizZUftYFg9HGkv1xE
nDncZqke4Nc+hRqWl0pfIhh2nZB6SiuvbKLiasJ9kj5mE9V00QNrPpFSWhl4wfO1
Tlo6oLJOJzbwJY01/uNVr8S3+tW852re8kOcGWGi4KffO9yS64GNQ0kLwFmYOYJX
A7wzge21uHYv0oU8v/ZLPotblfZIg99lNMpOTqzF23/+YC2r6g8ZrwvaO37jscHE
/AIIo4c6yAWe+N3nrucpjhSEYYVgkeXc6GDL5C5dN1q6fQETKfCHo9U4QlUomuSf
FwmRmCPhKoBhgWluVUf4G394TYpYggByo1+OwyoMXgJXBU9DY8/Iw9wJAI7Aae2d
Kb7KQHpDyQiQeFQ/Z/wD+zIJd//QYRvtRKwRYsaBfHuH29vPDVkAvGvrnunhqlVz
UI3P/d1Zm7nwevNIX05W6WkTDXY0CF7zdF/pfrafNQ/QOGxaZfZYFxU6VMxbUwCx
mIXH8RC3t4ophzlVQ0fAApYFH44PctJv3t4u6J95PXCSX+n8+T203on5SdPXC58j
YqrYQt2JTW7Oxot2tXbJrsokiXy1PbwEis+LEmQjT3uPdPGeGJRKO9kOPpc/BTFK
KBZALnjK7Szx9PNq6KjKTwqcPHmoTnkHK+o9OLphRf7Qn8lb6ksdVrf/zVGd9klN
j2kliNqnkt/W6PWK+jElfxozNyfs5UDfHj38H2YPvT0UPU0NispmCqH9sge6rhkF
QuP4aBFiRdUqKs780xh/9Q6rklp8NLQW4fHdjZcs4CLYW/qOrXdxqukcMUaoGNXz
ozCctXXCaoF0St6YB5YBujeeaFkn+iEAbXZ6O+OOy5o1LCoCb5M3Le0L/ZFnEPsw
qkJMssvSu8HTWMl3wtytA7W2LkNSfICUQpYDLvsqW3roTUkMcAD8Ki/QjXf8OP74
cztQ4nRbwikCuih2lzM8t/ervbHLnTlCdOgDdEBTd4h45uXo3sG+/1gyCkt/B/tM
LEs7aax39vqxyywW0d12iBp6F3woPNFsHE+W/xKIRzA2649sH9O+ueqHdhDjYim7
AEGO57eKeSnKaRKoUB6XnaLwOVM6jNNQm5n9sRnqQyHThNkzzvijALWTLBSTBzNz
J1rHfDQz4r5ipdHEGWFaagaZb200Q17Y0KtyiyNjjGTRLkZ2vOgg92Muz99QQJSx
VAv73wwswUPaHsDdHU+apHWF2NXEqvvoch9G26nvppIQ02aNASskRJONgDIqaOMc
wWkaFGMiE6YJPK7aKZKqO3jNrwcWh9dSQyF6gkwVxgZWQLLn4v7JVJsoqcghVpmf
SkUbNAu++nGIG/bcS6oCYXs+ZUzre6peBqItr0uR9AmLClBEZEXVGKngQX3zCy16
CahwsoVZJj81XaRJ8pgo1Haz3yfDGGaE2LqK+2rK4WyLFGZUlvlTvbSB6T0IHZGO
i3tzt+ynRsKWj7Cm+DSkXRhxIpm21Siq/CJcqshOJNM7i67MCyX8SYa1numctiUT
ZDlm7yFSzi1S2mV3Kn6PZTwNj9MJt5E7xPC/KfpeAU01VEUg/qTp5g/sPoEwOeAK
vR7a4/9n4ZeEu+wbyIrrf0X1JwDy+edk2mbVsvUM6S9bn1vsCPnGVQf6cB9oiTdv
V2NmyyLb2YdMo1KAgfWC+9kIlSK7PEoWOOTVfSex/PvIumTYK5aU4VKodkLguw9D
Kg1Kw9qoQp354NDDYGej4hHk9eenf2Hk23ZE/vui+1n3bgItBOgz0KGrgKFrBz+A
DF9B3zU6jqLilssrSsjX05nn4zm8Le1vu6SvKiwo8aOicIKed/txrwYny8tLVRAO
INX0aOjftF1gwCewjUq+nUceNSLzrMN3Axqg/D/cIq2bx16DaOK+RvCJgJim8Jta
Y78Te+5aM/Iu6yff6XVudEJm5cUzRFDrUe7hrUvbjGRoKu8s6Chy7JymKmz0TUhO
WjdXPfMM0MDw8EhbX08LeHHlPqJ/VZODTG0HkeE2WdVqgCUC0zcOtrm/eeECcAg4
sTI2vtdICBE1+792Xtj6Ym7VRdY81OXzcrpVKTlv9UINKxNhXxOMQZLRATJLo2EY
mZDiWkC4fwhIgPR8YGSoFclntINPSzT0iy5XcWRlO+6dP5LERxDxa25LBliLYdjL
GFuvfK/namRFdreQPAiW162uimYsruPt3QH7NUKnVVMhLVxhCBxt4tJ2Popfkufh
NIhA2KIR5P5ckolJagQTsimaB58wls9srqnQHFiwoQoqXfUgFAGTyfkYL0KvX82K
uFU4pkiGtMoqqan/Q2guWIXV/DYp/hzXLLTw09d3g3S6OqoTjE3Nv+4VzrD9W3OX
kpRFxG7JN1537nBKRgnPY/qtjZpjxGk6sBacUJ7TgbY82yFK7WKd6mm8EzQb3AOt
5qNoRmSxPilrA3OZ54GDgpKtxr+vmGh/HjTo93+GmowUphh9IgzzY00ZUjcNu/rL
sbSXDXzmZybgPPcNQthvd/5DDRZ1ujMfPbHXIZUbwlWQ8WY0BVxzCeNBLkMdeuzd
OHMdmK26O+eBjj92PhJtCA7f0tYLXGzE67ZxkgL/Urt2YzhNii8qnTgtt6KyccAV
seGp6Ql5PqkK4IADz54F+c97E/H8hGCvuSMcfw+mnDFfE9p5yabcCi8Nr9uKklM4
IorptkCXniB0DFBN71wHWkQZdqBBCKRAnMZVA0ubpuOpczgQ1bHLlovcu4SwmVvD
6iVkS1LI6DnLkkoXNeS+LKRxuvtKfzt8mVNTv4iZkYgvtQ+AXzzHbGWqUufN24ny
5kF0xuseGqkVjWWSf+HSyjl02OZM1bc1Pa93GKdaa9iNfIwqmEnaN17iYoAgMPdi
oWT4aDTpMy0L3yfS5vbfw4UQI1XH+xfCVN1j241Kr8EvUAnZYAUUnQKmqHIUvlxw
o6H7MNiwcZb9c+bo1cs3esGLDxZPwYp85fyYpjLFMopLBo0I/5grCWZUCwx2FdEm
e7TrVTbVtu1FWEB82kqQgjwoPqDXeRazJxyQASvthaDlyM+J0tdhT2zbLitEZWn6
WwDnnb0m4e5ktwdVTckNISqHpdY58ok0D4gGaSgFmUApntyvsEzoOYKXGoByGA2j
TN+YwwMWlX6UNxxXsPWrFMTz89d4KcJoCwvbGlW76qcTPgc+cHzWc3didzDrIh1i
Ufg5/+L42ptKzrzpmX6yDd6GBGFfBWRvirgrXf3etG8++H7Ft134DkQDP8XpAxze
12p/ZyLxuPMpWPERGha5y3F+HyRM2QC0uVVHSPKg7wLU5hfwgD28IB+l3s3BbZDb
wGatsLKjOugRQvC7dzxnwEm/3nkynD+0dsgdXUkX1LYd32faq2NmcCxXGTFr7C8p
SXF/raHPf2oU4ZAunPkI4QYreqbNlGBTiHHgsfgVOCEbRh3RM1jfNUN4PEqfMPmo
nKRPyyfaBjINkcHiqN+TiEueZDNyXqot81mc4lXkGReC4R5RQXM4u4ht8VB5PSPc
dw87sBCcUFuPipOf+Up//WZV1uOMKFkMeBo49UCs9JxNAf5U+x/PQ7SJSCpVQ4q+
B7wXa/X4lq5KajC/uU6DJmKuUmg8m5cHKKXcRS01obbP5aRRw6rfBtVc9enG5eOG
Q7FfxBrMB8Xd3gk4HiCiu8rgYPfgTmI3mPcKCOjdc5oLCwtFJ01bsUJ62q7e0OzG
dU4Zt2XSpNjBjjA0rIYZuj6wdL4M41syXjjozqP4mir38NKS5eJFiEWpaS91qdQX
CRpW8A0JBZ32o84wZymdP3MlePXpLb9ZRKEw696LDePSwDEqsBZBEAaHDiO9qk7z
og65be5t8bbAuT6V8BbgGy5w0H79IztKe8EE6Vpnj5MYIgNkL4bRokE0vx8K5qrt
/f3o9t4oj4YZl925BnMDO1qRZS4K12Km6IDXBrUpX/Ff2KWBzqEX5Nmqdzxa1chf
zsvG+K8JeOmgMT7cW8WXgEH4LJKiPIdhVLfomC+2WvvRh2jBICcfBvzpF/LXBj2J
lWO1gVSmYPUlskpZsp/2u5/4febrPGmvVHIOJf2vvmATSKL/uUsHR4VY8zKqIWC8
SXtNyB3gYNfAalK+zdl3wkXF4Cowxr0Lq+C/BLhbyK4ttQ0pK9b3SuoYPEjwa3ZV
TTX1PfUcTGN+K4CSxyP2uuBjvgufsNUboCAm1CccWFTUgwJpr6ynxRw7L/6h+Mx5
PKf8MFQMWmCO9GmmON7wVQfM5dLUbWCqV7tOh8midgKVSw/4rGmmu8msQxv0SyTk
mUShi/8o9NT5/95sndLUhOmvLY+z2j4lbWw+KUHMbMLBnjLKKuo9QRAJ8owCQj1S
uPHv+ncKRBIGEKQtM3RghwEn32v3TppmlDCMtH1kj+nESOu/Hv2TMVJqf9twz+HU
+GnKSVimxB6Te03Mu3XZU31Ql58+48QKRsaVKlFKSdYgcNDuycGkxIqTCdc0rwIt
TUB997+RKNK/n58Z+tRYNhZ6+OSuRKLNpKGnUi0aOndGhVbeeSMWvVLft/SvZI3y
dKgDcbTNxG7UnbS6oU7Lhkt2HObs2ZD0K0DuGrzPSdU1h2QOAc9+1hHZKhFTbObQ
CpCYYTeYTr1YyNkt4yWw1kI0SA7OUnP717BwHZht2EuW4aiwNGNpZqKvTkHY4rRl
p41tZcfIPcO+CIDlplTNvcajmFgCQFKwDst18h3W3ureOkmHLynJWzAxraLGLHSA
oMp95eagREiplCYpRVI5l5LKEQnIPbVwNJV1AqqaBma69VowGDXFPXF1bQL8uM2g
9wKG6ngvlPDlcJt0WoRoOGSISBfHJnQCjLuy6O563sOrW9cQ5kiEoXnW4k3niMSP
b0T5ZWS7A4anKOUhlc6+/3H/wBfrZdYLamPZM/7AZ58Vo3NvgQy0ZmLsmJhj6UWS
Wnoe/CqMumMsTeF0CSHx2mspPl3HSIfHHoEHAJqIEj2dx5Rw9/6muNEpvv8JIOfa
XZR1MFo+eq2yNja5WqwZ64VfkEeNDz3Caj6Umtcxi3uJWgvBoiFiXtZmswNvpn1G
Y1AGsqQ15kV5cLSFPkRgAlm99UsZFtdU0bveVo5khuiKKPdYY83VsPw0O6y/eBMT
gULtleYtn8WRXs7gqeV3eK06IAgJoAqsmrZygs6RGfzNvslWrHtuw7b93/mhLTQv
x81LMBYBCldkfO6gSNCC6dwck80N3n5qvSWqAVZ7ZPQ26gtTFOdgNv7wOL28SOeW
4RdmexyajgxESCzV2jho7X00gJ78sa/FjuLoo/L+Xv/jpn28kdwNsuCHsRpLEcec
0ni0KY6k5FGxItZXfaZB9n4GKVhCyVuxiCCFKABfSWMxHmMBq8w47x1QzReDfhQp
BQMg2+LbwEnfvfoWGdkYdnh91jGgwgov7V2FqKVvHq7FusqWq8Vj93WVxE9EhLCb
ZbcwlM6F7mnW6engKGUg8vI0CmfmvPTQyW2F7FXzunrRAsvj/sH14rjtLw/Mcb/q
PrGKS5JxAdOqZ6LLxFWzbpILYNkLrNVhD9ZWyfuuq2FgFZS8867CNPqAkvy5KXUP
CbnwmZKjLjVmZS8kYULrDvEKN3V8r+FMwVlPcXWCH2zvfAWwUHvXkvfG99H42tLf
f3BVVJwqrv5ilKuvGxX6MZkp0THdSktsrPysMaPnG3AHERFTt8x9Us3FbDM4/tQX
4SXUDi86CXSvy6rERtfyhfgat4c78v00/pfumOAmb34hMMIgbrUVlr/bH7Hkk+lB
re3GGfZZXZffLTSj/CEly/MUdnZM7s9yjVT0fgltmQK3we670tlHByPDsZvqLyEh
y/d4FJSLwgrZCi0LMH9ise2snpJCjUa2Ueoe/i+UcbFSyciqu1EmL8QFvn6ibmHa
lyd55Ohz0lctzJioKFHhtFzO7UuifCZKllud9QCOEbJmKcXr+DQbqyTxHjGRM/4s
4YnOQoymd+i1LP+UjxgHYd3fPgmRPvOMgKx3eoSk5G1pbDtmk2MUGejnVEsfwvRw
Mwqr215PE3O5X8lsPt9L18dMc3NO6jvF9Pi867U9uKJ56xACY3Hrv+XfVEA+ERPA
ExiLdfrg8/25B1sSzA3img0ChKmxLavGMxutQS85PqHxbLzLfjRzS9hjxOpRB4HT
a+Cik7jCgO4xJz90emsDFoOtcTd5eQbsLE9Wpu2WJ5ztyusyzoBcPuyOxae7S3pt
Y8xO0y9bqTuhuqbAz4D9h3LSTf9TsdAI36aO1AcxBBpkGgc8H4vzTI7AKfPHa2RG
XR5Zj+8ppD0dq+Nh9ausw+3+DFBsLLz2W5V4Usa4bhCPCNjmVdHrzATeqp/lS+N8
fOfY7SkWfAbfznRFn49UBIe59OZBza2aNuZS14Tof9QcGwZWGHuATaPzP9zHYTju
13kL9FHGxNS1Q7xZb4abJdhk+dCez1Y5/bPanZkv4KzEWHSa3OPz6+md8zE7iKl0
Z2bh1ahv7tMZoBYlJZ0bqczqk+EVshJd+93LFfKjxH3VHz+O+QSjSotpuga+aXQV
+C/HuhHyFaJ9WSqX4QtrMosdMkydPIrLHlR8tREK6FTJopS8Nx0ihYOsKv90BzwF
yFVoJSKjg12hUV18I8j8GwKV+t+VcT4beKYbYJ06yXPIv0ElH12UR97Hjh4pz29W
SS8wowfuFASTAjDhyuq95/0S5+InBGpNlP86AjDLJP2p3lgRO8qTaJ30BgAjzYAB
tJPK1EAFiv/50CoUqMlAweKEhrqe5EVrtXZ6SQok5aEsLUDht38jFmv0zZvZJACZ
GMPsoTdlUW+N7k8oCdONxUuhj8bK6lCVSBY38pk+kptQQK45UCQ46J2XzI0emVKF
7zYeb2tzCBR+g60dtrvnDe/sLfx/DrokYG+psh1MKb0bqd38yx/GKmh7+G7O+dRa
q2FQAqVut4RjR/ndUMkbzePAcGFwW0ZcmPWMRYNrHy/zac3Nt+xQbruMOCT+2Z6T
0SPBzaBaayrXEgwxi5tPP3we7OmVO5NAPAFSK7I2DC4Cw9Vxl+fx9IrEqHNy979B
F9y8+24Is8Q9O6VpcsuxgWMmo5vMWzTPVpjD7JIlShlUm4G9L1Y5bJvfi9rS0Kuz
BaKkv7sRi8hos/aiye/NK/oHZXO6tkmzQBGetdkkjYvlJ+TGij/Lg0n+jTYNm++s
AgdoVapEC+9/i0RdQd79yFwSXOD/myQ9u4LkejV+AMyrrv6aNT4DTUXvNfs2gh5d
R6grj4FCgjjsuAdEckzKQPSXsOYPyyuEpyhk6hRdLKnMNPBNwxxGnt4Hi4O8Y+IP
rwOQGyZy1uvEXxlP60vnyFz2IiWh9LVzgzmkinHv8Sl1CkSpTAAlRlywLYBsc14d
UxslDgTylWHQbUbWbP/HUyl9wWSvCH9XfGyOHHIhU+J3PbrcLQ3Yfuw4jS90RU5t
Ihxft6d5b5VluuydJd35aNR1NCPzzSC5rCzIPCKGBIB2C0FvM4ZeamTU9xNbYiHT
+WCnm8yjBtrDVvzNHANmWTrenFl2iCNJUBhBu0kfTDFmcl3HwpfdxfkBSKP3C02P
+D948q1b6cajk+gKObR5ACjLN2qXzudn2jM25ippcbgn6mo0J5y9qVhbRR99gPgG
K1FiE1+cIBe0X7FcTCylnOVdIvP/uD06OwfsS5oThXyKv0lgC0eY9DKDT6LZR4rE
G32faK0hrufPtqeaUXbUsczILs/3mmGPrsz5I1KlwjkNJFL/MANN4MWr1+Z3FYJ5
/P8UnqjCBnmJLnwVhLX/L+Z3ZQOrXOYelqczL0c3iWWOwUHA9CIOxYcPCoA5w98t
7lqqTyS3mJEbCNHvxL04jslkP8hQzvM5AugPOrN5fI3cTgp8vg6ZWuQoT3+Px0uG
8Na3HqEc4IZSodZaYa9Z50qa8ENdPJ39/ILZV+Qwr+KgUQo/ZuhPSbwKIA5tU0da
2oybKa7Yy/F0dqGDQ1/l46KZkey4/hxUPn+G+ufgsGuBH+eUmGWZjeXxZwfaVkgQ
8IFWPz1AAYmX5qIWqWXe6yMnqnrmiyX9ICewSn3YRhJX1Lby2LY9mbrvA/+PKpIv
BqNKUVkOaDFauAXYQuqhoMIsDxuvTWEjBzKNCc/QrNLt8/Do1ZOU11WbgxoGz6lE
opndbYbMIEnXdhFN+H8j17MhusT5X7EOrhUprn26S3DzmgHS6wUFbq5WlFJNydQj
hKJ7wCPPLZpTEMogeKNMphHszDGcKc0wSTrL8bxz0xkPwI6BX0HQPBHIyItITN8j
Ony0X9s3Kl3K1eq5wEGfgc/989qgtQz6BHVBO9UKIlkQUhGy+Pyjr/aAM0z8rv37
9dscpr236PJK+gdT0VE4ptk5u6yQrMuMB4qkOzv7KuWCnznA6Q6pVLzPYNvymZC3
0Wyc/VYNwXUTdB9AFsnKQwimY4De4sOsOfvUjkBJY4fSyfADcQ/FhknDMPDmjM4z
WhQ9VWs4wVp+EGt3fmmtGob2nAZnOFw6q0iws5jfJ6rJ5NO/SD5iOOUonU+waK5U
6+gT/ed/hp4GRy89lrryd+/lL4iNXngnFRwh4KM8IgUkKWudX5unCcwmL8OYgPlh
O4xmdsVWlWEPtg+x0dicxg3YAZukuMQ5U5+HptL22zo8U5ZvCvwrjbec2Z9D9l31
X7SDytWt3pFoCIAcux+LczC2RA9t8uH1okD6zv9LHcAub9rx0DCwD+uTh362TYCd
bT3tpLAtunbGaidZFi+Wa+ApVaRVr3vMYFEUXK57lhpSgxijDZEo0a1uuKfb3zp+
1LLjnOL/b2uzwnX9byNNK+py1GteBDBTq6ZYxO9txBCfqC8JRA5glCCb2oEG68F5
UC707tKZGCySKSfAgeWdMEK4wC8CqoVwUEbrwyWazA0tn+kqzjtSjbjnQKyiJSE7
fMZkQVvS/+v+JhgVSMDQJtToaVAHLA4dZOb4iJgz1oY7811/uxgmiG5J34/dhLOH
83oygF64bz3kXQqIHKcN8JgKfOw3eGYdv0sXgNfbvAySmRLuZCV/KZ6KQS9DVbXr
tJHxcMpd/dBq5tPAs7RwhLVyBYRuZczaWMUS+sUrc6zbSnAZfwxcbHwrZV7/8aNd
LJNxWDHaXkc7RoifPfYPg9DQYv+q+e2RRSvmglIwrd5AdxfBwVkgb/zL/73b8FIN
ck7L+67Yg+ZXT5y5mQ6FV57/U7T323VN3dxauOtIgHRL+yuucoGMP3i+7J3gYb6S
FW6cFk3nwjzlH8eQEohM/skISDTbv/a4xE5IrgsF8UL8svoUk91GsyFqKFKin94e
2AhlccnnUqN95gLK0souZHrbp7z20G/NCNtvArpwyjYckyITpFTWTuNLr67juY+N
PhAOd5i+lUa9YuQtqAlmSdD/cjfb88543mDYq0xtndHbx881g/BAiAoLUo3263VJ
MoAZZCDpkcTh8J2gMNtVRPKAV6TLWvthnVSSS7OCG00xjRDagnjTSrPk2nWork5U
+LKURBZOrTXt16wDa/3Za6I4CTnKxXqD2TFrx+jSn4uTlG9iLeaZsfCMjqyrntIr
zQnPYi8ur0Y92ZsbgBqSfFqgS2R0R8OXE0/NQDmags7snqvjq/nBekEAdxlShTwH
OLGEPyZr5Mln1c0YkmqubfUV9iOqTtet2ZbsJ+9cAAt0Eb5NiX0UwJX5XEMhryX3
pujoNtufTGN24UU32ql9/bFc1cnDIm7t6CNap0ArHhYbvs7Lh0bg1VCTH50x0plb
fVZiMKTV4Em9RkS5/t1jxqUTTepkTouNCNg+J5Vu5e7IQI0wI7soE+MGRIhnPNL+
rTj5bFsSoloe0dWkPoAosDka2W7NOh/4/oaeiiNpFYEu2U0lK2gp79bllCUFYlKz
/AF4YT1GQJFpwqpeo6xSbSTdu6Zp6Cm/smR8lkaYcFwJSf0Aon3pjSRu7absqz+3
2J75S1tnry9xfEyHLQGhnlWLtcuU2I514r+BhzBydm6Pnd5sqzHLutkUWFdEL2DJ
JAfVed1I1RvMh5/qHhceTiMTBUE8w5Rd06WfkvjY5J33ZiycQQjshwfLb9uK3plD
NTc+73jYvB7G+DrdESNuY/4xvy6QyFNE4QKc93fAsxlwpS6Fo4zgLgZhAGtuf/Du
J8m70dMgsNgJZGxuDvmhfm0Gtmgkz9aRT5xUEex4aZlegiyPbxKmrotiNudwfgz5
5k74V3EG6MyV1RdpU6iUNTK5CeawKfUSpUz2BqUnO9Uz8/Ji9vmXC5Cvt96u1Q68
U4No1ZZ0HR55ewu+clbdHd0hpJxA1RjwLDsJmhSqzvz/hwmHLx5O5d38++uwS8wk
h+5dATH9WpVEn3+ByMCdZxL7oBLq43t0UQWuyDQt4Wd8UPGLVG8t6HNI9E9KwE9Y
SwPGcWT2GFtAlYJ9rytztNrXoSCKE6MuKAB0fXz5parqS1CZpxll1gRavS+tO5EU
QwR+Vm/irPUtJqhBzyypeaXesHNGuVOWu7tYHcv4q4Ao6pRKgCDR6p6q9viPRbjm
MUmcxrBSsLaCwVE3BYu9zw5GlBWvBgy80a6qsmQXfsSu17wGv7a3qRu3bR6HxB3+
zdiMqvwCKgQOXQ6NNyWcUHO5UJbOq3IHWj1acbkJ9aygo9/R03kvnZU863qimtu1
V+BBHtqiDhiH1vviCai9+KoYiyjY1pKWJZkcAdvl822qUh+Vhd28Rdu9stFrFaPV
DG2PYatbI9+O6Ae1+54xWWdezNAm1Hi7ZQUZiK8vYeXX+Jl5OqUAxP2Ro2GCT3ey
85Sray9sMUf+A8I0pTRqeA5cvNRcv/O/mUcn3Gy5s3E0Cadpslixd9jXkfqboAY5
W+m2ilMSbjVJYKUos7MiyJa0TWUsVTCla214VXoDYTXidFUACaVZv2bZJdjfdx0C
/KiDp3nPnlXElAGhWxA9UrYWCasnfBvjiIWQ0pLvb7erHRdVjO6wCtss3uL9jmUg
FswKkSACGLzbWkr244ueH/s7VZ/doc4o0DqCl9ZsoO+1KIKf1vZ4HXWN6Iw5TEEc
XpWOBVhUdh61S6XCGUNZ7HQ/CpK4xtUneX1plZoTRL+QF1WDri/5kIG1fBJKto0l
enqAoerrJTEmmp+1H9+NViP2AQtfWDqn5KNTRHFkftNFsGi0u2LpEUqvFjx0onlR
ITeXPJkNkmJL6XpDqBMMOsnvKRwhjZLsqE8q1zMSGCJe9SOKJPiMjLzl2K2rTi8B
mfhvpIgVFqVcCIcAyAQlQA2kIn36Q7xoA9bavgbegpSE7Li3pA02P/8fxORzFp/p
09eCW+R64s3L9J/5bhaI4DzJ9QUv1VnXSJzTeKActphtUp3LONfLwXlwKLF/M6ML
5RGDVV8ydQYJZFtFwX2tMQLu1ASSB8vAqaVwO0spnHtO6DZ08+KVGUXpZprhCKPo
Y3lUeKuGWccNmxlAH8y4bXc2A+bBaDj1xdpmC9NETbET6tLc/UEUXNcTMIGBC2Zw
wJ7FU3yvG27Kx/R9YBwlMwhYaDCyXcp9b4UNTPL3NR6AMk6sL2AMne5YGv4+AlP2
luHYKY1MX380M0NMm5Cv6R6N3ex60cs9WCt2+pVhVxm3aG4dA5NqkTBrMl5SLY+4
2ZYyGg6IznKX5+hxVd0x+wHNgIpZIud/yuFpxO3sPLjiTDxubAcjPgAbSXlkSGC0
JZHht9vNzRm6XNIA73RFAxMrzIrTe1Jzq1mj2gDMfhzMZsQie8HKBKb593ixklKl
1LTN+4G8AF5ZuW14krLhU/12a1DCrK/XTOZYDIDqDdkFY8Kc1P74DAU5m/x2tliE
++JRRZd+N6mBHtU6Y5a/GfUMjtJ6mqyrBq6No6N9zUxQDtRjtXMiU6DG0eBGdF+n
q/NwFtJDKfksTBFgHjY4EQS6GDsRhTkEObJDDc9FVzeUznylPsXUZTdUF5YrdWbW
rq405oqyOmqoUX07z0u4OEWXZhMCA9E5MIuPjYYraP4FiVSQls2lzjWb5Sw2OVUi
FYaIUXXYqTpOzrNUEyhp8zkZnqwITw/JulCt/b/atvxIT79GErE5M5DVyNdmttWI
C3wOvInnSJ2ZPmIsISOgtP/hHNJJRXV1um0rD7BLEF4J3vHZX0SzMYmt4QmS4zrC
+U8DxSZcD9gkRbQovH+0NI7Np8JSP8mdFNL1ZKYliJ9p5SPnDlFGtBECl/q0pHS4
oQIQaYpjKaelO/g6JvejHyeegxgu+/DKmdhtO8EXTCheSdFaQ4UYeIvGNfuRY3oz
ABB+ii4nfGz+jqnwlUt86rPE8CKoy1i54QIElkMRxvdj0PtZV2eJ4EIuJsK3CD5J
8AThrLyY8GVR0sKwjnucdliD6xYgmjbNFTYUywPgXP7PGqZ4PiPGh2A2eABHzQRc
lMK+b/GQAZfHSnNj6WINOITQ4XvLp/jjcmRAo4Wus1s35Ap+Bzi2fWGjWAx9sfQF
t6sG6D/NcToe+0M3qgBFL5xzbF6/J3GUKoh9W/mcczEeCJ2oWp2sf/Fg8l/0DZ2T
wpc0LMmv7HcLx84HTXwB+JMZYmwqqi//0H/5JcpAI6EL6RUby2vFgbJr3ESkF45S
W6mjy8LHeLN17FNKUcCKZ7Xbdyv9lr7NypoBmkM64pZP3blo+JrpWxWd70gunrdF
lInrUD3rHMgs8mrRFLvkh//b8HHBCN1qhG2HZV/TuS2pdsN2nNDttx+0/b5aApSZ
Q/ilVPIpXaaRsETRML8cD3GSkB5twJ2EEEaCeRYlIrqYnlJzV4svK7MuzCZN5XvD
k2VAImZiZJVKSeAWpEct3eHOTlTsjVmddZVCU7f+wTxNR6sKX5JIMS0NbVICtuiv
b8VD6q7+mAAtU5cquc2AT8VEJTVk6VmyvjRSln0KQCaIU19OVCjEkCrazXFkgFld
cWKi6p8uoBkGrz2XSAmxrNsIcfgGv90PbdkpRH4yGCQ8nqJve4OQzQkrFJ3lUlSO
gduvpJryTpkDf5UOjrVPQvTGErTjq2S2vC8iZ7a3lvuuku/ONReUQsQYjARc4NBw
5RYjEwG62Pn4JUdeHUjHO0ECaZHwXeQJrR+ChYfCZcBrbwLN2HpiXaOCha88rkIN
AgP/m3RD6x4CobfMMp1ZEk+W/+8r22quBj1Cx8K2swp8xixYPuLIIxTfHuthdde7
YXJ3unxaygSfWfcwzd1/h7IhNw0E6u4lrdtjFxXotLoriL55VAKk/x+rDrL6Wz79
82TmRyEw5lVIU4pbKboA5EPoYzgaBXnCF1J5vHQgpW9RgvaQiOFXzuoKV2wumPy5
nlHIJ9uggS/KvNKpAEVMfwYfPMpWNkqqripguEONJu3gVLgumWvZkM+6FEXFV/zY
aVldHf7SYeywFoCLJy7//A70hqxq7jFWvUVqpzfyX3Sq5rUh5OJI7aJ58Wpo5y1V
UIotGzZi+y/H187nSVJCQKFY1JGhIorKH7qffFDnYAU9cQUDtz8BZQ7GCWT/Nqtc
o9BP6Hp/2HZHBcHKCGaeJkIWXFZBklbbfUrC8mRlDyHui1pDR79lT6FHElc2N452
fSWIiLz6YIqoLqcEDTdm84TOHkybNkVYZZgTyyahBhi7Wd/ZfoOrpGIAPE5rlJRD
HLtUv8jlYvGuj66fk4XhoqWbmpF623NoniBPFl3NW/BxTJJgFVHSmDwJ5swuRMm8
Ko3M9gTyphueFtQKrRPUEqD8kjIMgu6q3uI3y6zgyIj5OHxuMIF5z23vAccdlVVg
GqKxbR/K85AQWmr52A4KqUcle6oArDr7+Bh1ANcq1ac3WL5LsI51eK/x7WtJlQl6
/ghW04T0ct8C4ptgoqcWBVt6U+9bl/5jZAG5ClPCFL848KGi49MJs5yoT2rXLFOY
VzmRVR8OfQRAulpbOBqVe18MbWrd9DibxEBvcpE+nlHEH9TVKmsQtE5UfPTAwoKG
yqfS0vpnbPm2/uDr7NL0h/Jrz7/8QUjULjdur0xjx7b9qUS05v0nuqgsNEvgUGyP
bkW0gqElzlc62LOSyos7e4pYG5X5d6uc2L04SNanIy1zHdJv+vbgd4Q4SU+qgqXL
mvfBllq7U00ZibXA7wMp3sk2swvjHsjhNjgZ6VHwvSWHs5XLuWYfinwCni7xTh5H
4ZYhPgLmq4hb5Wq2UftvlFaXWy+yjIaggfNa9tX6fdi1F7k+3t08yUsqh+60lMUt
KNt0T2of5K/eBr0l+/+PpfMPpD2WGG22MP6hOcvXcfM78Ra4VVI5WCj7CjFkQzSa
Y03i2At2WlzMsxrg8a4q1S5N1tN2U9jfAKoe5+A4DV8Xf2BMWjCZFLBL3Vog7UYs
LWO5MG19/R8qYDIBUz0M2VFIH1VmyL6h682Z61soKI0K3hJWf7Oyrwpd0WYrsb8O
pfo+TW6qo6v3TwjSp0Qv7EOoK3e/TOdlcvUAJ2TM4r3dMux5oznCNfbB6P/LrJkj
S4Vgbwl0rf87p1na1MUww0FSdpVAUBZU7hXal6shQqyzHOvyq/JLlWSS3o2nSU4J
7yymjDUpHEW+FwZpoG4xICQF8jOTosRD5S5k8zBn/I0BlLQyYJXoUDJ/Lx+l/f21
E5So/6j8l+soujCEaGb2a21XuEsX9i+Byv+ILNtDAkGyqB3/hHRYC2jy8A+qhP0j
JsD0dtQ9lJvbUOrNFgHQViZa6cg6Rs0OwtmtMnWQ33RLVqM9+cnXk8qyXLKSSl7O
NyZENP2Urr1H8815XIXWPm0DWI3n3NXBbJOPVUY/rCYTBsvuuf7AS0d/HGQY3Dki
TZolI6YeH6KGFsJ2F56ZeBmlG5GFgZJJTswmk8jsZqrse8WY4Lu7mrmwLsmeQWV2
/TY4PSk+Ee2K1mqxGeshvSoMRf8FhvKdby55Mf0op4kIWi/Huzq6dnCDiaGGZ4BB
mG3Vpu/UQzKV3ceyh4KHixMiLgzy6nNVjMBNWqQzcnMmk3FKHSbh9l0UgIpK3gtL
VwScCci611oWofzJIYY77MqGukIxEZfgKiePNPEjiRzW6lbxhisgLaM6WKLgJfEx
bI/YeNcmiadC/zb+SPHicVrpBJhRtSskk35sPkJFKHDDIM57TZW0G2drC8hkYVtP
bTEJVWXSVkRVYcbvVbkXL43UUIhRNXBH4laLl1n/KDP2LwGnSHleccajO4YQi3n/
feXtghYz0DOuWK6wvscPLQ5vvcnusCfDJVIIHSLbDL4DriHIkNI0EsJoQqvNMDOo
RgjPfq5JAnB5vR/yqEkdP5S0sDpBJQMlFbQSQCxHV7APu4rOUyYAXPb7+0DWCFDs
umUrdpwjehkRwqfKkEmXr3QQqd9oaaRj0v5O80d6Ax6BK68SAH29XqupJ2ntZaPb
cDY/9qeOY6dqd9Q+4fxUNfFYZA7ZzcPVvLYmLn8fh3avNohbQ36/t1ARK2PJ9PsT
AC5s2TWKt75M/fS6nZg1QhgjdKfnAq4RWSOkK7myDwDnGPGVyuzByFevTeEUrgCT
2Atfls2cZYLvnQaFYL3KKErIpYn+DlqSyQmxfOrOsPY2zd1TJq0gGNhNW6c0bQdO
aTnXOdsq3hUfquQtZ3/IyQoRX4bNikkKRML7ep0rd/BfGX2Cl+thOD7pxeYOs/IP
YZb9O9CrrHAq4WrnJPTFKKEf+di7zO/um3rGNU8dFne4AIbHihdZIJet0bqgzjxJ
ZI9bwfHE3+O31PChMw8PV8jQjp+Q17mOZvy9xnxjWeV6LeDCICXj7Wbft7MZc6Ao
7LHC+g+33VyNI1KLZDfA+GuXt9dj2tSwpugrzf7AvMNApOphWblofs0yplM17Xym
U4vHPJoacy2kIJUoVMeWiINzpahfj2h35s2jeCgVmL5r+6XSuSbo+YLBc+YCLY5m
uW7BuXtU/Ett+doVnXK93HuQ/TgkVRZwMaMLRWcfuGuGamWGqgpHXdHjaoB3BpJy
TA7sof8CRoDn9FkRrPp6mCgX6HWSnqWAzMVY2nDGNIDgU7yAdafUgQHKJ+ANS/2w
oa3LOTa0e7bc91lVRV7R7t4/DUm7a5mkjS7zIOxwt+289kYS53wN/3x0oMULW928
G/EOkpQ+dXd0RayUJwIjN6FJuv3TJKajZ9DtpM8f6Q1J2RZgVIq50VttrItTugpa
tvbohGtj7OUMutEmrxNhTZSgiBeW66g6h3kZyiOryF5uz8Cu2Ugo0sk0kcn/FI6D
ey/beI5Pe7c41RPSjuPigudOTcUpl7oIMs2j6wwNZyhC6G2eVsELQuCZjzCwGMkq
Vl+4lG9N9bOwW1JXNgzqR1eNugnhaLUWiAza5BEHoQt/De9kOSDDZyjhohv8cwUM
ShLYsBCO5YkMf4jG/zYSlpqqQMeRhmhb5znbPbzOvz312MvtFuY3SrcBRYyefCjy
FpmeO4sBsdpvQgyWwvkoArA6TxByfwpUPaVb+1iLvziPFPnsjKzgL5u+gKgfHhBZ
igTURrSjzKQz9n3c0yH3jAV1v7SIRylTzbLJWxxlIvsZw5WR3YTiS074f0pD13lY
W/8ThvpXkZxI3MkUSEeyWBD1w1ojBUBkxPPF/8UK0B5gDae6lIyZh4Qqxi6LfpHA
3Sx9RDGBxyc7yjemqAd38oh93uGiXZgEtvAXYoICr+TrsfZr2/oGVzwF9IjL+uRQ
dDardwcWy5vpBi9X+QdqFdrzhDNZfqZsAnhuImRQPoy7d/n9I3uWHYLbtU40FBoW
5lsCf9xLYFxyIvY7KPtpOBIxDl97t4wW5YJx3awh9Dz2ISScb3HMNznIaNC5HIz9
QoXIJSqCtEjsXakso/J8ZKeV5aGhyh/Fu8FdWJ2IhZ4iAfZ+APe8WpEBK0+Nz5tr
08LUYg8Oj8/58lSRw6/y/QAkVR8C+LZtPD6P9Hd8TDdfooklI06wUZ5pbBPpHrwR
wfbeWKY3ppQiQLatUsBcFJJ+X3cFE5HC/IYB5H77y60ue1EN/WdIfbb8s1+L059n
BR4lZHMIYu+Kv+hruViy7oQTeQ4b3RymBANKrlAPFwrfn9rGtMrqhParDnEFgRLp
bJE3NL7kXXIuPgeR39rDxz5lAKLW44g0O59cAQ1g/rkUIDeKdVSxO069AsusaizG
XeN6axymx2dEV0lLFD20RozdldNpAkTtNe2axWlyOyaJFw1BCXX730zCApS1Aw0G
AQnMOuH3xvpdJfOXTAAhtTLjGqYNcOh9kD+WV27WYn6livqsxG6Mugo+c12Bzm+O
xNZYCoPScbz3zv6LIKOc0WMDt4cHAM58kJB1O8u8HuOHBSsXL6tlQAliojFlKIo9
WlUbDnw3nO9We/PvavfppeHN3m+mWKsiyZsYEeWI/xCqQdAq/1TYltRQXxC6wcLd
B60LL+GWUgw6u8kGOvQckEDYl6SvYSIqak4f1AkaPqArQpk74uE8PnW+3FC49EBE
5AlgZb2m2t1+usJohmFlnDRhlUxA/vaIsDwVbOsQZxxNyLIlqM7F7UU3pcTVMYNL
K23NhKL+3S47p4XcMx9Qb0itl2ZSXrEesdIg6oUPKI4CrR6+pKrNHfdM4R8O4hxZ
Z1zwPZSpii2e7Cx/Jhm7FWuTwg8/oP9KdkjIGQdCzzKIx9fZY0L1c073Bl1Od4yP
uyq62BsT51/ae9F1R5hEEz1CWDOQtY+w+VPehfB17ksqXW9MOxKWVYOE7RmomUVn
Lzslej4S33VYy9oSLj7jLF1zgkNWf+PBilGGnJUF84vc9f6a5ar4g2TmRzel/RpL
IGMQhiW4Eztq3tDV81iiB84SKOSH4IdfPNWNA/2A1oic727Nsgi+uH6ERmU95fv4
KmbOM/nOgzAxCU0VSaMWSBfUOwoysm5hunsv2HSNM/Kh+sRENOqRvo6+HKghOdSr
4UV7Y4wbWB+fS7tLpButnDeRhvRsQHsRGKho97UnQ0umjatnFSdxfoU6Ev6Dy3+b
hiSsr73qJp8/yz25nocdNxOJoIoCPXMeCHDCaKP9ZmZJsCXgXcIhCytKgFG7QYCe
bY7wImTjYTFSzmBBtwA607Ehi9FViAxvForoypb2LKkSXe8bPL/GlgjSljwyTm3M
e+uKV9lRFTMP6qJwYg7TGY8kHIsV44phmP4iml031zh9VMD4Rtz+HdSqI5BzXxhT
rBhxvrxt/Xedr4IHcP04sw/WzOSZNkqn5V4IFakc2QllsXQt0THgXUWjrWPcYs9i
0VALgZN4HskwuPSeobUPoFOYHOX3q9L7rSKf0wKiCK2pVxbg0LjkbY3SpnLd4XRH
iAF7ubf/BekQtplCwIP/8t7g3Ol7yLns2tBVO+A2duWOOlHW7fPnUcBKY2uYPGs3
ps+k7GMT15q56WVCiJ2MKtA8wMbYhgN3IWWEEE2J/ottx1O2p5aWaVxmrk9Do2e/
V2/Yeh66fFPgs/y8a18JYDzwrbZuJKP+C6fsVIgKcjz5/8FfIhYxzZAAOYZxN583
lzAg3A99ozBT1pT6b9MqF2SHLmiDBZzl4ak6H2Vs/MZ47NWj+U6CiMkGyHdy4aLT
CBEvDvZl0eITwYVxhMCyAbRVEwYdBRMCYvnI4xNFrxzeHKQxtSQXxm3dM8fV8oiI
XNfudhlP1kSs2VtoXg2zOE76FOh3TcVTMe0jHWXX39JaBFWltu2wykFlga6CXSk+
K1C+VPqtY3p0KkZ4Y7PL6fdHGZiOTVXfnryOdeDfF6oSGHE/g4CywsoePxkpmqht
Pv43iJKdcCkY7eUMU5Llu64lk/hQazozvuRc1ldNs6whGVOPXO0fuoHkRmCEc8Wf
3FYVON6f92pI/GNlSCaFtPw53wPxp3SPRa1YlJ9VVcY9B4CgD/Me6FQOy97Sj9/M
mtO6W1kbAmT1bmG5P6dn19+FMqKkmk2bTJFo/nYgtR5qvEqczeVzpVAD4JIFh+5q
urco5vo+0e8MoYqViPcXQRWBZaPpOGjFKcypOINoFYoeiKnM2T6/XN3wVSIUnQRx
lqvlch95rF2dWac2RsAGIZSZIvoxQ4bDoHFlhyQI6uITW4WdqAFWOX9FXFAH/cOA
XHGX4+3FiZuVPAvuwoLRgNGoVbMIXZqW2WgbqFzyyhdT3WdPcfEnavvumCSIpbes
aQHA3a54B5hERP+v6GYjr8HHlJT+DBqc3GPRCQtB7ESNq6ufmqklExJuaX13Wx2K
9HtTC5ghRIiirJ5SvkiqE6CUK1CW3098oyZEeXCrystjTGdwjbo7pvXeYDZ+L4qI
krSSINTMMjItdDDjdxGGBffStndVVwSjyZO4d3JhbwHE6Mr3mJuiKJxTikPqzAs/
OP4WwQGdTZGxAbTeWcnLuaEu3KQbjcIKojzeDbY99zkfUjd8X2KgjuYagOUiRj+n
4YY/e2ksSOWddad9h4FA+hvClSruGUWg3uZDE6T+1MSCHFJ8z3vKtQOH+2W0oLzJ
CsRtgWwXIU3IL9lZqGRgmNgjNZmTr2+nrm4p7Ash99eg7qyBtbbBDlDaYuE7FyYL
55YbCTZ1eWl7viDOOEvBsj+iLST5ll6a5G/AZ9HeYq/WbAf1wY8XVY9ObWMj36Du
R7FN8UsVyOqQJ9I1W0VV0RFaXGj/WDrI2beXHeVyEP5QiQQsPuo3WZO1WiX+muKR
DzFsD7HYCTCBgvXYslurLW86/QZw3ZJztVjHeKTEleVLOeF/2sozqeBfvd7gXxZi
FhOsBMlwbDGs3qxsku2qPGUhONuQQx2lXGz/1uoLlhNLMlGRJEtIUtqG86xSWOAJ
up64itdOCdU3yN4B7iYMwE1FfLeU/+ygEGeAfqRpfhMbqBK9hnmUjHun6m2cq6Rx
L3nLpJx+U/IPIyWjUTjBdnW2gJqKl8wXG6WiPaMc5D+/gq1M1JgOtXGnAWukSLlH
V7D8k/wAjlqdj/PiWG08Z4XTVg6M3UJpM58Ru7JkcAatoCXOKmcXnfxbP3YX0dDV
q9IQtE4Ou4YsAlGWGbjrG7OH2PFdEiTHPSOl4sIzooomOu7en/ok4Fe0NWNiLrM5
USGi4mNx7pUQUCA7+gL8mM+JBlSHk663mg+EeFb/6XgZmQREDfUJ4EiVTU6l43jp
vpCtgCuRRm4edUBl2MwWW27sNG1eSOWcXDAlN0eKCJoEwqt8uoxjX2FX0peoe24E
Oko/AIQrZbDsW2mQp16ctqWDgjXfqoDo2Be1S3X4Tekmm1eIVndaVloNpELePjSp
Vhfr5qszSzXEbGhFu8juGoK39dUVheHA0S0gSVj7aKLhdQmp/3QQUNVPUv2QSjFM
w1KlDST2c3TwrZspRFz9OSqVoVqbEECtEnsaM8KtvTdg6bamjN0KpJUXGCoCsq3P
Qop+6b3fE5B//poAstSem6OPXfIs3Bjz+3w3DuY2uLYjzFILLQJ/VVz5fnebDjuJ
g3gumOthbOLpQUVnBWXZHdWNvRSVS4uh7YXgyod+6iJ+6p9L/FsPwWFMWXdBPwjs
SB2wNfoU0NnU5F700rRgk3Mchgrw14jvvKn2FPzuS5akZL0qOdiN6DeDtnr35s4n
B4Sbsrex9b668Vklv/jE9Y8ee+DzN+eRuftg6c33kxkfwrb1cQyy5hJRXgG9v3D+
PDLI1xalaLG1Z60j11vCCp4zPrGpGQPr8RE2DQLBHXGoYfrkG0jb+jNQIvBvPLRl
vF29zLIZlelM5+qjWaJnuh1/WtM1X/CsUXuBC/iSFTkaG/WajukdjOaPSuy3oKtA
td1pyf1pP83eMZQV0iQdBU0eqx7oY4KMRChUIiwfQ7mp6KJoLW3Q3MVsHp0z+XyJ
QmRizvDZNNKKbqH8iLQomLtqLLNbU4uOUUKMpEPo9JPWYNa9hdZVP9i9BSxQ5NgU
R8S5Frqb1qplA7kGAMysHNCF98AUEpeSUPkwn78dVqMboL7xdiK9ANzmPMBUk/6q
K3gI7DxS2JfyasZ36mCm1aYM6FuAnb9Hy4AYZKoeSeo93E+cOLijuPPMkLZ2Vac8
tgQ+hCCMe0y3PmGj+ZC63Rv/bnL1k1+5Vo4eDmFSUzq5Hs5e4tqfrgt5NPQ1CCI2
MISfsod5LMod3UcN1avTpl05qvVO/iE7XyzWLoPKAwyVJdIR2o7utFpM8TpQU00U
jtmgYrgEa+PqNVOX+/tvMOujrSY4LJwBoS9InVuLu2n2W6vH4Mozkmm0SHrINRiJ
LyV3uD1XnMoC5XxDaWh4tFspfMUKKlmluH81NwrZVSzWu3Gp/32uCD/55to4WtrN
oqH184T9dgNd2mh2Yr1+tSh7Swl0oFWYzpf68+gXjv7cpc9FWqvFBV5PL8YdIS8z
1HynYJ5QvILRs2ntxCGDAT5YMzMHBf5oFcsD/AUCDNOmIw+mXNgGEZgs6SRh+9bk
52YYP2cOqAMcB5Rmb4RkqTifaAq+HoQ574O5Xv8tijmTibwXJZEDIZMkUkigyJLU
T3eatO65VotALv5g34S2IxDRyAPKYCLBM/q6nixA30+xkkXtZAlH899wo0tkdeyc
vA26KHbfZ8A6RFkKhUZe5AtTlhO5REfwz61TQ8U5FD6KLWZOSG9Xtjo0FxR3+qbG
cmXYdnoxSldXSIfBN2XZo+nHvNPBWIATsk5Qe7/9j5UGmxXDciX521HQT4I2r4tC
MF6Q3mPGBv/SCVbmqZR3blBNdNErDuF4LCBL5kGLmkoxdSSYL2zV5Ccjt9NR+rGI
Elu6dlcIDe89yp0QmH6h5ktroUhV5GUUepeBoVR3OklN52jeX6U1CDi2JUVC02N0
XIb8inznV38kbD/pjNYpPtX6nE7eYz88tV/JEUJyNjjF9bJGMEOc5+y36hwPVcJF
opharycbhbuADU3hH7YuaxqhF/gctrQ7Rk432L0YJxckc4T8Jcz4J4k+nM9Mrn31
ywmKlCyziUg/7kgKExJQLYE46SgisiHMSyPWgFGDVNbT9AW04t8TV1yLDzR3pvMk
uquZF11PARmYT2JPgmdzoI2j1AWYxoQNDpKrvNV9xshpz9nelXkYb63JgSorP06a
2LRtAAx11fkozQYpdk3vpSIdWc6wKJ4PXbQVYH9CuJg44utQiUAx5OHyQmJx0V8w
iY0GAa+sF/7KmSEYPZi3LYJQ6VQuGFpe8Tapl5p6bBZqy9a9KYVi+dPYWJysTv6o
EKtu1GbOKIIvQ+h8upYfOsvr4I6fNsJcy0SJQByQz+7l30EiJf+HIObRGHc2AICq
oMFrltm6QzpvtS0g/g7V034v0p54TXBDPs4WIrsiXQImlw9RJDDBno9GaOEHVM0m
oHqcvxIWK4E8hQPE/eD8uEphYjKnUQkcH7kBy87shVC3cdTTblm44bmWARq8XFTy
ZscoV7Cik1pbDLg8OBSdnxE4UTvrQRntVPARcrwvGktZXELzFGPtodILyiRxD5D/
6RzVzk5YNTOa/68br1lP2lc2494eugcwGADSuHNLAjzUel7+s9gt6R/oPsYCS5iB
hK2QGNIcAQ39TLXdmoS+gQBMeAP+7Id2wvfRZekS5S4mr6hmjcqD/mVFpXXII1vj
DQ6K31b3f1C8NSOh7m7a2wG//09Jfx715uCY4MXDIKz5bRw1iOoKxAi/XJT0K75e
65PHBgOBEhK4dycA+40o6qUqpAczaNvmCE6scBO+sZ1umTp0Mdr4osnX2S2gGlWc
BZk9RX+A8PEt7nOZRzgu7t9uHZ4Fw3GzSS2uKi3SudlUbGIutKNa8ZXKC5Kq4N+z
ajNAkiPhx4Jh+ngl+Mod0YTeKHTCb8GThbh+zHCcdt6gVIKV5ElqokdLsMZgOy8C
/O4wTWpUqQ46hQ2fxhfRnPOqvWPt2HsoBHdQbzioNKjEb30CS3zcvKfEVfT7dMlf
dR75BLHEeVlQTiQgnWDEgX2+dXUKyByiVCAOqoszxV+QRickdR4KMxBFEzJuwED+
eZEb+j+H2oQN1lvDkuQIsuDsfuNOVEaf/mxO3zbbF42qYLB62aAoUfJrNmYKxeXA
EDBDuC2g5eqMdET+M0ov8CvinnaP2dTcKe88zLu0AW1FSHmL6G3NaoXrR6xSIB9Z
lH5trkhLi4maPDslTeVNhAVy8ov8gN/ooRP8SO/LvmA5jD5psZLYTnlVvcb1zibP
XjFdb96tnZshphsCnXQyfElaPbqYRpxGPPC6FGLCtSSWKVLAKNRI9mIuJWFeY80W
5OR7cHDtuw7DPhuLvNga7z4q5QjGd+9Dd8VvtEGaN6g8lw01ooi5bC5sllxx112w
9hZ3ciBMF8dsoJv9g0VnaW8zpu3mOzs8eBMnJz1/QB1jt3lzIGoC0okYt63ZlCQz
RWINkoPY7udoBUynFUYT9I1A/1D0P0lH9prJefkhJmp64Zx+XPXkSXlc1AlaUArQ
bj5/JcXpBX2sBsYCYsh1dvRV0wyVthIrkD6t5332Ol6LdoJqZWFKr8lUFiBvf2Wc
hOmHUDBQ3mEaHcYXByC7mq/E6HUCVbCfIPxBgVYO+5Tpwta5WiKLVjH9c7uY61of
9x7FnrQMRYYEb4fbrKuA24fBSJfVBV6PTspoc8waV5k0WEy1iqMfGXujUub6C8ne
XtnoRuf2gMhqFMAQdrRtBzp7n1JW+aEY648YN4DrdavvoHwmEmafwPNZibng1Qtd
/5Geoj0jETN5VBVL2/LLCaJIUMOVVYlNzbG7304l6VqBkiwb7s+/V1G32aoq1GXO
aBehi3Ei8QgCeRzlrOtLnvwXGTAhnqDmfzy++j2Vn988uy+Bp4uku8PVnqpxSQRf
6U0MDaWL5uXInBjZ5rKglRAGG2TF6Y+SgoLk4EeN6ZPeAH4KRzR8nURyLnagT05p
3eu0Ka+QjIIbSKonNJd4pDfjq20aqFAiKZwW1T7j9lNenbmYRTiuMGbsNdH+uVzy
7nHyzXJBW7fN07yUvqXZ7tL8U4DlceJVuD2zMbB/lzFX+bg5uydpGQ/T3QfQxACs
qf3xjjw114OQTKjI7OAZlRwEaH4UEFOtnzv6yvb1mT+58tIBHQzOmPCNOiXJdaJ9
ZVpkWe9Un9+NU4PHr8HoV8m+HhwdViTpAiq6cB8WkoTPBlaJICpFATUdvcmIGDFX
xvUt4rduG5QXLwMTW6cYAEHBCfRi2WiQReEB3BNEyiT83O6tjC9TtBmQ5Vg4lURj
E0FwUAPJj4peaBBjNmwpCpYmXH4pVOPtZtljPM3Zi+3KprCiGlUMKTzRCLKUgv7C
qd/oHLHjaOSPPsFYz3hLSpKL+2aVTO1LRwDDXzh75yif1CBNPqRxszbMDk/WOkLi
AXUMOg4AC03T+vG+FWD4YMn32cjCRO2/lvcfDQHN3gyQVL7m2YJL/1o4BCMebxkA
nNAxnTT4m2/K2xsE7lbsqE6pUSJflwAeff+9D2wJ+degmpRvrFJE4dCVC/iBXBLS
aax7nFRCVRepVIPB2ivvrqwHaJc8rlERzUiJXfOJE79xDzKsdglqGntENsTCzLxY
S70kygwLOZrdjJOc0kN0uC9lUW0uNq9zQKiXeFbmTwOW77cNdvgtAru0xmGrUswW
rQX4i3cSxVJo5Sa0ejr6HtsYSd09hEAu1iJZ3Egx4wLXl6kjawvL3ZP90daU6zXO
rdOmbBP1uYvY6BhaAQTdqyrQGz7YOQ8cK8YpzJiLNgOBPCz+pSj786TMN2PGbVU6
KzI7YZ4OjaZ9zQKd6ePIjr2iiM9Csqk4l26T9ugysBvixPZm0r6HSHCs0CzT/fXV
tUaNSgAIQIuNKzzD2bf1VF7oFjdXAW+aHrbNd/brfoaTWf74hN8Rv6EAfEeYxVrB
ztldGHRjuw7LFuB4V6GvLZ1cecFgPwirG8gO3rLGbr1oO0X+A2dHbX0/QG1f4orS
YOjrrKCaP8J8xVGdf8D8JD4AnwlPh1hRNK9hVVbaLa2UcnWwXfAwKXG5OYJm/2JQ
ynMfWJJRX8cVWghTVZlvT8aDCUudrn+WDR/8fk+NywbM1nZJsLVv1KfdLHCSO9u2
NillP5y9XOURPgAb8ujwyYx88Z7F7jnO3I8GLpxRZIeqI7oc0JiBkCRd44HBQfnO
yc8SieK0QyodvjfIJeyHMyP43rbmiNEA197/dh9JpzFjILaYV2fuLzniKiovzAYe
DRo5Rv3PcUc9+y7vgcu5w73uvQ0dnthisGmzLZyWLFPNf1Tawn5PGlDeJ9ra/86n
AkMrlZM4EUmKljqXDwo+fkP+uMSBsQwko6DGqugE3ggVt7nvv98Q6r7gKIFfEq8m
QKuK04etN//vsB2cdupSDtm+dHzB2FlzLCjRtdOg0FV8mMn8yA6DVv7H2e1dDyEY
ofr/It6ftfdNIOMosbX5JJA9DaGZOEV0InAMHU+CbzymPbZ6ZF8H4hCMiWQU944M
4HRMF5hKuEGrxGNB6zpJW+YNn332B0Xz/DZq16HbstXugiu6Y4rSWdvkx1rzSkYf
rK+pdzFAoNKtrZ41jOnZpI9yHW3DzMoB7qqT+8sGz+wY8aPfs3cyxkw/7kP9e6hQ
TvAlj4aonAkbGYS03ooWHQ7J8jLMRffB9beJm7jCRRQ7igehCaFBnJ3YN+iKZlym
oKYSM0IS6wFaJ1xbkEjIVEtLSzCfu9AmXNvFmgLeTQ8MwZcuusHzrAJ2DDGxV3gu
15R60gJKiGWaFrRcDALpoXRf1uqFAeGu+7SE7aTIDoq3brAuv0C3NnqyBdPnsRd5
DoyxMiTp7pr/RFZdGvhde6bg5YG11OwkKBWrgUNZzTnIGx8Q17WZRaxK3g6IeBrL
V5nRrIG0OZdE1mzai97C+yOfCKI+Em8rX7RX784g7LhD/PhC7KWnyUxA9+rJDz+x
kLfQwrcrpyGIlb62i/Au6cgmVG1NCIXzdUWUZLOqFXmYY376P0blsFI58vWeLX4m
PwhmMnmHOvnFnux50nQsW/pDig8fjEAFo8odZMMYJ57e/EtVgfRXjP+J977OIgb7
kQ8dEEYSP7AIjw1h9dMQ6mlhkLF1RIDSt1nHW4rh5LV0YrGgetULjdSEZ7MPR+Id
hE0nyOyxscuoOafexNnaFyMbeVkR4YMT/m5i/v4122itKNEc6Pc7pvlpD5yLCm6g
v0ysdLAYkMBPxNvULH6tCCJeeDsXxPiwABcubaFPGHfsQrtOZwG0jand931Z6iHV
umgJDx2dw1BcdgzpLcMmqj1jZvq5oop8NvfhhOlbl9o80q9Pi3d7VnkZ/qmRHV6c
tenT2wD88sxkdYHXMz7oTxygAn9X3XyEI+OucpoWJvPkBlrwGjxBQf2hUPDOBV7s
1L9VLUl/BX3gNqI6nXx6NosgVwuHnyFIFNr51EVEcfOg6t0UkdehD05arVB9gYet
LVU1bugy7GDDT+IVfWEHlvF2Xw8XBzPr7qgUcz4ifDHf5RtWsjhTss9LHeFlhVMq
z+K1ClP7Jn6Aa+0owhsfraSRBrmpZ7niyKr8qKbsEZqpGfArbka76shPfYZafC6D
4DUAqeEHhkjXPSo/i8yiQ32RcYpfKhFDTflBCZxT5zoEhyQJJME4poQHXnueXM/c
0HcnL7aU3q6zjW3+ylbmpMSdFtQ/KFQFzNoApQvU7zIyOv4J8UNujXnJhnUU3DnR
f9Q7DRAHUdD2hqtSKZz3n7//GjWzUzCoMCMWS+aHceB5hh/vxtOGeWyvKR/Xltq6
BgEpOQisID9Kt1/j2u+EcKgl8znoYMSr0/XqjfugBJ1oYOrUwY59/hRGQ2emyqOa
44t2OsZfpP48HJoI3ieVlZCXigB3rESg19d+jMiFmELR2CIAc57blopuVQUr9CpG
MrS/CX3XrI/lXsMhDt8fozlSv5Ah97L4XGiiuEUCCP24rx5YMmFtUD2eLhtGVtM5
HrXuvnUr17vhUaLQYZxuMP65QrETS9ooyTVXHNWzIgUg7bNMQDyQ2EgydeyJVUEy
lVxHJ4UmThYlh8P1Nyq4ZDUO/qMXX4RqIbDsJGEV6PIp88Zagi6Rlv41F/abSSdx
8Hie46DsZ0tWmnL3VgSAg9sahkunbA2TdWuTUg/lg5v5bsyYXTOMqEkf6KL1FXGn
VCc6pgsSzm4lBE5auqEigx4apXusVRJUv+bfX6U6l+Kg7yOZep0orWpu3CkDEsfn
aAhpSp+X5KQ60y2ru+o5R1zCc6oDLYpXnr3QrNgCZMIU66ZdmaMjeqEwgpUFRzGz
XPqdTFHYrILkRgH34DlmGHEuIaP1GPHxkD4szVBB7WbtKgVyg+weTbHMfpxkJUPH
yoxuU4alJAEGM20fBUM77tzUjdreDg5JflL5U6SI9O9e8G48SnODoHyhdyxZ5MmM
QR1SztUGXVFD2su5BzkWeNjTNR+w93g7mvcUE9G/o0JtqbJiRMyGYfV2Qrvdm9ij
VClzZDOH+Bd7f0YQL/PNhQp9INn0RqI/FLw6MCe4XUCI/u2DvsnKm9OUbp96h9c/
xl/F/TzQS+4XX09aamHmaJu5KC6xqx1vFHmXwveuMcm/4sLwEBOusVpRUBoYJH+U
nTF0RQc9fvsBoghohQ+c+2ZVNtE96WM6Eg7NdPD5z9YqWSZbp7k93FaeqtjrOUCy
GC03yyE7Co1foe/26ulv1oNDhyYv+ho6aKdgFP8CnL7tv+sH3b4RiJFBOw7qR3qn
fX11zdLq2wxi8sK8oJ44w02IhyFwZHgePCJ0Iw2MJI1kwHzQfRHojQiWDONXHd8a
F1hHHcoVxVqyxsc1EWIt9J/zPthALIqW5NkPvqfUjpP2u8Qvrwvrz5xsc2qOAoRe
LCxzHyWSyRDBliWIk8rUHHsmRqo1moIJkMgfJ2n1ZZrYwC9dI3LRq1DOWC3bq6pu
0OeJKFCjHafFjmKd+/u0k0WqS/vu/ZXvw2DHgB3uuS/eXDSNbYV0sfRfIBfzrndV
Rez5D0kFlGh/JUnEPiEiaG/etzRFXlL+K700lq4jas0DtW1uHQgeSrNbBLulKAyy
lzDYUmohwy6WRtOs3yyoCj9J1IKEPqmXY9+px7zPriAAUUQV0FkjnrFLNZKDrUZb
8QoInPd0wTGt4E/EHkZJKTLToKUvj+BiJU8FVKZDhUdcMobek3fmHSWOCckovyYb
tRuG64afD/OkbPBvxMYj1lXK5ufpHeoxWwVAdFJYuF9xVO4vZcD9RcGM+E3zYYr1
r9edr6Z/em56+5lcPtw9CvT7JC5geX/u5YD9bAdd3QvnG0TCO0iDe2RvLGgLlBKt
4MxAb5zif32k9J2RD61F8PJpbAuouy4rTjmIbRi9hFq4joU3hnqHSo6Fe7s8y3QF
fYzLTL/r9+K79Vm3h/uOtFO6lzXJG34naSPvUAf6gTVgP+kRFEYZy0yGPF3UpzsI
XBRvKgt7rP6AsdOmmS6nxN9VzS1Tb7saJ99ZxWot0bB7qx6SB+j4ctQ0gFlFmUMa
4HFuXzpup1wR7x5RH5nyJV/G5ATCHOEJjc5BffNY2xkM6TQ8+jdJhMvw/COJ3zZ6
4I0Yh4uKemMAvyk2PyFBO4nl4Cx2qoaKuH4Do2S9Cb+lY0K2DV0e5QlORki1yE28
VwvlkTMcbgCDCiNM1aiGwDSXB59F4acFUsOJ4E2I3FLG0sqfM/W9pGb8DykBJWcR
yedv26vG8Qc7r14WO1rYzcJlJmy3bMSEbJEmBB/A4IzG2bmtdB5rPdfTIY47mBm7
YaNRFUj0fJ3rk9nDRwuFwIMLY0/rvSW1HBYLtbvJD+WNS3cKThvnPigrpiJ3pBuE
/IeDMO+nD0Bh1vtmxo7HYTJ7PLLa7X60valSbheZj04y9XhShrHGuwvUpccJQW3w
ef1vYSCvxPH62qzbA4umjK6Yg4gCOeXhk3cRLvJvRbyshipOZ+IAG++/v7siITXX
D4E+EsSXSBye4+g3cfoIjz4ObV77D8zz+4aikhYieroA0ZaUD1mO2CqwB+yWHCku
kBj549ifq8A5kp1uhQfP1EXZa4XW72v5mi8VA2LB4UH+X30YGdUr4U5kueQFYrWT
WlrR28nUoUMGYEKOMtwJV24hOwAQvGzx/orGGEL6SMYjPyhMcuUGHnmuRcrtcNLp
pLZoJnmpSo41J9XUt4JQ9DPO9VVDLM9ousOqTOrEuz5w0jCPNVXrcssBeOLBmyA2
qB9py/WVxyVvBceQCbMtUwBzF8J9s8ltPiW7y8EWLULU3Y4T1OYMhKGvOOPqNx4o
6NBxjnhgJPxzT+SfkEwXjbIk2AdSczhADmu6YtKl/GtjT+ieVYk4OXUiVEFxECqN
CJbZhdVQyAyT9wODPStIGp1MsZcmn2dxO5SWVC5d5cMuIoxqQfSgzNRXLJZhEstq
P5gHIoxhSbF7qAdwB/6WSHcDNdRVOtR/xyqr4DVg7sWm2VA5lUZzD8kKC2o1PK8g
vkjcezfb6ZVTu1NT62rfNRFVgq3m/yGpiOAmd0rOy3sXVuwGlM6fjt1TTnzKSMzo
jmvYPmFdue4vvkuOKuPtHajSoV5bGlLzioidvdBT5Mu1AJlz/LQCxgvd9b45PIbd
uE6IUKMh+HzAOYHQGWi8+32cGOLVmEeW5zqX3lUdqXeZsDRCHwHkehYvGn8o7QkH
KvJIUGZbmT7pEy5wDFo/4QUQYQgYh6WRr7Q1AVfHqC+XPI38nHjaPxskoQTkIG8z
kPgqFH7e58EATAGXFR+xvFgzCzN8M7N9eRW/EP7455G3pzdVTU834b27uGFeaf7M
3O6FALdffwt91e9OYcyqU2wS9OVndJzUiyCAxvExRYMPrx9xQnoqJAbureKdRXIo
4IZUdmdomHfBOcsZXysr/xKQxs4xJsgNacyobDYpR97LJiONldHQfxD3YgGpd7+O
43w9XalbJxeamB6o9zqDeYBnq7TCMp8mrWtI4q1K/dtE3pnj1sVw+HuqRBhbDdXi
txZtmDODAaFHXcgo6hD31BUPlynIMcs/AYk3XRFlH36+aY58pbfywK0pOPagAywB
iZQDSWjr/TOQXb/wjupZdTZyBpx0DtCFm9IQPxGZXuNk8rqp2Jb9V1e/g+POjpfZ
CzUh2+SAB6KUkwXzHwJjJEzzcBW3iVrqfVC1KZOV7C5EZqR3Xqg2xcxIKSuGwGaG
nsepHKVegeh01Ydx9CTOK1OQ0SscMeqRDcuiEJAp8BJtMBijhljRuxrW3cS949iF
L+WPiaDhujQ1QYSHif7LMGteqm1qgcoYVMITIK5BzGaBTSB50oZYQU+9hiDy+q1E
nHV8Y9evjzMJZMMw49z37I7TY6WNK4MZ+YgTBdcX8uhxff2VbkG4UskDbKLB0opu
JNkSatKtwzB4rY4OavZrAGrnPqvpdL/7sPbg5P3ESktGhMqmo5O9Hc1WxsoDMbvP
F+MCgF07L+GF37LitrqrsjuSqu60X5eDGUNZvMsrhO7dwnOYSbi5ijVT64bDLXm7
mfecwkCIjtadDF1AoqJ+Tm3qS3kBmGdhv9nfog8pdcE/Rt1QCuSmQONCnTdsiX9x
zK2CT3FgUu05Ba6bkIU5zSRYa0yg0fN45oDum5Stm2VGQH163XKR1cjf4vjQJ4AB
s99xOCaYhb/m4SpzAWbk3t3BmMmRm2cKipljpJOhxm6y8NAr/GksB4BQ9UgQTg/p
UOl8tLIahcZZQmbUXi3N6rErSMBQzXDdfPFHzBB0aOr8EQMpA1tZjrBwjUp156XN
5ui6u15CGULicMtrKUWSVAM2etFeUPS6KbQlq8g92jzccJdVja+zpnbcI7Ndcffc
7A2cQoMhKeC10YcDzTllKfJe5x6kkAIiEXk4yVMxvIN3vtrG/I7s3VW75l3O+v/Y
gmznDTZaRsCdAkf4opD+vdCd5tHaDeE/99FwTFHVrxHRuR+ev1uJ3ba6wjCuLOz1
h2DGNmllTd9mNTiWM66Ajj78lAmMjY+gtJXQ/+DTS0U4kSrOcDr25cL1upOgjwT/
IrlH1w+Z03zl+WN09ygfBGknUyoRuV2pJwfXSwl6DAVuMKscpwPGAvjGSA6YrmyE
PElNdhe8cmpu9VxRW0tKwOAEPofzsSGEfb6aV8FOSLiZKWqw7Ux8VDO37tc3ppwu
yPueBffNbvufzs0k4RabRHFU+wQ351i8Psje7rS2LWWd4hViYoXgKHXPVoJDjET9
VFCkseu0Cb/Bha7VHx6MRH3x/NvVU7v/B4DuKp9W+3HPUog2rLUfb2v42Ij4EtJM
tlXKKOL/FCd808H+vegT231+JoUbZh3hIHxPpI67Q2G29p5Tflr4MolnlGfS4s+B
j9rpPpJ+p0fvDTs+wnCNl7Phg3Xk69IgyN5kqjf/4w5Z8WS2fQDYh80K1s/CqbHR
vMZXeEWm3U66bNbcd7u6FL4p+8Ep4GoczlUUx+JkmqsQuIwlliHwB2VJEBF36GgJ
ukl+WWsJnPSsKaW7DlNu4S2yme0dQjRwe6cIboWylXQO9Uli0TkZOaUEnH8YpAjn
MQ8/dRQ+Yx2MSBMLGO18TRjouqG8ZvKqaJw8PppcT54vEoB4g8G0lp1FW6J9qi5C
9eWyflGREWvJo/DNVBxgS3KrBFK8pYbWxEvIApExrMubYbmjjoZ1M0RbgQT5hctt
V8kRI7SOwFfQxOiLCexbkw4kmUwFI7A63Wutyce31CkXyA9Gy9TR7dL1WRseC0aT
sGJ+iskLDGPwJtm8pgHooDM9nDlWV2aCnyvK7A2PjteoXDkyP3GM9I8+FSSlN+n7
A1QAFR2vMuE3r3WDuLnCB0UTjEE9jJL1Zq04Xx0t50BlXQKnFRsKIOwT4bGRJ1n4
N0TuwQiK/7Uw2gHbwhiYK+aOi+dMtaftbL/Q15esJ/LpKTP803kp1dAbfckDBhFa
PYEsTc8LhAH4+eBjTfjdWjs40A5cm5v5nY+oAZ1ZFa5n4JcIHgErS+QIjYejvaud
9RFNljMWxqOnwEcBAzc/GoKgxWje9CEOeRzzIp5ShgQumxbz8RDvuCMl3PswkU9R
p/1+b7OelNWTWQMlG/FaRTOTfnRgZoMoLIzAsELcg9xddEWJcJD/mx1RNLGuF5XZ
6SWrzupZ9IrIgmISOiflgaX9AaVP7bPORQVMMbgNgjdeQ6WNwiHwrENwasjYWI91
0kBKDrdnCfsUPD+1Yrrz4sQGZIgqWoD5ll3bHRZ9dyTTqFHooUvMx35uBTDtE1T2
cXwJGyGANr4X44bQEKW7SG5ki+igC+JMS8wjqPCttjQGr854Uk0tUw/AFO2oMw/n
4h3q9WO7LcXxkPPFZUuWXu5KaeSbCU4Wv49vE1SLZoju0/ar1B3itRB/8gEQX4lc
t/cwfmx88wf+yCMJWdlQWs5pUOFoCHJvtA/fnpP4zaUDibSstJHbc2MusYt+/MTk
5tQTBXC3ylOA9MfoRR43eFpNv18FlLOs8raZY1VBd6TwFPviCliKwydFQK0/adH/
kN0pr4/Jgkc2ha379xBBxHz0DWPYfjCYl5l3c2Kulh1tDNgeBO9zdTwmtwAb+ZZa
yEWvU3f90uw7LJqWb+hpQOnxmfE0Ic2+mjWQw+Fy7tUS9mujuhj59SWYtwGxvyiJ
/8cLlQDxL7i3gS3QPZUkMtIXQ5iUQGKayn8WkXVMrDzZ03DahbynreTzmMn0tcLY
857WwX1CyO2k8pnvU6fj9V2RqtTCxI5+88wWuDMH8O1SeoAwF0ItQj1fkEXTtyNN
/b0ERX/NTUh1AvCpZpbIxmVhbdZof/EnjjIi3ozRgcKTFESn33CcWwsA2MHv8dRh
IAs1DG61muFwnKvFN8aAEVYa8DRdMV0JNIjJD/2WagmvWecCj1tYL+QZKMkPdQV0
IqFD5Uku72SzVfpQcm7/cx18YuB2h7ODKWLH5Jk12cn6vmceM8plRz/ZBUuGaBkH
WrOLeFmE80nLNi4eVp4PH0Xh2R124qZp+BoEl5c9b7jEFtBAPKLtP1rYiVjynhzQ
ziHRhCKnym5oSJsiW8fdxtXjkylILDsZTl1t/HgylrS5s2eMxoET0eqIn6xxfwjH
wsIQX0kSFHzVyRn+S/z7Y8cuDlL7S2Modt67v2javv42hy/zrGWZxlUMIBdfsJgr
lTjZTn0uax6DXTIQNKrsAQzeyyd8jvbHPp2pBnEIhboXh17j2xDXlYKTMulXaV75
WT8wj+ota5axk/pkap9D7gDoFKGddDfqkzRUazdT+36jui9iF0rQHF3BWSFtXEbN
DzuJcfZQhe2OVDmiC55XXf+B89tJWu/jJhOkRaYfzyQDXtMcWQHCdfQJ5vQ65WLF
xriWgcqR9L+uuOFgFCfYkFAxgMVdPiDxrog7aElO2ZaYlrpNLeZpWYlyFApS9f1w
mAP7LaSYAT4M42LxJS3WcHlSkTEmlJLlQHol/x/+DVLuqxw0lM2isTI+ONOObSRh
/7IoI/xwaqRr5rhTieJe0w9fkE4nVniaKjBaA0EXTRn+ZfO7Pd7AZv07KJiZUlbi
oyGPsC2Nq3GZSsJYHCVfSjWxppqitfhFrNDAW8uuJzhZ7R1Cqk7QuGLSxQVk3Kya
B1uCtq9X8W62XVjEOYUCDQvGj+XNiHtBNFJ19NOHwIxK3qv0b/ytzstfn2D/VIb0
lIlV3n3/9g+YVrNX4rrOQBBy1mDKPfFExJZWNpFgM42of8sE5pRdxxhS/IHXOpCG
+lAvitBqrW7b1y06iozGdgd1FyTt8S2Jfp1oju9A3ZUamNPxdqL98Tbj1svNs+bB
7Pc8qorjnhlW/a0wa6Egk82ZtDk27trqh1pp6K2pfCSGtNDdiWsnf8yCGG0fpAbV
G1fFCJcM/AiWQkUPBr4Whi+o0stU93p6660CmXF9NJ5k4KfTKo5Sh6C6farQPz23
Cb/J0+8dczBpQ2sOR2IP1RPvB2sn+lJt8htY0dnZK9AYwKynzlY9tK5mXcVPGJDx
hwkn+bog2DfYC3vv3CepvOooUxFW33VJPtXIWTPt5A52bHfkb5AoFkbiXuxY8jqW
3Cb4ZiSOwCkY0Hz5Z0No5UdEU9l2JPaeYFQrnc7gLKmqe6lTfRLFvcCmwQDS2OLn
E0ueWCwW8BZ82b9ECwWmKNk/2iStZxhTTIzoC76gAYvRZ2LOBktaWahMYYLLuPUP
1B8KmtjVu5lVE7pQHyh4K+RPVi/SzxjOen0DX7meMovLxgyicdQSlCZm++f0I+JV
ni69w1KBPw+yecmDkoVR+0kZAu0Y1ht7dZTqrEag7oJlMhrEm8TxtBhFMmsGntT+
3ksPMrXU86gWXSqgjKrymnV1DzYNDedvrtsbz4XSGzG/syipiuM965cKrAR2abHn
CXj68RXhO8RKJPPOUru0G/W5aQABsUOIJwkoCW37F/utZL4cmo8vHeWrZPH0FShw
RFO2hsLHyOTwFY7Ss0s4hvcV/899hvQpgDG8U2WoQr19rzMG3xtZHWDY9tckV/NW
w7flYn0F4dkNKCbvb+UA9xmsvv0wyfVxeydOSepct5AsxWLEcY1oYzqEQ3n/rz1Z
1bLPV6Tv6B9MnoVYBhNj+TtcVmA/GaZsb616zTQzcUeeJOcaLOFRMd4hhtLEiwyy
IjF/HRAiD7yzXzFkdMQBROlPrWKsL9bReSiVpYuJpwgWI00PZaa90f8xq5+hGVuf
EYgQabumClWYacDvk3+ZhIfQOtN1ABEaF7Cza7kyp8vMrn4PFxDM7eEDKlW3OgQj
vPYILaTsAe5TMF9yBBb8lsefQv/DOG+5WNjAK170zz5jiX1XQQq+GRB3QTuCjc1e
yNruM3845gB4fhv0DAYc7AHLZVn8yNrulpNDC2nLNXwye9gQLGEZ8Oq3otyWo70z
ubSjK3KKh2tX2vTkU2+rekgIclfkorvO9Oyb3WPPGwlDQL75wB8q13GZGgxevGzZ
ZYm0roR9bqkKt0+FwQpHQksI8XLKvEwdqZUCt3QZ2rotrNZWn88qrm6vKuoNZyVm
GPxuqkQ0zADHHEjJevAVJbphnAXNXoy1+bS12iDkgy1GoykZ3wMY4lxyA78CRPK2
twrv6Y1kJcNQj6GirRvJekKXkt+lmJaHtFXFX9NNZ8XK5owhT1Vyva9FFoXcpf7Y
9tnT0A52py6xjDPXYH+YpCDgr4N3bViekZlQgDL3ZnnxX/VF2CyXQMZ9aKZj2zGj
q+JtcbpQn/Wiq0Va8in76QB6TE3jR2s9HWtpgwkzmni3S1Io1QsjETt06/81CpAh
5KGZenJhXxHtn0W/l1u4RZ9qK9S6GznyzyVqwMvjbXoo3HwTGqrCry69YEphMvnT
17PGNDghAhkJJA0oircYHf7q7Oj3GX2sPJqoG4Q9KIEzBCbV9FCYhd4dj1+mRwtm
a4pPGdeW1hzlkBi6Xn6BwjgNcZ+1IT9wdvi55K+q4r9HP1NjBWiAXV0hElitvCpw
6PvRgnAuHUAM72hD2FhskXswjKwSNNHvUQ+r2dDWfno5c4ShYSrxmH7Cr5JpqGgw
W04uf4Jg50c9SIgkSZa0gWYWzKwUJmPheC3gDr5IYZDx+ir92xAmu2jpoT1e3br6
kN8Nz0VSGPrjkTtYbyGECJ0oqmpbInMO3uHpLPFsbdu72OlcypsYHwGnck05+YLy
vgjL+W9kDGPBeJYAyb9N38yznm8vSkQYniPypYNE0POjQQuIVMpj8oNSSzHRnHED
fdHCPitp0sHV5OVDVoR2Fuh/G4WG9qnD43OxLnrt81vl6V5QiBf/TYtbR++qKMVr
UJiWhDPO18/pvIo+v3Pk+jhCYg5RghfaKfqwKGA0Dygr0ezoqJ8awYTsmbFTe5Ds
NfdXwLGaN7DMFc/k6bqWe8V7i/Si6Dfzq3dMaorSgRZ51TDMU1yBpBimaYgF1naI
wU4VrH4GBu7qRfF17y1qtiArjCAZLuq6O42XAJSqNKnpDJB2ymHZmQq47OchhOUe
JnDj6dY/+impMJJTEsi/mvulIGIjPefgVHKDUrrkpTXfctNXKnkP4QoxILO7qExl
XrPDsoaxeOWJvRdVUmbbOleQAh21V1uJ+4EYPEcFmbTTgvqNtEPHwlRr6+9620o2
5rS92T646G48Myn94lIP3TLA/vL3zGypvyjHJvFU3G4WSbqxx8g9q7UMJF7vx3sV
z+xM0jguvmgJWYoqUhZ8gpOluVihT+7Msq3Lni2KAtEhpxddUXEPIDUwY/WP4Xqr
PJWxprxxW4cAmVc3cksFF+Ooc6F6CTTZPXBC2YnSYD9wk49nHEWG97NDjbmHRFnc
fnaYvUI3+tWjk0oXoBfax1TfSrxic3ZNdMQyhickzV+5dc9ecOMe3Wc3MNU+/0Rh
Pljf8/L46jBfi6xH9HQdp4Jxvy11wpR9a8aFi8Kg5jW/IbYwHdmRzpTXyBWgKZrC
43XUMcyOCkXa9gHRm6N7+rD+S22V5MYruqG+cOyg0G26mMyY81ayQME/VUTY0Xwi
Ajzwvmaop0630DZDMyD8r5SzlwhzNTugbVVDehEQWfuEG4gKAt78/dpP57VLGNoe
we43anwHa3JlQAvUQOdCCLoCl/d11EiakFCyTtdKfOCn1pe1SATs1BEcRUgvoukD
8yJEvuPY/4Bk5S501OnkVIHXcMTce0Xv1fL+JN1sakxMMwRcLDw8n9NPYmmSjfhc
nZcqxpl+sIzx2nObftnRUjah2xHVdhOs92/WXUehw7yBv358KnFUFXrBTIUjfXWT
smBmAtP1xNu680IKBSnqLBcZn8aduVcczrTfbX0SyN9y9SZPaCnMX4ybZmQPQaGL
xPwMmKJwgWSo35CoL7eOPDeK5V2yTxDkOfumMgaPnbHi7w53tsOKNq4a1avgU1Iw
0iqqItGdqb3g4tshIN5foZ0yg3Fq0MQkrdFbbBFirmo/Z8x0r2HVeqjxnn7+DFls
/uuYsR12PriU93UtdxWgVPypiFaGcu2GM3dOnSoM+Vz1iuZOmBQJKqrzyZNXONF/
8dqPDftzCSKbpYGMcs7+42nmxRxN6vE3W6h6S/VvP0zfQaIfETlY3IXnkKcse6s+
a3d/y8tA/RDPPOagBBh/buKOdhyMcXLX5b9DYgaLwluCXCzE7b0d7vZia7FQKSOy
RztWFTpM/gqZb0Vu5UwE/ztw/xHn3Nf3T6PkiTjXSfbJVhOuXdw/SeDfIK27kDbZ
X4GQmAi9FvAQ+4xnBQbpekTpVr35Dw3HdPAdFRER6jq0xUGLn3iV+uZMXAvOW6Ui
1A9qVclwrZBOdny5RpRl1z7TT0nr7RqZZVqLgpJH9fNPYIJuU3d62J/I5MaWL32J
NMJ6g58fPe56OXtx1VOtOMb6l8VcR+/aXIYoxi3DY8xzgURq76+ujMhaqtuBAQ/f
gMASTIN5xUWCVvWTM00kuuR1G36NnF5QV/hMwUpuvhzh0DHGTRNMUFQu0rezyTlZ
aFvF3OBGSEYmI2/GqLCES/CcIELkQjB8Ih5DnDGzOk8AI/umkRVrkwn7whmphYOM
f13eljww+ZRVg/kdkyjqSvtczou/kXCL1cmn//AcCw/HH/TNqjLvTNzW8SJf9mfs
sTuKCG4zpRD6F3zCrg3n9zNSYf9IeN/MbR4/45JJvWREpoReDAseYeDlzuR1osuF
Hj2DhpQk+63EpyX629qmczZ1aji0pNrQtVJPtomcOkU99/AxmCRrOXS/l166Y4D8
fAVkXT+rA9kwMU4LpWGIl4nqDZmvtZ9RC5Z4/174Zh9h+654BFaiwp9xp3Au7Z9a
oRRRnqINvZ0sQnbaHvK52qex01JIdwkgURgW761KOB81uPdfYxUM3/1BbOXjeaQq
m+a+N6CAEnswpQDBbrSHq6v/LNwnCsYK63pYI4R1DA0+3MIgLfi1rKj9Bs1Q/wtO
CnXCVzsr9MdCk21wsewoGXp3WsrM8Mu4a8ac+aSY8PSXcNfThQ6lcwD7ZUVBoP4x
PaS+hJiptJy8C5aPM7Q8Y/lRq1rRInaViROA6ka9FC5mVy8iXUMepMhJ3Ggjow0/
sW5M5lJKf6bVQg6tNwd0rIziJDNUJjDCJSMK1N1OvR3ZzwO1LirboATnh8j52YRo
pkeMr9pk69siz3jGja03NyR9AVuMf/c6bO/pnrWmZa3cmmEPhiJTSM/iXG4231r3
gT9ixDYitpqiKC66zgsP469Bs82vGSu4X30h4VfSKolgHv7SEgglbtCt756r+EAV
f88U8F/BaiMC9/ZIWbaL3wjwhG4DHywNZUQvcJyzjZsVFlGXfC56UTaN1dXG5EeF
mKq/6IpJoZlScxOtCgYmullMx3K2Vf8PG2Wdi1l7mU714XQh8IIixy1EB4SiB0dx
PV6t2orEmCcoqG1t2SvQ0dd9sLvlTSB/mZSqEVEYlPYeas8nadQR+w5jbKKnOq77
11rjcfv4XjdlggyfH+OXw/RDWNLJ5yy4P0G36QMCRK74ds80DR96b8NDs/d/cHLE
5GFr+oBAcreS4gwvyEsFYfi2ZIfedzrdim3alQhPIGmnZUMheLM+bWsM+K60lgU5
p7rE6e7rpCDsgI7DFdYouuXczfzQjEwlkUkOdrQFhFZSeh8Lu6x4qFNM+azlIgCm
45mKjtcW+7ojGXorC0UhxF27huwJAISePmDi0+32q1MxC/1MoIy7Syfs7CH7ZsNe
l730SqV5gnDHr+3oaBnNik8NlMNHmMOCsYSj2yY3qHypKddlV0nNc8ZZF8JtXK8T
Aa7ESpbHWxp03Cgj9P/dLy1/MUuuBZ1rTD70poMfXwkffr417c4n88bBNmH23Jr2
uKuQjFCMEmrspHl3iY+FHw432CBOK0o1Sz0ZPLVbvkxht6dsJtCMnmAHP0Hn+SwX
8ODmLpOEIsfCSd2+bdw87xXnfM7ya0axhcklRwts/bVQHnsfkIP/BA38HcbhVwwv
KzgbCyphJKET62SpQJDpvwPmOoDQpi5oxXsnDSLxu4GWTQErx6ypWeLhzx2sU66q
lkpu7XIiAirEKKsth7UpcosRgIXA91Yv+I9UFWb6ircgC1lsfRzxsMXGTFjRRvr3
TlBMCDNU2C+uPJT8Trqk800euh/1+ggpyLF/Qq9wWLM8yeIL3OFkjGn2J53S5D4W
VBLsGT2+Djlh7+HdmVIV639gIC/t/5aR/T+PexzXd65EQV8TaDL1j2kBQBkSMtqc
Je+VmrK1vdFhbGx7/bNlDQ1nwSCNnNP6o+uwfQORcDCgvQvNiNbSaPZQp0hRxBli
kjXXToE8l2+WXBAkFnlqqtjV54p61AdM6VSpeG6PiuvCynZvf43BQdlNDv3b8NSr
Fk9FiAMhNHyTmztpTomIlaj8BLW3HQYEwMao8gkBm2eK+ayx69jUzJZ+dpEYC+1x
2kSlpNRYvAWTNPK0yeXUBk8Xoe+m8v67FNuoBAvB7n9K31umgtMRSdDCQYUNoMua
EYkg389asvHweF/WzaFqDDvWUF3gK3GgeEmr4BhDtZxwHQQ7ZBgUmenewboQFKwJ
wtkbZ7zZBQMdF96sHWp5sooOnGfys/7sHRnu+XlNtBv9i4vJaCCwsrcrUq+P9gev
3FqeQCBCfMLNdPE/3dSEdvrMb87sUin8Ghu3UoJx6QSXoWfkbmoADMtU6Kx0VTCf
hyFOyMBwKWQvkfP+/X56FbQTgRLS99MDZo9onD/ZOTp+lTfSivqZ1esUVl3Qw0ub
g+z4WZoGJUyhRbl+m6s5p31v2BbquJG72AFyu1XVmA9kGsQzAzXApJDVc+/RRp1+
XMbcgnGAKLhlx/Z+ghCOt8rwfyMUBLXd9SibDH/Nu6npLyc3y1bb2Yz0dx1L2eI4
WCdfFLOtjy2wmeSUd2InpqTNIo8cSh+iNk6dfPyq4lDDuwv3BGCgKljDWo4OliRy
K8KwLaZP3PwPYY1V/wM5XnAGj5tH0I5nW1UJcwNV2RyIaurcQ7cH4uVeIRwTJiGu
fJDErcEwUaharN1sjXPfVey6zD3rE40OljjCA8jjJL92qta9xK9t2Aph+f5Z46Za
O6Raa9lzBLDZMe82b6+115DUxKvwqKy0SWY8odh7ZV3DiPZFOwhcSskMGOLJPN96
5Gbl5HhClB0sA4LT0VTQ3yW4hV7xvkaBg+yRdZhbY8CNaga/gTUYniEw37fFLF8O
v5v68CcHIffCT0ANRlU971AUl0tNI5WEnNsuvKeTZgGUQnlCtj9vIN0cK1SH/8T7
4tTHIwl1/afhLYCW/HqdYx5dvOjiPzoJFoXebOU8uH1zmQM5OdjOgbCzwm02tgws
RlRu0sVzXdUzGan0SDQFECDKIV/e1ALg7mlfC/UGqCFuFpk6FryfrFfsv+clxlt9
4/eWjRlk3OINi0A4TnE2SlMyDCQ1sy5kHNhVOGl56C+NNO9qMeh6OL8Yl6HL22OW
FvXvNXtYkPfPAY04nbn765DJisethhJZg0sJkowj4tjKvq/mTcrbPAlYG0ia8JEt
YVULM3inviF38CFUr5NfYiDbZSYQez4CjfdPtfwXMfwRXmz52sZfXhkzwmUeEPw9
ac0p2mAEEj87i2VKW74ze63YlHaCQXOJ4pXNTWuhTCyYmqj+qJaGt3ofpGfHK5BM
anwST33BctzYsEK6+NSdigijTqWgBwDdtLN3IJlxbFLssLvke3jdFtObEsYSaB36
evugjJ5hXMlDJG4cYcer/HfKVWL2Eo+eVSpluNorGEqpL/a5X45PNUCBmeXGmzg4
8hUNDn2MlId7ilpNBY9wGQONC+SqzRj+ZdkZOP4m7GQZLW1r9oXxxb/lk4XQ7q32
sIckHNAt3qK8GweoJtB/ef5+TV6bK+kehNfV29KHXltQk4RvHQ57K6+hUofMr55q
DqsTa/QtKJlf2HEVjP2PRJ2x1uWkmmMxOaVnjCHShMmEHs0YtDXF3OWrDfwnOrbE
mgRtNX/LApooBpDhVyZTJmbRxvpX/Y1Yjy1wjzLdr7jMQ93+ec9sxySae/y0xKqy
FXgFINCW8EG7n3Dsps9enNO9JhTFI1lxocSRp7aOAEl55+GEIHDPpEoW1LL0Q3Mo
A7/e6jIaKOtwD+z7CYZ9/MRcb3bO5PtDx3Khy8Ylbv6oAgH8V5mmRG5PulF6KoU/
YXhFZ90wY/a2Ei7Uzyf08GqsBWiQ8qAjonoNufrd43PXyBY+aX0hrVD5t8s5dnlb
O64V4FnsiXr8RMSFfMo/mYqYXPL3MKZ3QIgG96SKP8CS+UO/UFGOYnm5Y8zXClyr
7Rym5g7RpgRO1EE8ysZnMudHsaX1aW9DOnkAQ0nJFShpXuAh4jfQftXe/0DR2iWH
+L4HxG76Bm1Lv3wcIhKwENSIsdxp+irCZAX7X4mgm5R+WmlMIvbeBph25GAQEfzn
4Sb2C0v0d+e+nwg+7pqa2E6nWiL8Y6f/r0LxHo2ZtV5Q7sslSHlhOq2p779lZEsQ
wUsJ9zGpJPrvvyjdMhfPbd90vbOOqQhKuDehfnhPncMErnMKXRbcMgpti5rQ7M4I
wxbXpdmxM7ZdAPMYJg4Eb6YhPMAE13BGsZmKfDhLM4j1W3aEkql2Z4UzlDlOnNi6
vNXSKbElqk3bMpvs57GUoB7xTG6TQbpFu+kGfOs/plz8aZuHwdLvwb0RXliMWrK0
3T18wTuRbO8nHqnQN9f5QAVDmZrvBCWrfaOhLAY285YwqTqbw7x/7/55iSnRxVH+
Ck9d7lymwF1e+uT+sA+lOtu4HD+url1jQCzgD1aUFtOdQ/T1chXmxBagb5d4OZiY
I+aCQStpNaFEu9nZuGSnCEg5ehc9e24cNQokOAU8CbKKZzYtdPDJeoCs77DduC13
Y99k0DnYpNAZddNTpRKQAm4MlZzO/hSjz1wzOZBOdoTM79mDkFEo/Wy5y/djDKus
DS+sQlYmhtmCmNAOMfCfag2bPGwcYleApoMM6nZ+RNAcoE1aot6lxI0uKnDNuG3f
WNLQ7Xn9cUbyG4CUhqkdX8BuCNZnk01cQkXWykzN2WfbXe5PGRA356Xrn/2F5P9E
V+j2oR2YSONrOV9ZEEBc3h8M0J3BBCmzAjXG6DjPa24Pl+MTQGsLF/gB9NQ1mYyw
adaomQ3R32m1fsnnIJan4H1KD/dUlb/14zPFCnGuDqUFpn+TDGht4M/QuSWemh6l
njSq38egE2z297nNElHMru6t37RRlRH4ahYnQnA+KNi4oc+/qd37Ye2Ap1Y0J6lW
RBrQ/PDkFL9PMtFBRc8URK9UOy0HXEVg2CifBpXLRDe7zZyVKqava50byVwT+LIP
+8rwqxLssqv06vy8bOrKY8xlJIbx9IGtmcT5Ls1ZOGARUJ/Mwnpx6mkOCJPMJkZw
IRglLzxbIxAR9aQzntq1x+n4w+EUOICYE1q2D6cfDAQ5Nv2Hlo9YapYBxwcm+6ZY
HD093yQzf2L2YpRDJthHmdWU5ylG5xcPIreWkBQBZJQAqtgptOTWMPaylTqnLePU
UzXv5loI+nDwhxobKFX8ZhVrMa7yWpCWPo5yhEsYbOwDyxYfP4bY9aJC5H3/NaRO
5CzMahYyKyUBb5fZyvWVtxk9O57hOq4SkrA1mxIilNsfvkACw79HEFwSTaqBiv9f
1h/VkhzhGSLaacNJI+0zJK+Nqhtl95kEwq+5queOGDyBXvv/irMmbtohGGy4O8lt
JqgTSOyuNdTlO9bCI1+IPT0aJFkPL0zHV7hP3sdL5PLbXh5Msbx+nvpiqq1L8Wjc
dtSuseetE4n38XxHGbKkh7sUuI2kFhx1IBCNAwVPBOQq2hrUNjkraBwwiUJBbxkW
3PqktYb+uQPc2gBehwAf3mszL2rbKRZxovDkGlPZrAp7Kvuz2l1glptzzPBHmm6x
GQUCe3iLQG6q0Zbv3Ncera3CFu8UD434RZuxerrontl1WiKotyQr4Fc746MuqNn3
pJktlyk1+oa6dbipLPBKice03M+zKCsI1Ps4evDwxScM2wqGcZRCDjWaRi/EE537
/0N8+68UB0rG+NNwD2ELdBvF7uHMGzx2MFdVzMLR7C2GerrRnv5iazgTIAzjdC4i
jZW50ihjSKHewTxrgT8Uz08/A7+edWPVnP96qs1AEp90DvqHPMxGeNgG0eD0x2iZ
XObGx+/p6YDg2fZcR679UkymoPZzRK98quy06gRLfWlML1MnZwjngXvT5QLGidDu
pmPzLb324f5bDeLRTABskuQUKmjT600OwTZVnr8EU8F6TI0irm5xkf5rRtBKTZtt
usvjvAXxv3aZK6Z17ErgnGW0ZF3hLj7MQ4xFlu1ErgIGgaHDTF5mIIzJkBRL8iBf
G/Zdvx3nYTFKLNSzuWeEpEGWnwpIZ/JZfc00fcxWA6t6H4p6CFWYYPNNvJKExzCS
pj20rEOHJTEuxEbd5FEmdDUs6xErxPP4q/GmUY9OWZNdgKRn5NBv82UDW/EwBuBc
hqoslTm1OX221sXw+SU4fZFZqig4NLpfjxDQG3IA5Qtgyk6IGsXYe6l31KFkDRjM
pUXoxnlfpnmZLtCHa49CxFQA1zp6/ZbLRhIj/Uh/3tpcFnGTLeqbCrDQlmatNIvi
Uz7m76ZxPKmnSjFo4H2HiJ9zzHh5wnmk22f5cCYGUJlCcwts5jEQ2fXIqN9T8BkM
IvFzG93vMNyY2VsUHHCxjBk3REf9GjuhEQXZm8fZhtTsxemNd7h7k2BWNruIa/CE
2iY4uWB5PBtW+N5Ndgc/Jt0ApG8aRDwlZ8KP/wl3oN4J19tyRzqXtw7F8lDfIEO0
b32FDtjUx2uALm0F5TokzCzWPqxG8XmS2ppmVx4eBMLdNT6RKNmqjh3YlBfkjyD4
vMh/CLB3OyxPkQbuHymbKclwZEGT8xHRAkn6n0ZrusawAYHfb6+7JMkZM/3loFTv
8ikD8mgdrUb4iKTr3G0lwtVImXlVRFDNErTxz5t81kzYTlMlnNzlL1kUVRAI20hR
qcxhrRkkV6MVPHC08AsofptaJo+302qWlFKN0t69qyG3ilC10imBr4KowBX6B5UM
9j7L6aIH5nFzsxUIiev7E0MNcfFKjpuaXDZcYWcMqQGbzPhD7XoqMZAutHMEY5Dg
i7RgKW2VXSc32X11zcHG601jrm7G1S9r38VVqLumzjZrsclNFTwYWyooTm8a5Sfy
PnUVrT8H6bET9oEr87wxfIgyaMKGxDkxdTCwV9GovN9z6HH9b/wdkOWFGjukx2rL
n4lR7KMg36VAe6Wf7jeazHTPSdWaQmAlbxVWHzbrZy27DQG7J4Cl/CZoy47m1BBz
8XwiFQA5px4Vkqx15Cyr7217twYY1L2lZmvSgwQMrTnol8a4L1/9GFVZ4HROg+Td
Mwt/siDFkLTyzfRc6p793kFhIOSNWHO5i+lHCYsBTo53G2WoC1JJH1T2zgy83zKp
sda259oOViACxYqgl3N0oo6PRvnG1iOeYE58GFrZL5lSmPa9/CtNDV1ePY6G2ZL6
zF5G5hfWtxmcDkWbGlz9zmW1a3b0H5ElJ3IQ9aqh//yAwQT3SxfD28lRAffnvPo0
tCtpQ0t3PG4WM7tH8WRhdG2CyAxThD6/+0Ps2T0uh5WsftGz21ByuFSN1kan6I/c
SOF1tDcpilhlwnX1uNFZpV/HV1qTw0MxfqgFA7addBYwepMrkR2i0oWhasJsGxVO
FR26ZHqAqw6R+OTBBNnSJdhqV1szvLHylzgrypI8Zt/rRYFJpKE6JkzKf/8jZb0l
kXBJ0djqM8FfV+IELjv85DoGeVW4pjfUyqGcx5PD0UrKFifC4+I0lCXPX7xbYImX
HEZinzDVTNYKWtVlGfwbStLFM3clBgyCHPgM3SdAZNiYLYOjxiHLvfDrpGkErZtU
L8PGpWGYhzFoImuhYgyOwycvJMXJJ1Ah2DupyIw8O537cWVVkx85KdWh5XB1LhlV
Y9zUuQrAiW/PpH66URkNH1VOF/6dVDGF8Oh/LIcPn+Vkt1Ic7IqwtB76POCpog04
/iJM/SUyEfVjltAGkvGA0hH/BIUcRQPAV20UtUSJ7cSD/ebcAY4RIgNmOTsjtMav
pyqeyilD/4rQthBauCxoFB0I3aTtjgdPJqIrLJzTluqp9orzii7QxOpJ23ipWxwe
qK4udoaLLH0QMRSw1NbHORZglCTvWigqzL7hB3kFK8SU3g1GPzHoT6eEBmw7M9iL
MyMz+9b9eHujZV7pz3AazdOAy24yrXdzzYPBDHjMY5TUsIVXewYYo61rQwDKMTmu
zDm97LMeomwYCx8Lo+LXuIXJ1l1mtsamgq8RIk12+7LbY8Kavs2kH451gHOy0bHP
rA7jP9xV+PtqCFOX66zcI8FkbsEQNBIMVAYMaYNdh6A3JafYYGf7S+GGPmCunFGO
0PcYHxvNLjI+q5TDOb6+A03gNJZ3jdRrjsq1c1c5xHVf5bWo5fTtRApGsneJUu3Z
tr2kSYPEFsfc5+kmG6XwcDe1UZLI2nrdPaEZkVTl7kg+8xatkS9+tzsZtrd7xQOu
iTGLqZWUQLbIVjvcss2WXgkWm2HCJfLdVk/Kpw+Br3T9IA8Oqa/8i9agd2Vl49WA
GA+sUfcjMs4Uhh9QLXsZtSJVXq3paGtKARmsx+sMyKWv9U4cTIWgjP7A5e6JU0hG
BJwqgKKhCIGVEsy+vRhLaTcL3rQtysYVZCKLhqMfttEZsYQ6wVmRAGXYqktr6wE+
fFig/3KmT9a+r+sPrpB/UoUxJokGzjwrcQoudKQOUTRZnZqQkaPzY08qKTV+DdKt
yH5PL9TWjWZfv8usN1EeM4Zx5CIuNdOquVgQKvh8Cqd6qICP7QdMtJCZcAZkuN18
Jm8tdeOnaCFxkHHhXwp1gyh7GyO0nycCHgrg37bUs2rNul4RgxP5s5MNpZ8e/Pxs
TXmSEXY8lJkD/Z77FW/weOSO3wG0RWFqXUVyAdjBVvjas/UCh8V3lPehv6AI9v9U
njwhSjfmh34ocTektsRbYeixxSqvLDcZVdYwZFh71qdwffDORwP+Q0Po+oxraxxq
G7MKKZuwZHB0ynJCNgDZg5sdLqJjbg+sI/i0Ocq/turpScvHdxq1J9mDr43ycMox
2U0WDabT/eWJmppUmIKv8PtWV4krLhDGJ1UGhDjj+2GqFGGTyMw0bRET2hy0N/US
5TigmsQX9PgTFi2ZtNQnUILrLCH+/Y/uYVVBMz18jk3HgSNncKcOXVgdWnjk+9mS
k7pHhKF0k/IMudCIuO7zemyhkiCvU8PlcQiWnPeeGEOe8hAcjK3J7L0Nu9e8INvw
8QmjsQFBTZa1oAWN5iDlkalPQ9JwiOXPOu1U/Gm7d+Ss5mM9ggK0WetsJ/8m/K29
C8jcSKflasVu44SWO8dbux0v9GhiMdNmR4dLNcCVTgmgm16BtTEA6GnpyxwGuNnH
UcT0vboOaongv28Wj9DCQ9xlU25cvvNZXEj4YUAHN8NpTKL5/hjkN8EH1BsUNVSr
4Q2gYd9kw8tKlsFCaxwppjy8YTAgGlDrPoVnKzF7SBbcwWBRKDfnlZHFIxViHruk
6V6ay3TXC98GY3VyfmTW1hogsFRAWAC3+tDeaaGoOn2Y8jObCGb/HZ5hl8XiUAqW
THyAKc8hGesZq+dUw7O2r7PbZ3VBAvHV5aRQBTe1lhvRYEqkCb/NQXbPuARfY/nD
YglVXsQ2Ukr1GsLJ5qhnvFOLOvB5hfGzoulTfnPHCUuH6Ze6Ynisv45Xl+zMAef1
hjclQDuZE/TzldIyrOnLLNPDqoVK+YIgysceYfHuBt/CoyullVxgWIWvIo5Fzmil
ot/TPLS/V+kh4/TXimlpDAdACk/1ARDufsdwguI0ysni9a9QXvw9HM0ryKLJwtrT
v0+iUqx+R+l6Hd62gXQ5BTaJWvrSVkgx+okGDepV1MAY3q+BMjWEdkj7fagPvxk1
Rj8fst9D84cHpuN98xxUVMeVzHtE7Rbho/8iwqwxj9WNaonkWzyuoRyGCGAkMxRP
rxvytRmPC+70QjKBFcSNmWsmsYaFQ6XOfY8JbVs95k3vAPMcZ6j+WQHlZ0oraCza
Q2FWKRIkuGN89qKcZcCMpzbPRQGLVAQ3pnIt7CSg6IG8m4TooihPGmApumad4NEy
bwxbsZbyYfmbkPu1WzM3GUQRJLzqSMrF3VHomFv/KD1XyrZbOydgOUN9sZe6cUJg
nMYQWA3DWY1Ui6ww6g4sv/n4LPyNj1scg7hcReUwLmFvpWIh+jh5DAb/w/bJdJZc
ANcvhbOu43Vl0jTckkjguSWU7mOH04i1NLazKoRFlrkpU/MKG7214vionA4y0MHU
5tbpzJBqC53kreBKgPIgM700HEAVj8qSJ7RA120T5MmgcB7mMCvoiUM2zccApD1+
qOh3VHgzltII/4GikxFi0UpFrRZIV7kpNCOFcg3Rpo37igRYRYyrfFMAVUtZkmqa
TdH7Ilsm/SEt7jNMO4q9S6X164ESFE9iwHmu2v06iZ2fVZxa21KyFCn1PJ6XctpC
OHzrxt1nayBx94mRhTPnf803sjTQhbZqJ9w9CIdACU5tA5RJKawwUbE+hgHwLTwt
6TN/JoAia1l5qd/IQYNdndB9EjUpBoS/nsGWCcjDLr2eVmgUyKuJFzQx8lDjvDhI
JNwPTzcSti2ccz2tn9TUMLh06m1qfdxjj9ZudboyNHx5xrFhxI5+rDaV/8QhZ6Re
l0/AYRQ6RIFfDyU5BhE56UnlNP1MbGD++Mv9reOJfLDHVJry1aKLJmkwyxoF6KDB
Uel+ewnlRjRIhvruGTQobHHpYbwzcGL1tmiJYw3AZ2IfB27Fd6T2a++qlrc0/SsY
h3XxGXdkCMJup/c82qA3ITIHU8nPBkHlpxLGh93oZjcmzTcL64JZXJ9NJlL9uNMP
1kqaxu2SMKfXgEWf8MJ3dsAMERmshOYQXYuqa8DkmNTAuyEW3faHA0ExG/8Khj/H
nwzFrGNPXnG8VwWbOnra1cf5TwPxevSibtDxjCfTpYmotKzgP5YRF6CVu3ke1D/l
iz5t2HkhQq1Xrw9E+KhXQrh8gy81AsaOOEsk5n9gcFeNi71BtZQ706jg5k/eYiIF
Vqcs0FuYscbB9qEum2jRlYWGTAAoJydkyGpTaSHH+hlUOf6lfBhTXlHZ+znF3Rin
4kCwK97seXs42m306JxBLnj4+RwFFEHW92BxlicLobh6bpeEDxAkiTX0j6ttAH8h
AU8KrHIvEPdcKL6Z5klvcXHJehmU1ViS3S41haiMTPY/+5wQYHaSUoR1B3EdyOV0
/SAQB9F9iQNSUCzqTeipVjUstTCtX23PA9Fs5uGrRwg8RuXNzcS908pVsRH7HhBS
nqx5cTTSPwxYdA6IjDSYag69mjK9jXZSiNY/fl/s3YDouRE7OZbfYYCMvvtueVqt
qlLb8hxrKxkeUQkXrO/ObtQ3oRIIxHgCLkJ/as2wwXn8VoQWu+Z3i9OaZRMgP68B
k/9NyA22nZBmV8LX4xvlqtqbxOuP6lv4c8DRAOibwEEX2cFzeDdxH7QnJFuzru7x
5ySqWwhiUqV/aeatv7VNTX5VyC0wmVU8vtsg7Q/yQOYTOwcZZZntlR+lkQ+C4JrX
PZ/Dzh2+E3Uw5QcyClp1usjg5zVfrQq3BdkBd2OtiakmMPKCnIF68nlDG84Helvi
ViNrUo/rjQ+YVMJ1cMDRLnRLDAOO5YN8Zfq7OYIjqQkblcV4ufUH5pX2TojuxRqR
eQfHGOQZX1kI27M07QJP/xtwykP5fULgVW3FTfONGd7dmWauPO/vNx4h9tI4HUfr
5rmSgJC451r/xfRqMRhPC4zDLOFPW9OfpGKtUefbgv4UdfcE1d3ACYBH+wLRvsJW
DIlAb1bqXsQ0Dv1xvzSEfhc4yYDDVNHZgX5WwxwLSwtfOmswDAc3pj5Xv4AgsQcD
NVp912532Sa/pYa2Y5AsuGEw5+wSpSLEfXGca3oOaUsJ2talzW1RXA4rIn50FzeD
TKupNfWnA8QdGVVHvr0nQ2X6Cr18fty30X1IfgiI7WZZGu+uT8c3VDeXvVqk/pRW
kPaLMt2GRPl3yGzVhAp13u87I8R1J02nm1bj7KUZB+hBA8hm+VDczsRGwnhaWOtc
XKYX6LtjMsUPdhD7+ee3U+pVdrXmI12SogpCKJRkUt+zr/pwUpNDQiZ70nX4qwPL
PBV9k4ZsCKuDvcBy+t3Md3GdNJYxFIrLm1H58ZG/mtefUIMY7ALd3IwE9TRpNIoo
Vy2SjC4MT2LSXpn2Yu6g0rZd3DI4m0GSt23NaMQAlumDZ7o2xhrrZ2GFUxAoVUKq
uM7oFP/dLar5ItLSpWZ//Z/TJOBgM/3YvkuFR5EYSOyWZXj6yHu5kpA1qztsXrcV
TOC+DRYDORGC7kO63DjgbPv8EQocRggyGb7YD/KulUqtkGK1UuRcMLKfO8Z/6KgL
czV0wdc+ltxkGAp+iizh7x+VeqmrYLf3NTHQoGv6b3qZK7Qy2Q7vNNGXy8nWXE+A
UnUPeJfsLuEBtPleGtlYjpI5Q7cYyhNum/E4TKDXEM7VCzTRwAIE/hcPhlzY3xTk
00DOYYPP5+5p+iUvQ1uN3OI+zkCVJh+PvPFZ8uY6uQTx8wTgvYbQEkZEFyWHCWHg
AnPkX3C3Wp+qv5cQ9OHJIMJVICJd14bjjx0US2SCcWICrqgVRuPL1kS4QpqOYvGB
DfDeZEfXtsA5Vv6xr3XqNn+BDl5dzAmsl3ElR2nHTEBeAMwxxrbNcB0M6jsTJcqc
IbhCVx6BuKvOKaIbi1gJzYUIXf8fVm4oswZ5UsTlE228UsL3jHqs86TuNf1M9kHA
cnr7y/C7cPI/u9MJ3XMX5avgiqdW0TL5fgo12Zmils2ROasneWd2HQQJfesH5FJM
a9+zJi9ThMsqLijmOPtnyATWS71cc8JCTTf2iORQkQQ5BDA+69BY59VYm/AMt24Y
Ei039IKT/6uf9BzSs8htdwL3YaY90MgObTDeMZfzZqk8EisgocTTig6Xhm4OygYr
ARJZoVbTXSmJSiHjgc814LuVFgLWDRIwnRQ1nuaMAcYyTWx+O+g8sZrdoyYp7Zwn
UrhwShjD9KzRworCLFCq+Qxay21Pqhccrisq32xKm3+hjUsEYqA75uLJSBh24vPZ
IvWenQDw6Qa8OjXoQ1KleM8Rm4wDzuNXl5/0qnOX6tjnp6K6RstBqrkA4GOQ1iTt
VVxLln/prgUn1OlS0AyQ/qMrdwPDjdT3AQUc6CdtvjDB7EKscf7pvxe5sTao4CNQ
v7nZ4P/1QrcU55fteqT9F7N9eE7QVmDn5HrXJ+SrUSC815ONdRK65dM6WNEwnzNo
vdNjCgm+UGSeZqhggqsuTwl/fUeoE2iI05c43c1lHwUhYVqaO9YWsWol0x9SSSJD
i9F9+gDCSx6lufLS3f7Y6GPilcECW24/gSPjx5bCQpKg2orSHbyeaaTeYKItfmGC
cOZ1QHgP2B7ciyKmBGub+QyqYX9+UrGqx7ggsnvCWFtqWI0Svb9ya4Qhq3K/s3TL
JifTxPMp6fRS6vTLNlhw8kAK2B3gZVyIw3qs2kQhtpLbYRB5SLg5TOn1xQt+2DRY
oHkj5uzFfiiGgkPDI3YlAtGqoPLbnHjR5dBDYang07K9XlhKbD25K3/Az9i2uPsC
uBHMvkAiXpOh2TDLl3kVn6O6WqlmeXf5Y1F9GK9sCNyQGOlWRzMlaphQvi9cBYsR
C3LPsKg7bB18aRk5lZR3a6j/BtGXW4bsFkN1+D124zEqS82xXxKyd6fGV6oR15PA
Apethvmz6SM47gxCEsJfK6goRZmDhiRRzTLEphmzdsq7Nm2Jgc6rYj+RPX04NxKH
aG9ZEZ6b/M9EHVOup1jR64smu887ZqosChlNBWhaPUXkprKyo8gZUrL99xLVizUT
SUjQdDPS66BDgQhnQcNeqDwNhPPKZjPfhysVBwdsOapIJ+jSSFXEb8GGBzvP5RB3
NWJ+j3a3LRJShwcXC2fM0PkNh4ILa5rSOAhQeWO4vMbEWPwNN1MCkJxbMoh3FVwd
KMGNCuATDOUlmvysxYxYqjp5n1K9hJOkP520bOYdV4TH3Jv/YxXqv3OfON+HugUP
eXnE/AiHnVdnlHs7I3pDkTA/ZveWOUpXTnlLXQio1mXard8dpAfBGEtwi+LG4uR0
BbQWgaYE1bhl4lvIh6pHt7OForU6OwOmGoZXfodQAs5zBQDitrGVjCr3TxnHMtph
QTzDGn7ZxMBE5c/TryLPctKpFMazwNxJYHP8lkFlgbsABoeZRucT7PcEfXJf1yyF
FxF0L2Gqn5xHcacMIwWAWQYSsOvBhw/fixjQMrs9LQ6f6CeDS5s/d0l5SRKYmcLJ
075X23T85kdfYtLCqV19HXYTefi497eQAXlmYiGTImQOb6lI4Hq2rwc/bJSDnSB3
SSfJmx90iTCXV4be3A6Sf5EbJFwkwoRgeNTIKiIoF3rqHJJchQfEDXsUdAbqaskZ
O30CJ8TyfBKcf6RuOk3cOorBGkCfSZeXxyHGXjaqgSVDgo5scAi7cNwPDPZXPiK8
94Ox4e97xcod4ElgHgePomuoJvu+ZFk25xGhnSFCOO+U+zYS4IvE6zl60MOI2wva
uKvcOT5GWdefJJa069oLeXxXvQffRBpJw+tnsPLIdOniXiMsAN6XIRzqbLzsI1Z1
hV55JseoE4XfK96NvKKbeid1XeYYtKRetGW8ZObUrnDwQUb9ncnh7snYhGiclC0q
YQN6dzGBRrmQ9EAF2VugWU3OSgPl9Jg6o/ptSQnOzFykCoLkRTAMBY0WnHGAAhru
tW0ixI9WVZ48KJdNYRaKVWKO+i6dadgJkXSg7wqtQR9lvC6MM23ZOsquIVN1JhfM
MfwZ+1Qf9DVvpJB0/6xAf7tFDMiNVzhImSuSUFs/OSzAwLbZzk7w4hCpnTMrMkXD
gfP6zLTs9no/T/qBAZCyHLKN3nXfv2oklkTPr0jEgRPfjqzKhLB5Gdz2xahXHakh
q/nzoBR5ughkMjuyuZj/cRGyOH3516+n1NTzuAr7l4KV5vZSjG/4nVwRJoCqP+3h
nXWZ7JAHMM+VjfaAjxaiQQpPOpbIxa+hoMZA7s91w8/V0dT34i+YdDPQA5aksHsd
RZfG7/iVPMPZODRFagNNaBVXaAkPmHLLxjB2PNGM+pSzPMN0+daY0tDFiIg1D4ko
q2ZDnmUG0jR8OuOWhXYwbxa1WXMqrkE4JrCfv0kRxhczWeGFvFGUdxzx7MlI1DsG
u6PKKHR7OhyGJZYw3tTd2dF9LZfATrk8SyA/+7BuSBXLyYlMpnh+s7bLrTzb3cxX
BFv45SlIlf2ajCScoxM5AWdat2GEa+aAwXVUmAX7yfAuNZdHKZMJuI7k0EMJfq25
r4Yd60izbvnbfWRQ6865/SqXtuUXJhJGiwFuAzBBrrwIRKqJRSUjnA0Oyd90sp4A
mAFeo/4Strc/4SEyyVrWfA+NHic+AEZR2rrXVV4MKQlQccduT8Pngvkl/nlz9GR/
3H2Ae8/Sv2nYwrCcEm+QMRumGIb8Exnogfi3qt37LIqniVygAIvhrfze+LS7sEnp
ovIWzOOHLeFmCTx8lRl3xfYgXR+/224YP8DodoLbOPH4UuBlsTSJu7FsDXX09ght
ysSVU587PcKOsUvN9G5r5oaaUAEICIFvi5CM0Bt8VuF+fnsixCMFs6QnPJEYJN/h
lWq7EfDG5GpdZYTEKv1ug3/P+1UVEcglhBvuJml2Xr+KeYk9G102lB3XRJQxlZR7
99XCM5mg4XADDpHtN4cBhcNDT2cOcEObh2BZrxtsI3jUv3y8ReAEmVggXvNHnEJV
FhlgWYecE/zjFg0RPL7hl4hEqErlSC+exXd22+mMKbDUVHwFo7x7upSFw7WxTwib
paqdLtFNGSUj5MCkfQapiv2KIYkHemGLLWMkvjjPq2CD9f5KNmtxBIozP2AB+Yh3
e8WBR7X7D68D1VnjADg/K0KlHeuYejVX0cHa5Xh2pz38DsHB4XGO/FYwUkh2qM4l
yZfGMw9Jmhenq8JVGskKwfPVGzT50SaDkif28czmAOs7Ej46Pb4uRsfVCADBmbYA
Tf/f4o5dL2Oho++DAL2OOTcYqF56+Ymm27E7gREcD3+MFjZn6FOLnnxxHxIwEwKm
HC8rnOTvOyLhRHqiMomiTmRG23CunzvKjzRb09yRH2XezSqmdQSEL3ffjk1Q3Re8
GBt+8ZURaLs+iF80TdOr0Mv6zBMwPrGlyC0iyBC+zOxvSra9FisakC4lHMeqjigO
EmlcX+depc+ptkUNQ1JyAUd4Z92BaTC2A7oHmOx8yGzb/trQL0E1hZ4HamuIEQUd
iBL3KBUv+ZsQEZ7RyUYtWIH7c/Lr35YY776CdsabpqH/yIHWlCu41vGePPmf0IL5
ztbiw2U6dM/yu1G0tBmj1++td/4/abz9yqV41lm1Lq5ZkYcp0F8CQDcYq/y7/mVn
kC9I2P1JdY2Cjuo9yOxFu8sUXiQkkhI5Ov+EiyX2w6mqxrzz98TjXDZasGoEV/CX
bHXW0vTC7gn+PfULNzuOhjh3lwYF4nd0QtCP9/OhPXEzq+xykOwe0AJnfMqHwQBh
7D8rnmnScB7Geq2BoCxoAEhrYsF/ViPUNih3LuyaLb3CBQqLjSDojpzUBcPpOiEB
CjHLcsrht2BkR6SN1k4piWLH+4c0x5XujXyod4M8aD78x69v6m0eTxpqNAH7Hmn3
OM/65WL/mT/Ho/msC/sxNeoGtyafTEEK49wNrNiRsTwNszEWBXso2tkHKByeIsZj
3Odq+vGr2HP7zDlsr6cHkFzo1WbdrqJx0WE6tdLjJDTA+boLimaANh5/cOwEGDEw
iikUTmeub4euo1xAcGTPj9kfTLnU4Un3btKAtxtfNyu4FZi8IFB0fDURv1+lQx62
OU/zHCxdUr5XbrDiZtjdOvvkRYk4hFPPZ2M/OUQDMXDIeT/cSUYO3nSbMFSo0v/7
V+NYUapFeR27tIYIzsCiCj9ZaUBXGa66dK1HiejVPxcA4jQ6abNaHkxIZqcnBqaP
wQli7lhhmKMgOwsI2tfjxgeJ48zG4h3W45aYgZSOm0owcWd38N3GEx06a7Jxzzhd
AZ5iUdRoJm0G2bwUrIP11krUhYem3pV61mr8+3nrDDFFrYX/wdP7vkbgSs6sDs6p
dsvKSX9+ijxXXHsf4BvkeagYGl5LRihvWHivm4SieZ2RyqOmyXt7cxSaryuRBvro
1D79hXYI/YMNJYXmwcKs5K+IJ+yF+1v6d9v2tg8sTPr7jL3XhIFoULkNNWAMbarQ
ZF3qVHIb8s6bRXMSQqbi4VfDHL7WnTwLb3ThGpo7DsAJE475rQ27XrgPTobSRI9t
x6wpUQEz3JDOjyxDaEy/mOYwEa7/jqG8e6ju404HqHFX1FVzO/YynnmGalzTmc6q
iFqioMe4PEMBHE7QGR55Gg5tVD1V4L5uwpmCFusZlvkNguKc2Dpa1X9F4rzcMWDP
Cw97s4LukvoaH/7O3on9MG2tO4SqpNIR8dMrTBfjcZ7ESHzngSLKxG3gS0qrltyY
S6qii5BUyQ5WqtlUtaIEDUbm5M8yUibMkbs2hAfzOgRjdq/UEkAw/eH9NkRUjGXe
yQ+4kud6elNgmN5wXGsz5f3s7YwnoVlDZYLn8yhP5zGdRr0MacnCf96OuTnqVfNX
8AgNDDJedshxvJpdS1yIsuDcfLBoSXR3PqX8/8Zm13Ks05YkDDq/6Xc0d10LXtyS
+hJwnGz9ONrBhpQAcpSaZ8Ar2JRZOYUupXUDKtSyUVv4imj2lUxHEYCaakWH7CEZ
SRsYOVI6TnwGJe/wbVPDTn1gVpiUVn8hfdhQ82miLCRQSUehgDGDRdrJBFzK2rfe
+NNLkAylFSZ5qtpXvDjxaP2w+eZWNoii9Tyx/LLEy/GSEcyQZGFbFuYqKjE1g11e
tV1DK3C5Vfwx+Zvork2kT8fzO7O8colcEip0pWehoptVUQUN0eWq8VmRrwzG5G7S
E+Wwb0o5vHVhmAupLSI1UWNbvDuYeJyxYtHgIWijF6ZIBmpKrWx+9NaAebWjvX12
swTpcMrXJ/5LARdzPnbe/9HdYA1rgwNVaZqkLrNvzqg5U8gB2crOFbMgd4ppv2Zn
aePyc1NP2F51ciQSfupJFTbLhZiEkuM5vddjQ+hpCGi6j7y73sBXantuqspbuuPb
jFT2uBMy8h5TQOjmrd0ysVoMi2twOnTmQyy1Htx2lR7DROyrPym2aXSd5nYnV2A2
aaEtDiU9zWbFZnvco54SH39/Gh6tdD58f6EP35HkyHJwDkk8ir118rpIGzKkYW2Q
YR+N519zdkMbGjFCAMxNjfLXCtMW3c2MdsnMdFWcLipZIOphYpAGLa69m+M+yLgy
uqCn5iJtuDWJSrbtqitJmGn8OeR7GSUpzm5Zlm1L7z9+3vfd22A6ggXc8F8DPoEC
vt7Z3PZRabMK3IYvSiuvbGdTM2XYdqhHWPP9qke4bbj3RtvFEEFYR0EY4RMzZiT7
vK1G2IP/AoSFu0LUXA9DyZ0g+Zt2hAltpQ7ZUU2jmI/4IYjre7X0+J01uKb/AaL+
UABDVounuBNgwDHdRCNUeqnavcZb88kmHuQCvGUdxNtlJgzViLNqBi59QfQ3DL8E
1rroYdhT+gsduFOw1MmTjRkl9Fgwb67BsQaekqBMenNmmGNHBtZQGYJ8y3FkEMjy
jhzxRm3nzRyeFnbSTJ7D6Mem0+OWVR4Sualt79Jek9oz0HF9m90qUPG2bsWwxAQO
R10RGmC5p3v8Kxp8+qbBoJXdL7gTYEn5xasbZ4bPJg4KbW671nx/rUKZGOlHZ7/C
DjAziqKFy+3DevwaGHLg+DBd9gh/EWUw2z/Z26mPU2YCYkaTwNhaqqWwuTq+J52z
FZM1eotgOJM2+yvsvOTv9tII4j8D5HX1WvFciyt481++s2E/HJiFxFO3CpP5CAiI
CUlEWw2xg06/2IGWrkUp3i8RbtJgr5EoetjgMHduEIFjPLvJVOQAiLrKbGP695hg
4SGkzQeQXJ37aoBVViHAJqjz4ELdKDtZqD9Ef5UB5gX7UJmRBF/H8qvNddwVA8MC
arJ4/RwAEBwjdoeXYQkoOcGsEUt8jkkJ1O3cb6blH3MUIXJro3o8MlVLR/10Sswq
0djSkpEWbgtV8/n7PpAdwYlnKv0an1UJ1je5M1UfBuy/3wtK9Zt50As7a/qN8zjh
T8sxmLNVF9wGDKg/Mpn3UgQPhbqz3FVfZH+IKib183yJjtwT6LUdbTqShE6EaRvx
fybG4l5Y+ysWu1cWVqQhMPW9+ph7JpZcv/QSelY1dczQWueW/ER4lDz0cChiuasF
heLcItdMOUT/g4Ns4orSbeDW4Am/8K687g5gEf1q5Y7zBTWuGvdYdUZ7A6Gmlj19
fLLcfSb3hI5mcqxUFIwZzAUetgP2sZzmBqFmpglWLKjmYMy/ovWiTajgd1qsO7px
JA+TlhS5c5Xb2gMvlQUR8ATUjU+wlvuClU41rtW7JmSP7eS4mVcFJ/ItGUg4TUu4
b6JuCEBldBW5BzJxLWXHcct6fVuo2Cb2/N6ldtV+TvcDJXhUWfVg+h+TMLZrtoDA
mYPX1338FwkPt9Ssi5vGH6IHEj1PrXa14cKek1D5FwVyttBr8YYkQ8X7Vsl3LTsS
IZ0bR2Fp6wG5dsOk5SEi4QWCEpSFETPoswOg7kFCDGKDn1khmp9jnX3aZJXoJpk1
468hgZBa4zL/4RShZYceDgYZgI//E9PCx1Xnhjgns8xrbRdZ8tmo/zxDXO5IkEkv
WaarEDs0iCo8aBl9tUdokWunqh/FQ/BGkynY9Xs67QEOAhGdJQ8rUq17HJelv7+P
EFpX0py4YqcmfeNxrGPf+o6k9RvWZCiztYIOtAFMpid6qMJKerrnmjFhdDw2R4kO
JtD6rRWMUSdz1s1iAowWNovGP1UcH/9HKtsT1sR20uEInO4fgg9Jw+RYlmFZySld
TUOIB8GSqmxlNsMhaSjV8+0TxnRV0YMEXVrYpVJxYt5Lkdo8PVPwCtHe9M6/T/p3
xdcyGThAug3JJo0GoNJZaiwZdPA7UknNhtVGUEmD2pmBUHORezoHxFkDyAfr8GM+
2ahY5YS7ifMxRl2wUy34sapeqlevdxsfiQur0cNIt65XDpMiQhu3pbeC6RUsrYtY
HZMH3cneu5DoroJPg8hxSVki8XqO8Eim/bJe/G/cNbQF+Qn5NdgJbRRK4SsZlby9
l0gLSd/BUPZYl5y0aH0Hnhy2b3JD5lSN5AGyBr64FlV/aWwUtT0UoWOERhYwuJGt
IkY67XF+h25HKW/hKWJThO4tUlKrJGfHA8denKA/jDgUqRbQ9v3ktYzylZ9bfdB7
woi2rEclVKg0OeBfWGnkTQOlObTAuqa4r2F+Pq/Rk+ZFo/4fuIz0BAICvFAkmqwk
pj5TF0KyGN1B6bjiW6u5CCjQhyIAkZp+UG7RvyHu7vKN6RMuCIZanPW2WuX71dFg
YNE4RY7zNUZchwnVNKtKZE4R4E/XuAV3+0l0h+dKgxrdgMGmfvrc4co2ER6BHYts
Z49vXyXf2jLYEhFYxrHKiR9tCJyM+zi+S794Of6TgukN+QvsdOPCGXyHbPne85mg
x+eWdVCqHAtVqInu1QchsxcHZEDVtizmM7oaka/GmHGILA9OY2Un25uiEnKWCxs2
4ZRqx8zKejTpZN0f1qeAV87JZYG32peljzoNtw1r8BDB1RDzlyFPO+SPtPr7URPQ
3i9C9Gy4yLq6Mews4Vm1KOHWgXK2uRQb7gXKxqp30knMNPE0UPLyyq9JWKDaH3hZ
ThUgLaqocOITr+9Zh8xJzc8G1rrOpKcXyaqaa0zAq5Ujlti5qFjRZnOSelm7rlB3
kQ6XuFs3ZToHVywWde4h+ofbNibX0bkjyBh+jQkI+MzuSq7mKxTUNInxP/JgZ3pq
bcasKU65+dZSZ44pF5qVYm1pQb4c2TzzcrTXjr7gxb4tFbamAKcO4lt5l2EGWkqc
08za7JusMeBJAbrXTVIqLPCF8M1bYxSlqn8HFomEiCqa6BKHBfE5XldhFvWtizj9
X2VbLVNdgHNTbBLMTyaeC1FFYI0KvgT3nv+fjbTefLeRlavVSRICvGeKf62bIjkS
HED46yUU+cRi6kjQkrjYSyMZoKkqJ0z8dlzgHq8y8xJ4f823Xe4zobph0Fn5oNtN
NY9AsbydFtYwaIQUmLGhjUSw8y9DCB3igNbHLaVSvreX49Th8p9mojSJqnsOxOKa
qQr62gB7bM1azfhxmsjH4YkKgwfLLYuTd4PfJbwfKwfmizfcGRKD2hA9ZpuYVTrN
OOu9UcjZCqvLO2Q2qsjDBSP/FkhjtAGCz4LmLNInxX4BcaWl4QkC4whPDZgqFt3J
iHpjKgXUE8x4s4F6xG2ZlmyOrQPHXZ7Xe9o91QdoBNqvNBYmhp9ba8pzgND+DJLm
n+n2GgvRb+qqj1N64/SnM+GaS7niVCQCMv8XWEIpztyVNTy6v7+MIiF47GBpp8I4
p8dNmWiIuPEMXfbYt5vAi5ech5Mfs+2BKXxIoMqMzU7TLf9NR3qP8033b2My0+82
oHXJgfJRlQ6QJfGS2dRQMYOLcVwXSki86EVpJlP9QhigZBJDZKmpCNovgZUJNryU
R4yHmLfDEbN5BjGzfCnXPyIaUd6KbKX2np4kYv6Jww7ZdhIPBkXFNcgVpqHXaDT8
FGfe226/gt7dM806wHo2yoPVm+wKtLezMjxWy5KuScJAdJPX+QocC1KgvIKCa3DE
f1ahi02BEuzGauRu53xeZIMhrcE/ENBEsqFZOQ+bE7jVpiPvhqW19dzxr+EzWbwa
20V+Rw6moeNIKa+WXoiN2gfaEaai1GlvTLpt7SeABAm2+aabNjXSZ4kbJvMyhypP
lpmhWizLSz9XfkT/d5Da2hIIzVDKF4L9I2JrDYnCRhDpS4RxKWGw9BiHJClEJVMs
9lvU70WLD9WY/1hn98fT2follMCh0aQGAGiKRsRGPE2ZjJ/rLbW7AywgJi7EGens
4yrExCJNtQQIFsnHPYgNzLrCddH/lVxvQPtuexOoew3q/SoJCzzNrB9XMJIT9sSK
4XCz31L+XqaA4/Brd0J3QeqZNf/QogEufnFZtTbP6+5N/HwjDa1264Vyy7MrHw4l
HVtco4jSGxVfwfPJSBApFlCMchcvwk5zKv8zW58NHoEzdGz0KQ3y62EFDV18csbL
oXrYU4TGACYaWg/yR27A4YDwpS22NrXxNCfTObM7qHqMwb90WWq6uPnR2psZQR3T
EhM9hUDzCNGH/eIDVvtyy9olXAEVNOYzAImJ4IPLjpCzbU8t7W2Oox87+lMSoZJH
I+rHs2pglISUsbd0XY59NlXtsnNy5jcd7KdHdQTKnLd82vfV5CsiGV1NBbQM6M/R
/wHS5CtFnV0WsXqpivzsLjJwwWrvoQLMmS5j7YL//itp3cJxbCLTpvMrazimrHoa
KN7vUZv7vosoI9hfMmI0jJQER0zc9bmE93OaGjlyytkIip9/AMT1TriXcL7fa1WU
Lejd4/nxbsa+6gVfexrTb3I4pIVXiX3BkibUxsWTINrjC+3hmjyQ4Qpf9SLXcrtB
r7jOXMPpVHvbsHfUbbl2URZ6lQviXhcUlhJUC1WJEXnQmwsdyuAyCeEzjtCZougS
kAiI/GOjERUiZjkGzBqfpuK4QWA+0Bgwb199MceNSIm5MOKfuMXra/u+GIDCIJRK
0pF6K62HXlkv7pFTRvv37JaZLhJWGI4EvA23OY5CwDFnyyajrkFCxHKS0gz8YNqC
B/gsG9oy/UWjxuVi/I5r4kUqTG28sACAfZ5QrVB5a/G+rBlubkNFXsLcIOn/qHav
Ar2D/ewJFw4Qh2d7TY9zqqZ0FP+VImNIJUkX9xjIoTx7oxWrpzMjB/5RGy1rdLCX
pqYG5Ql2EdnDH8LyxX/haciwU5Vap1ZAYIOxovcmf+kDDOX98a7l1gaj8hwhA3rf
PyL/dBoUSIa3LYO+U6XuXktNU75wKzACJo7qg3vGCTg79qHWWGbQoafATevHzic1
ImpWZ3acMQe3RqFyNwSMvv6sGLesWnHNlLWxtAPpYtQO2ZqBE54+bRXkC0Lg7lX+
9X8Ta7x24q5EkRH1qZHowmWnytrHGDI50Mvh43Qc3yx/6vmTb4egOnh7UWZIbyPt
vPEa/o0Hh2+ms5siDkismXnsqFLnX8B0dBylFqW0EhZCCF3eybY92niKU5k1Tw7U
XHgWJZnU49Yz+Tj40w2S3HkPXSI37kMf8P0z1HwlDWqY2M6c8zsvaZquWUjtTPIF
u8OB7HnqdQPNo8soP1jAsZoPq/1hYCV3QswqzMkxMuT/UMGfaXbKqh8V8swu1PUz
UBUHaUfCtVBw1sIi4ke19D6pQJs2vDCHS18+NWW9qmUZTKtz3bUyjp2w7qQtBu3y
XomkVvx2eW2Cj5MfKNg/bgcDcQwgYmYVQFacUOF7+cOABMnmXvezgo4bFv/QmPFi
rAwCBZGzcgLJJXja+vhwnxTKW9KVmLANHkebBwJbAnCrCyaKlqRYDRxxV+qrjxYC
snGT+0DRkJsMxH53raXsQW3CtCB9p6j6FLfFJ/lJj6HCKlH1dToMC7lo9cAnI1wP
QrAaIHx2FOjyr3WLHUOG3kA9+JXMZo7WdA2b5tlRw1CU6MDvS2/+GZpsPUstG9+l
Eeb+h3fMVR6FwMUdgMPF/kU6pGMdvRQwvdIWvzS+OmbR1fM75esh3AqF7kW+0/XS
ooi1H8vl7DECK/SOEuJrcUW7I3/TD3g6dU2jX5Bp/wmQSwRYlzcLb/ftjhxC8XT8
0YI7RR0W66eEZoKVhO3/rj/EZ64xwAk0hZxACU9RFaKe/kJ5dNXV7J1hJzDsmAjU
0SRbmpCGYrbLXkdBAyX8drJ9sEO6QhFnkANALTZmDp3NfS3zLneZwRFHBWhhacp9
kwpTMgOU7mlkLywoYzNVxF6qZK4n0r1IUF0Vcp2enFpB0x2RAp8pvnAylcu/0VYV
T3umtPIe36eeViWHjjzL0UaGhi7ntl0AoG2UEYpvjtSej9y2fdF7+YCb566rtS7P
tjR4HRn4ARV66FEN+5HFwpI9Gymq5qM+G9dSB4Mh5se6FFuh45F3Jd0upq00NQj3
Kvgn1NncFMe5CFF0lq/CNKMb5eogyTbseypggCcHFtNm1dayiiSocZ0R/0BsTEoE
nz5FlfrQeR3Vqs9nHxFiv9JsCa7/fGDJTk9QXTRVpNau5BoyjdnJMG66jlBssMgB
rzjU5kw6L26JeAI+8jssjZcyvRjzfI52qKf+PKj1rJPNEEOL78HlMbGDbJSQ5bZ3
fch2W7VAdVJb5APLdn68UZeOXzHAR5mGTnRaI5nlU9KBvFeEj7hzAxi6F2ZjvWC4
eo8WOcLEES97JeTOK1dKYfT4oWclULFM8pAkp8WUOChSX4Bx4K7LujM0h9QiRaeX
hSpYmEWevwrN8R71Z/skyEJroDQDTKfzCdotbpcMJcPZDoCHvDMkwx8MnPumstKn
uQ1UK9E2Vt+0NFKAS65XFczcK9M96CwSfA2ajDYtqdI9DfApzDs05q7EGEY3j+JB
3Iz8OvFCn7IUZ7IWXwYFNKTccnST2OSLXAi+C9fye4glTtu6YSUFgPJtLA6A2evY
laxNP4yOQVLEx/EcCd0HVi/dZmBg8pgWUL5VrHvU4xiq7gIJXdvec8i3rdyAz/6y
ogyRuuP9LtFSUEYVPingzamtXGXmRMk+ErF+UA6lrBIV7ZgZNOBgcpfgcyuwsp6I
nZOUL3jC9IgkRDYYgjTFjySvgn0nY37T0/49/uigQghP+1ldi93NBxaDtM4c8E0R
FeXQdjhgpc1zhmQp4gOZek5KmVufwMu77ALJHlBvD1k69cnqlyGVNbjYJVJ+xD4P
KogKlA1vS8owa9M5LLiu75lvekTwv0EsmN+UMDz9lXdzyFwDbFJfP0+zeM6LzXcv
lLeEXenIHP3fGKlpDV2ZhP8Qhvu0fbexWrvPg/o7J/wd7kxvlOm5jb+rqiXCVmvl
JK+E6KvZ0TYjJD4QjDtO+89EaRcGhboguW09DQAcZo8PUeOsDWarbZPjIcz/sJNg
kAeZSMkJwKVXikRfyZtXujo0roRNdwV8D9BdqZzW2ng2f5hr8zmddf6z/FDNfIUI
bB1kP1vpsP+WSlGMZBnmeN44odmA6EUyhrq8OwVw+wSpDwY/Vx7YkjAePxWxkw4L
E4Xd4m0jnfNMUy4JUSL+496qhbjSCrOYpzRv0AdskcQ1abuLZmFgzVChnZV427F0
kSwi6ngRFH1ooGh3ufpTh52C1OipbZZhNDwE5IyAcIwFDXmDNFRbpNOmwTCp9VHy
LiPrValILcFlbcq8hImAw8+XhYI1Z83HEoVo29ND9tJojKeJP6m0kl/xzvfxSPet
TGzJVvL+UGdICU94PtxUJMCTfHVNkV3NnFuHncrYfPsan+9XxLlCdtxLbscEsLIF
vlxBVSIj+Xttdw6c9yqUp8VVYu/GnY8rq9HpDMA3sbQ1B0MRu/6H4CROOLU1GC4e
ZD8O0xQJQY3S49SN+IsHQVHj9ouC50KLvb5ZA08z/p8LLC6/SakD/DYpSoooznJs
ewd0I6GARK2v0uAdPqUDfPvEulMFlWDOVaM5MpsW0I/q5ozZiiunxXlZzISkIgn6
lYYYtwGumDL9SWaElUiyxg1sGKuJUaK1XLjczNQjUQUeyXrB83YCqqHWWb8uE/3Z
D2w50GCaWPsHj3HQFPr6rslqtDOTnv4fvC5Ode1j/v92h9cZx72HOK7pMyiQ9r4d
nSTT4jC8LbegyaPGcVti4qAbMuzG1a7tCUvrxthqIrwlt8h3L+HLt+H93eGoqK9J
QUoc85V1qNmIy88LBs9kJLPcsBazLVfbKCpH1QX7bMtq0JRhgqy2h8bmsoBn3whX
rkq5mCMiWIC5Xc9qJrpRyiH8L+lqGh1V9ga9l/gF1pz22Wd0p5lFVLN4GG7Gx4Qm
QF0dhIOEt6jUMThzfGuBkmegkqHmuGzilGiCz76Xz4947HdrrfZY6NPKyWioLkOm
jndpknEYEe5HtAKyM5Aya1XPH3mE2F3tTN09qojJjy5cNksIJQ9uRBlroriMtmX1
Zih+nop2xBz6a3m/N01GqAbgbmP5s4Dp+LrNDqaq/lSzdvt/pHU8dENso5ZOLMU0
pcPjFpFfKAk/1mo9JxG2XZKx7IIhXQjQDnAhfWgQUB/5aXqsu6zzIeU7YBlCnxQM
C00NQHdpwGtWBxWCKwKYU0GqFiSbEba2MmoX2Q4y/NOLGGBFYDOVO6Xi7/scM1A3
eU7Dcxcc6uV5NLdIpDH2BGoODfMr0GX6P13/d8WWYWPCUJSkgwz/krAxfGCP4CLN
o8fzUXooIebTZ44N9lg3tqLptc6eJ4/0J9Orw7lrw7b8KAgijODSZtHzn782KLsf
l07D9Xa4dW8xPTILFqjgyq3oUwghU/1fapyxww/jWAVv7E6PSNNXbh0o9RT9tzWQ
C6ljOJziqwqhhPw5ZHatMrNEPjl+n63GzXKvdMsJ749ajw9NJkMmwFgVZHGoOi0m
MvVl48gXEml3B9+95kCN0cJvSap7BvQLU/K1NuYyrmVNikWyqd0sREPFin/hDa/9
mhGfC3cNRK00yA2knsvoUNcNMQu5Z9NvVo7bST8+BQ/7tRSuxDmVuV4rIeq6auas
QLOWtpYpCGRMSvOZZhHAxp3JOqFkShAIgV5ARQTCvhDuWiI2c90UfYboYQCExN6M
UJpPBStG0gbC0ftKaGvBShgpUIbxCJpNyaYi0DuZnb6KDfZdQprebjeGZ+hRGtC+
ojwOpHRlMH6S0wN2JjYQC3SwHF4XbfBbs2RmPz7DLZP4jQoVGTE4mww61FVKNQPd
iORPxGqJr96uEzHQtXLtY5st8a80jZX2e+qZVtBmo14x7a3qhBGK/KzMfSwdmU/Z
/+iBPUqaVCBt+LGJH9u3oNbqhQy9UUXffN86n2rZy574zlNQUgctw4/r6UHfYfy8
scTTp+Z/J+C+f/N28WutUdzmX4O5+5X61DoKxtFtxkcNn9OxytJ5DxpDmUdpkBgr
BfYxhvJ9XhTmmXkko9y5xU63oFQqqerscOFnnq0T1AsBhV+MTFb9baPhixvjJ/9Y
5EcDNqA9Le6Iygx6/JcuGc8qxtErtzZV0q56VmtP5KH223gMK6MeZI9emE+LBK9r
wU1lg5VZsuLu/j1WB5Y8MInLF2S+1VNDURWAn13c6JEmlHF80LDAPbfSqje1tb/G
rqs2CC4V6MvErhUvsspHloJUc5iHGQciJvvJN1fv0b4D703rNafr9irPEMEOY9j1
BeFDYcdCE+21DA/1frxpfSUWo25grBiU+BrqvuVyw7Ly1U8uX5eeXTKIKZgy7o1g
EUh8GOrj3QzQl+42En8lj7oYwfbsqzrLKRqsOZ+/b395//b9KvvfkF8xg831g0ar
S67IfK5Y3AyzCEgWcHpQfrqaahWTyv2cPFfIonjO7fcBiYW3MqYZi4jpYIjgS5zc
HGCaxskPVgkrCCm+JGxo+ZxVtyh/eFpg9jtZaCNN1wMSNEp/ZYOa2geVtPLiyG7u
WgWSj+/N/t2Rn1uVBA+EST9M01o4yJeYDZCa/eHTJ6NvImg6K+R/Lq4Sbf/xQRc9
jwnOX4XSyUNzpdizHI6qIIxzcmzpuGFZyOfE7QV/3nXI4xkk8tGXtydYBchTuEFW
C8sGEEjmi8hNiVpCYkPa4yIXnXFJUaTbLEiDs/+Asuqy1rQSWhhsYxM/PnjpmcsH
cF3myyRiiCUL6Lre43XmmhpK2Kv6WCX/rShjGCM84G8Zq0PjyWrPNhbbx6sbwhBg
HbdfgGYaohw4QKDPHOYLgaleBst/b7jgdSTNzmDca/caSAs3j58OEn3oDKWeGm/O
pQGgtBGrQa9tQmGkNDGAX+scRE870AS9Urz7f+I8R5nx8h5H7B9X411vQFDB9NBm
wds1JMDft1YmIR/48rpS7qI7KsftomT2O3J4tEmuWy6Fr5j4XW+MFo7xDLOtdOVt
C0leaZV9XWmddmrXLp35wzLNwCFAobvB0daoBqxMLmbxsSzGqnD3qQg6QT1eUKal
uLsyqdRukguELaLUgjdD1gcjCO2PaM6J8WOzA81+h8AxBHnieleEIo8tUbDw8CNw
7kwWBZRPMu7hCrEO70nfmSLGdviLdGCUY50c8ELYlz7Hevj3CTKFhmKZ71/MVicG
scczimuuDBJCnwZnYoIPfI1FJ8q9c8Hz4QSTwdar4+EWscInRUXwbT0tDNCDnEtn
fCkL9i16UuRHn7dwwlzLC3S3J0LslDP9wWwPs+hLtIEd405buj5jhXwBSYcjNY9J
Fsf7mMhnpVmETKmy3/JguRmhsExoXs7OrjUvUHM6R/Zmm61WHCn0x5hPlKZ9iofp
n+LHaOsyD+mtGThily36FMds00DD3zm7HWxjnqAM9iQtJxwD8o7qRWHAwwTlbEcO
7/naLQ+lAkEeK1rWWIX+VbJw0kAYkv5pRNVeXgNDcNe+hNP4SfBAVGWq5S3+/Ons
7k7oHQ4gKpdbFDqZFk7p/01ETKZ29w7cUr9KMyS0x7vMWsEWnkITPr/F8QiiGuiB
0SrSex07PHhaFpP3jZ3zN5Q7s2wuq5afQXuGOfox7COgaJDx+qTpIoUB/vPPeF9s
AOY0keswUg4T/5CeHU+F2pyPXhhkGejkUHFzNQsTm7zJTvPgZOS+hgSzwG6ZC69j
Tc1ZvRNlZlhqpfwFJLcUEzgtrqXA6lt9yRIlgQjiakRK3TU8drbt1FHIqVZSaGYR
73puK9kQ2zKtscqYgUj30B2cM/VjQrebyxkGNA+sXvHq6ryD8mDEiHYdlNo7dTd4
RS6Bq97p4tmyHai/2yR6YUJ5Ftpar8vLPRuPYBLLq89ry/hCW+OxQmjZPgf+J2K9
98RwNNumBpZo301lrD46b9Xs4Fh13con1hQW94yQdAKpiNPdBtublM+8zALLNMr8
TcrJ0eUepcMg8pH23i15hQiih8nfaEj9GLYCTZApAdA3udFHcqz0UvffY5P229H1
sr5JEfKoedHB5/mq8L5eRR+BJCUQHkRfZ9SOEkEPuPY2FhyWAJG7LBw020dps0fO
hVzpnl/F5QnpblFzzAz9Y4Ubk5e8BBtcxkRlYK5UCxGDNs0B1di4rdI7d5y2FIg+
5xdxTETIEYLKHuYls8j6WZ9fg9xe6rRPZkV56qF7ogbtr/k86EhqnJ5qnw7CSxcL
xaqWDNqVq0lnILkYdwh9npWyKcZ9NBnfiGjHddsmYSytK9R9xuzl1owia71MebOZ
Z4JE+PYgYTZrAWrMXVIHV+KmUs2BPG0CnRrw/4ufrjdK9C65et1qK1AEfhv2LQnZ
Vojcc6l/spRqPWJibrJ96pjcPMDMXRwT1YqffiGNOy5DtlfMv/rKSfaPulJQa/Pc
IGYsFVxAhykLRMbXBVVBv8a4vcD+fqDnTMfK/RPrBzv1HZT7/tKZhVToRHYAdO36
9jdXF6PiIeGbQV9mLSW5Ftiif7E9HW0BkA9sYCpNsq5rSr9hY9ZQSNFWFLBLfoAn
cDBkDzVV96Zsa9/RzxDZPcvWZ1MjWx+p3iQywSACV4kqYszQ6RU6u/LtB58+xK/Q
OgTaQll0tz4pabfaoPglhs+2HK05QWlnYiO9NqiVLNSgaazVtzXVHwKSi6vgpViM
Q2H54ZOFZtxA7CpcJcyuvlmALHWYKMaYaovrJPsQ5xYp8WktWg5CHMN/fZEVg8vu
N645JIfulCGwzVS64efqgtkT7MDesygXSbKdXjgxos4LpS5rKS6kUROnlY9fvryR
RACqoPvRJnGdAh5S65qvoUwhxqqaLgcR5wtuK/dol8J/brVuZB/52KUq/952OHzs
gh86LMfr3Jt8x9paoXHPMjLg+p3aIOMIzy24oOceHCO7jiWkorPSaJ6YViGRBRvi
RdI+s+uVpSjaVxBjXlDo/CXsm2fYI4l6uqS++SCaOpZklzbjiV7FjebgQaelcuXP
WlK+GHUjOdl+BNwWQR/du0iopZosQ0pTYWaRrUFSCruHIRzEc/R58jshxkxty47G
vn7M3lqZR64tPAyXHoyPgWkgs70t++YAWIOl/JAcYRdV8Om8xhkazWBKzwO6PBSb
pJ62p4r4f8dGWS8Mp5WSYA2A9OoAGIarTNV5k72WnuFO1yCYMbxw3XJYbPF9JeZN
72VqDRvHEUUsMCvMlfFX6dbjALuFcUs0RYeLFgtQTr89XqeMH4Vnkz4Y5HpZrlEz
TtAfLVYYL+V8bjg/waV3jy+FswKKrEssFOekEhpcMpDJnxcDsGyDvJgavzC2zUFH
3Rlt1fKKiCBeffRQmeKks6JP5xSmDzn2OCJdqQCMzASsH5N8IAlFmZXfWdt6H597
b+4uie4WUCt4d09g2PZO35OyX+Rt9thQYO+in4uqcl918+rz/WUkVnKJdclaJtRh
7ygD1+4zuUEYteWKPw8BtBSWW9a21zkbCqDrNoJoOlFpALvV1r1PNlcpG3dD8zIR
IHG8DAKUDIyUwng4z9mBMwrewrvkVTvq2rBMdit9Dg+4hcEwfYIILeu5zBGwtwsN
pOA3xucCBkJzoAS7134SLQ98kQ0yC9nvtNWkzJsEO2o+742o4RzgbL2p4oarxpx6
MjA0JzYmNiVF+mPDh9p/opO3nKtJ0VnzLe60/topIpo2W43qieBXyT8WisSWSsa4
SJ/TXvZ3wlqoWpAVE28/WgcGRlITJsALZgCVgpqPe5j9eScb0BQF8QghcwkwotbK
KBRIoRaqBYISUOCBJuobTltObE2Z2hHjVc5SZLs2Gkjh1g5yC50aHJ1x6qmrTem3
gt2Q+INr2TkKSzggsl/azYtBo9pp2VhGVmDD4uojAldJbJvQ2UvVqWCgwW1jVjF3
ZjtfQ1n0oWPvanmPzTCAwtL1YVNI13XZeP+zUPuMd7AabhG94KytEYEF0158rJSn
VTu1rL+9KYucLKbJRQpsNjhGI9jWXhSM/2sw9Bgb9gKwLUIPqt54R4hymUYG062v
4RAcvX1EgIxmVc6nDd18/s6Fm/rQ3pvDULKuHx3sNvF0fX40gxYy1Jagf3kpxntl
PoudwsATzCorCZm2+cVvk+u5X++ULeLuNtNDYxRka8oERFNMUlGMFKrt361eOa8e
2aFdBPA0HxmjHdk9VVLJX5DN5n/edfZqYoDDiLXXaD4V4j1YTWZPRswKYtQyABqY
QGoMD1ONCTc1RicanetDIwU0sDvVfqkz0lb9q65K803br2zAY4WJdBtAXZp8MoTV
9l76djfOe4qsXwdeCFuOazX8m2NyeKITdv7vhsHUmM+KKKremAYwEsZR41gyPcDJ
uAmgZuWpCWPpmnk9i9lMfaGzHopG5ucC7LGCNq/xPzuxcJoglGykj6l7tFFeeYAu
cB31iwHSb+EYtC4YWK2dFROlrvuSu9zXb4JvNNstD0VVttRtUs1xsCPZHWJs2vUp
dWCfl8mW5PRo5qAFpSuXvSkKBKOAxc4a/Zpg69qIPLqdF5OdsLHfKUHbUrnbiM1T
YhYSuzn9rZo8zbqS8ea+v/7y2iq9aTltLQ68irr/Fnur2TS8YU8awoEx66TAEywe
ZnUjIYonR4u2JEPZZZFwxIZQCWvmTcT6yl8dptrwsAekeX0TCOnw+XCeCqtli9/y
Ku8rY8x+btdVKTKr4INeFAfDfB8sd0U6OKWcFIhP1NoSRofLe9PbZTWFcMzj7NQj
txf1TbajOBgwy4j4v5d68Hn+8p5O/G9gTCmsVlzhAPvX7cY3d9Rx6vDxPZLw2cmC
O5rN9mmGZ2/hhKgA8088a2zzKk5ttZS6nO2nJYQAWrlZUBQ5Wq77AJnqJr0a8XPA
q4++plNNLbqt4rVM0YhIfe7h7XyTooCFmkJTUBO172lbNNbC2aVfpQXd61OwK1Xc
3ZxPR6e3XE6TV0PCQFvObCR6hjQl+SiQIy0I6QQMEA84YRcqun4GQsbWBY2OBghZ
gsOUZ8A/XnzexEh0pCGd5WV8WQiWOqxQ4vwdiy63i51P6WX4DPveqzRPzlacYTt6
vAJ6GDxLyf64f6inQNLq6ZW01zlg1iIJSogBDQtBtxAKh9fz0DyoegqbQJQt4yMd
sKotkRJSlQhwp0+msxUCx0b4nRPThKBrh3+ks0WI0+L9TLGq3i6TEHKKMJeyCCN5
qoVyVklBL8mzmjghUNmO/nsQ+X7HjH3RobzYcjUxxxgAr10E4jex3SQP1CQLrRsh
kTSOac8hcmVUhy+E6drhwf1Kc9FQas7ubKl1rCtpHp8v8djTyJxNEzedf4KfWMyC
dlTzRNcSapZkSTBOTTDEL/q7yS45+5I0oEBSfLWLdmtJ5SRHQKbWGOSC2KFiy9iX
Q8xv7zzELw/MqO2LoOHWQveMYOu7jvjHY39mc6cbZD+EY71GqD1KGBzHDvMcbDFA
0a6e3RgwrKmv1WtMgq/MAa9ekBM3SDEdlG9LjoQgEiVNE5znEI3meouGfyDEvkZW
gyXSQ3grhojQmcqjs9r2GAAa5bkqOWJPerCpbDgQF/T/+ixu2z2oUlwfyJN9Auq9
oVGnLEdPL83EDQcS6Uc/fnHhVsbUOT/Q1YRyEp9ptFu/ULb+ZiIxAOyM1RsNyf2R
t2a+bwobt3t3Loc3B7wzCCwAIr5PYDHOVL1wy/F1vSvKoeGH/vNRKZmKvzVVYPDv
aP76lkgEplyOsN5YTfm84nFWy9z8hNTa6U95rPxLKVGTUucGaqQ0CEa1aLQP2w49
g+CiqWH4W/9Ibwa1nuFRG+HvGEtHjPcEyJONHjMl+/CbAukeoIzpSZtXXDZUDxdH
q1mLQFjDayib1yNMgq+l+uZMmgSiXFA4nXs2IZT7/FKpL6Fl7htN9bl6hm/Egw6z
7YTxqFL4/eST2iP0GMYV+c3/WJwVOhNW2OwZEVdqxyLwPR9K4RdS9SHRBFGbh5AJ
JOYlZ448OSm6/sI8OQb3sz8nK7/uwANi1dxsvAJiWAoVSVhzQBKF3y8t2wtIvkXc
2Ol105dM62IxTSU3IfHEg0E7sd6tHVgEHE2s3XtpxmxgaPddbyqPYOC0vEx7Fk3I
WO5TQmz811R1zml+wyhkmQrxrLr6dctu7lH6bm5oYpIgxklzofj0ENADumRyEnzp
tZV3g66eoxx0HfirOikMVZA5c0qUNHGGXzUfuJCBJ6HhvftGSARsAyTSMcZX0JhT
I18yvCmGLIjEw5ws1yCVc0wCqDyVtBbbqPruQlclsi01hKWM5Bkh+am6a4jDUepR
wQAqYochOQVvVIAqjgMIZG8AGodWR2JL7M10Ezk3CZ3dTeD6CzgFIq60giFaJ1IV
WCZd1rQRHN6+JFdK42B1S3/XOmf4dPCnZB0sV18QlTa15JdbkfBsQZ33sxlQcjTB
z8HTuljfD3E+usltgGAoOOSfGC9j+DqBpRwtWpFFgbICGgZHSj6gwRd2uu47kALN
GDyG7BfuorBPigjf0sxWMcclbls7NeshxOVGjlSxpV+NTYkt1omIfas/Q4CjW9qK
LhqKeA6Bv3UUuuqr40ta5Y3lfpqELahCuhMH+fl1/Rm97JYVEE0v1RSiXhKHqH90
xymZNC9oDwQYkeIsC58RgjckBrJBv69x/xTax1WdXPVzCSCsLsIwkD5asAPfW8Xu
lDRkQanVchpNa7PyFYjS+g9g965Se9N1WddzBWitYVt8sBjUpAHV7W/GBlfMLWZK
NOByUiRplbeEaG1vnBf0UaRezKeJmdSP5rqNCeJLsR62eJ91gHDyFis6862xkrs+
VwbohyPbW8FMs3icAp1KiT8opNW+KeZS+0Q0xsyypYRn1dSDjJEzCgV4QMCeZK0O
soCeCKH0Eiz88RdhTc254lq0AVtdodpILuJXLsWCXe7WPQ2NDFl7GqNT9MDZfi3N
FY5n6ip0X/Jrdt1L1ZNMktVRYcFVRG/pf1eA7JcBTqQQ/rfgY3I7ySV99KBofRXu
JaSxYDtVJwt2mq3/TfYEBUzDR66Ybl9Q2+okSbHNChdYQiFHlG/yGtv+cyM6rbnJ
oRHXaHw1QGjqbDXm5rD/N67qYPeof29LtzK0YrEgfgkJanBoWI/OMMHfQpxzgoUW
E1JD4IzUABdRnw135qSe6AY4oa1wJv/j4IlqBLgplvEgTczIWNFYAO816YCfvg7R
5MJ8vYaMWTTmAcLuFYuxGRxnYvgB2jYWwUzmfc4SLBEbfBSuH9hMm+6yhSFVAusv
LN9V8XD66pM3ZbpvAceSuJmQt/L9NUVc2NUv3umGK+SLv9IulgTRa07NpKl4kRzn
KKoDancc3PXzo3S6AS1WRjma59VsmHDvUsMuIPF/lBFSLZifgk7nfzUfEoXBxiwX
dp3vudeH4iM+n0uNeDsTrD4s63VFiYse9z4hEfVxdg2Y0ERGHRD9gt284iGHAjjn
+3wErOW7b4WeTFlCDnaWWU9FvJ/0Er8FWHPO+hrPZHZbSWnJBiGE8TZbnNHlDWat
l6VoceNLdO9Q1iuG6tyn/EPDTG1I1wOJXvruNjORiUG8qYIMarpXLYvzHzZ3QOmn
IoxwOzviMP6Oc46qmAj5Omn+cmH74RWCM9a/4M1wZEFeS088PS1zPfUMDB13S04h
ooX7mj+NveoFLU+7fwZzGbtVr5JLOvc6/oy9FqUOYWalcSoAlKge9U3GlhJ7kXzh
+n8XEot97moa4eN958H5IwZbL4uiYwi4/haQTirnDFdrnILUDrZtx4OxwOlbtY4A
IISh4GQ1oZ56+y3+pU+81XBB6dU9B0AXFL8UwAJmvsEi65cyHOvac0ohwhnaiNQJ
YVkiNecio0wWYDWWQUKxfheCMvcR4TXBqFF8/8POPUWYsqBmUIY4bT587EV+FzKL
48JHSWrM2VdEpjq8CA6L3jsy4rQlnDUUy3d3h+50MKh/XPkN8w+N0IRNKZSD5Vgk
azcTpsyUQ35DasuCUSXzClJylQV+NHQNjYlJmrordwWY4sr+Ub7hMmfsS0D8x8n9
HFKthgWLwnqzBfFoRpa7BVTsHvqvZMjMsWOK5j0eyF/mX9eGM1Iy3Qv2rgI/GtRt
pE4ZmM7rq/4MY+73g7yGCtHjpsufTadhzVMPh0oawJ+6S3dj4wRd9GlrSC6uM2h6
ZtrvvspdPZjM2VQKVWewpeRpvJ6B6HrWKicUdq0MNWQ2R7jQPknbe4oQ8ZzaaObT
9Y3AbRifd2uk2/Q9Qcr2PejU0+JcKXS3ktYIIOG65bqldc6jnHPlS1nJNMHZm9cb
U7yC7ha4EwsCTJNMqN3jSc7KGrnV59sVFolDKZCWEzfcFx1rU+13Cf054f74TID5
ubsK+7hPuiu6l/DzN7EOqcfw8Hm9U3uMOc1kjjYhHrxxOfWsYR86K8F7crsvThEu
4lsFGkModzvIvZ4rEOmAVD9LqpxMguyUFbzZeIoMZ0WDVwTIkal1nhEPQwekqoGl
zaNpT3d19bQWi/8Z9mIslIvVVVpNt1KIEImI17yNkzU9A7R77q2w7OrjXB46mGlm
JCgjFg7reDeyb0viOKn8uXe9VYzcgWFIExuYea3YuuDz45WBcqS0MshxZEYcAZ73
P6Gq8TVta3hQx/zY32sQxk9R+gdVDNFmLLbhHJQiymNLx9Iw3jOwK6vd4s+LKMzT
CaZvlWOaGOwcJDhOHWzDyRnMKOtfACqNJU7lm/hO1V7v3HOgb6K5VVy/1sDIAond
UPFPWirN4wtqKs8KtT1Trc7j7BfowQkAnpBILqh/DyIwA78x4rpEdzG/NfE3/WJ3
1DMPOk5uN5FrKChIW4tRMpu5MDg6YuglosfBsGIXyXWTB+AmWRkGOrJI/Mn+9jT2
mehyM9+3cfSLHlxU2sdbC3Tn6sa0LyGUfLNC1/+2UTjvirV4PeVYeMaFejOcRCf7
A3Z3b76sDKkdynk1J4ofW6Sf0HgVV4ZqrseN6nQuSMmSYmhApeHhCFlXAAnX96OK
NJqomtPA4Dz7ZBn0IQ9AVf+BhRTCzOpuYz4yRBTl6sLhoyx01+uF0AxvA4ZhDjD/
7LA4B5Jygby08O5ijX7S/+s+IsRX4QPh632z0mMVPdkXZfjk03y4dW6uIicfCMs2
pFHYmPStq1z3oKW3V5Qz0Cp1tcbeyfm11PW2ts7F7jPoPaBwIsGJe4YPeLb7og07
rN45rkxqjpnzHYZat95dUvUg/s2l0MLlwst/q+REbPoF0sLnBS4dLMQIkFSwu1cQ
d5eewGtX5ioEZ3ipbY7wmxyMbSmIL8hqQIAAb8fQr8w9gija2Cn3tK+u3JzlnS6n
Uqz4zUQHI0gpFD3LKzCCo3AtjqIFr6bkTfx/FBMGjXmahiqyB0aB2faHSBFM45AB
y0WFVmmU5HY6+OxVdVc1KOUQ6NbzAr3h3uCW3FR4vqOdt+3zBmUkxRElyhRfKfHZ
st2qedN/so3/sbzUPGKZLLJcfoAWfsk8sJqdIdyGFLOaH3aXzurL2Jj0lJjXwpQA
PRocFo28Q6muDCytESJZp8wlKt2jMJsYIKl4Eh5B5IT31i3zaw6EUilb6Aadl/jX
MlTuavSARcODvGkaebD4+ePiH6yxuvoOxvPCJBTBgwPzSJDXOrIyvf/VQTLbe4G4
E+Tei4+01KEhzIbuZcZWLJVtz2Dt+62szryTTau0boOi7HQJ2vAoFiWiO8BtsslV
EL2gOsp5w53LlpdIN5Drf/14CLME7Bzg2EBiLBPHsL9y1MviN5ujW3r9t5qVBmJo
tBuXKnD4lFmdU3+Mx+/bO01ptuOQFQ5tdOPI0BNH4HI3rxxF5KbdlgPkiEhw6bVv
NXHT7p8BHZTJcg9T4CLNTYjCcsrQxOKsvDuVNjk/6CKkCn+AiX4I6c3BOujYVv92
K6OL/NjgfFnt6tndjQvqSR9XQauqTYdXE3eTZv87Ts+kIUEsTTNQOdMru0sQqyz+
9WLyRn0rxMdUpKKVjMC7eqUpYD2jxrG8xoqWggygoBEwXlb3YalkVdbFEBz3WoJu
8ReVAnlmUfhQs+ioNqYkKe5tGeCGEpk8dejuSXIGqiYRXW2d0nBlqyyyL6ybr+eu
H6Ll3WsBGCBRj7/YZC4qi381Nvgis12Q1Ge5SA94g29FOBCUCEGUU/WdTzCzjA6G
NEDtT664vIU1SI9mytWvCyrC9hNkWgRqRXf/scUxA1TM9qGlQZSVnUyRp+jNu5zg
8zPf4x50Ve2fisdx/EJ3wddB0rzvwhjzJBiVZcO4hg3cEKYd0dB8/8DX0/FVypKx
ak9N2OFS/0wSC40047LVmHnTP6bc3ZzSEf5pC5a5pUjuqo5AHaQBS3SjjHhwWj4t
ExP+pozDLvFOSoUoSvCHmMdIdFYeG16JTUU6QC6JylH9qKJ3UuKhV5q5sOw2Lgtn
SHDVxy5tyOkOLXNtMT2YcgOk7iZag9ghs8ixBazX2AWLoyKvJNvUHHVdqlwRkBau
z4e3OiKl6R8SFH2l4T4+acFCBBLGDByet+2n78AZ/T2AY5q4nfdpoc0xRMM8DFRe
G0KhiyQUBHnSedVKTs2gAAewM399ZA9ibFivxqqNmmH75dD1NjxjJNQPeCHStojR
YJsYlggdhQLXZR8EE6VWWl+bBLz6neRLCI1IKFbrqRwJkLhL6SXDOCN+OOv9CHdG
nEwZOAvPq5c2+d/8MEBiXpnLmowyqkFd2zGaAy3GiRw7QUYA9cULuMdSxeifyAbr
v3ZzB6zZsSnWSg58eMvEkX/x1ZMZ00b46m4CclnmJtXeXVEcANNZefCIKN7LFChZ
x35YdCrLWT7xKXvk7kv0PfhuOlSAcXuHNyr+gYPUtEGWrwz4GaAfu5uDb3umwo1S
GN5TYJDrHXyUPlW7lCChX87yI6LqvBXWWQVpSkAdGKzLik+cgxBZHYb4pSZn5yu5
P8Hxx8zl62CRpf0gWy6wtVvB4O9l4PDETRDMKao/yzL+H+9JQlvbvnTrT3IxOD5F
DfDfCU6LMu0F5QyvWFRFxIBKaNubyp+EU9tZdhx2lGC97UVpnFTcKlyJ2bzeE+wZ
v1M2O1cxPITyS2D+YnQqUDPOFP5+RM+Us3030e1a+wTacEotcpDO8FXkC4mHioGr
Tlc7lXLj1o671+rk1IEvoTGLHjM+R768C+h2xGkNS8zEHPe+KC7oYh6tCQsd9n9/
fBHN/+YIy27nqn9RetV/Ynr3I/ALCSjlLkMg+r4tGN2qMZXCdKa0jUUgCiweGFmL
ZCYPnZVJTslrxAgUYqtrMPLlwcWzETihyFL2YECzofI8XJgJAs02VEx0H0u0pjYm
8jh08H6tASLwRerc9kj3WUHJ6wttfUsAO+LX0JTBO9w34MGTNzRLEodAKru6ylul
OgnqryR5QWkSxcLUJSrFfeOejLdBBl7CKpyMlWHMZLNbIVrEzLx8tPEZrsCL4WK+
fgZEwI6lFPENa3cm0cEh+40hs/oOR1/eCMwlTeT1sIgSSDzpjbgOgMhjLGcBpStW
nUVtDANA0nvJptR5mMOfngboTwMrLHmvWtFJ0kHXHkp6C+IrpPeLIyyafurnsqk3
0esuv1+x5rwv3xEVX+ennVHBREgZxNKALDsMnE+k6zKVlwiS14jwqE9Er+LaeNT1
s9+X7yErEn5lLq0iNaZo1DG5tueT5U8oPjr/T6LzMz+q/vKGqnmJTaB2fiy2VRlW
XkyXpnmZa5SFXTbH3Q8zzc37Nuj5J5SCcgXGAjNGyZwQcmzIkevjK911+gIOOrBP
8qdxS3zgv5HQDgXFrGPxCUYe5s2jRa8IzVAgi2AF4o6HRYxZXdA+YYSfQSMcX/Ku
O8TslyyBL/b5237OicoCJ2lINUPbFUUqoWibXBK9GU6J/L+xiwBNoPGLUKpD3YTR
gNaPkhWM/LSvhzvFqUVakmOI3R9dTaH9o79c68zYzuqOsbpTZ0zjwk6WSohPZFMq
NDpW0+WWDqY0zUWW4kwf9tftr7QkwPuEMl0mcGi/j3xHXa9Nblxxg9Z0+fySURrZ
EFv1vhb/v3sE+EhX+92yGxDpEL5r8l1pfqKXbeFjRIP+0UMBncYLhg5z2waSqeoP
hviWIFg5ER34IT8FukKUsBbAXBAzZ26YRpAS/d/8BLQ4aa1awOkUFaHkRXYIJ5Em
q1D1irWfEapqSoImVLVp+kGM9qXQsKIweUYm/tRQbQk515cGaRN8RxaZ9vxnkoe5
UtCCRb3HXmc2e45YPgt3c65C96UjXFHdYWMCnO3Ll/2DkRfLI2gzltQAjxIvKry1
ddqggvzVfflC6jNHAUNNsN/NlLD2ny0auSt9cfqBBnLWXgppoMX89mXRuVCELNaI
g4n0cANs2/m59ZtJ8cgFaYdHJTTsZdEokgWYzBS6ocCjShcpwOMaziHXEkadtnhA
X++u8Er+FXZ7+NZ0UhKC3RO6AGnlEmztSAEEu6nc+uhaAT4qu0tbcKYMRXt9EHNa
gU68rT0wMX5+IQfkPYJRVPZIxvJUu85CJhGbCQnPXmkbbFpUkm5bG31ahgf9Wmfg
E9duJGLn6LbapktCaW0h0ogU6TKojHYz39jGkpHSPMaAzltRYAqiOg6oYNM5mVEz
5ouALDVSj5IKvhFgGqaSeBNbsLa2mh9Ww/PL6b3XHri3cFWc1QU0wo2t6prpwiMj
DtJTlQxhuCw6RdJYkKS6RLdX1BFDDEAwQCRGGgL70p9MxMgJ0UTI1h26E1UzEpQx
OMSTnb7/vgA9g4KE1KtW/atzvSM8V+8Fo7nX0/Gk5FdalLsi74hnnIE9XudP93B3
I8SlQOCiWV/8pQj+/tOFXXdiiBOJhea73kgLn+MXXAkS3i9A3Oy4cSAwUBzXIT3w
HcGUFC1IjOW86/XjbEv2k3CT7XVg5NcGC8rkoffpCdhPa0Q3zuerMu5dKao5vZ30
AKtPlCd3QP6AXCQV4rrdBl2R1+2ANafy+/c6ZWpval8YOW0vxAyeEsQFVt1c6WNG
8dOzb7fC3/GEwov+eCoEhjwvLCxtBXvGwd0jl0pBSvStP0KMz87XOlc6gTjKM8eu
QFZmvlzkQrAEyvI7mH/oeHONbByKsffqkmq+A3vIj/AIwk4YhejkCt7WvYnk/fXC
cArw7Q0+gFb+wtjcV6jOGNnx3z3n41SPCKAzHraCYAMnU/wRIwtk0JoR/SycGuXl
RacKECrg/00yWCmB5uG/FGDwjzf+iAob6bEDh8oPtNHkgKF1EMe2LiitU45ahEQF
oteqSyKqmYDEfOyjgxkHKl3nNj2beW9tAfD7yEzp+XSg9i6gQQ0U0ebO0iSzDTZC
wpg/Zp96RvoMnlE2gOAubMezNXv5duypjsv10ZMVyWYIYF2DgHf2T5RkeNsiMVJe
xGcEfYWs5DJA+NkX+mXhbEb6VJEeZWJk3xakkWNZFoQfgFFLacOEznk0GQMrfW3j
a2Zym6nIp0hypZ7wMwD+zkMqdu/jkpbY3I4DMaZUTZDIZ+XDVWk+0RT62Nwuqo7b
JnYXyjWd86UHT8+kTdfBq+RuKMybNNVKwaL2I0i6F37i6cGEM+02EgBU0hMEM5j3
R7IMdt5hxsBp3foGxnfAPcaCwqypm3P5tjwbjtNwFCwgbU6EPrIabGKyP9JaxJzO
LxZ3LLGaDKLPJBZa/K+ANXHe4oJbgIwyJGszmmueUP/JLlWz7ZmZXBJJtLVzyZay
FkFd+OncYJUsNNY8vo4wMLi8TPpCzOa5Aw1Ha6hnR6KKtikCVxU2KqcIaZxc6j5l
/lEhsKeb0lhh5Fo7ZoGoyk0K1/kEOlcT5+JvFsgxd/09Ef+Lt1d2mLSCYsQgZTVe
ssRRTVQxqCuYPCZgF9s1kD6Ew2ELutADh5+AgjSeuxLE+W0qrC4ZRyFVqO/u4Pvk
x6zSv5cQL9LtYBqYscBWZiZgX7IEeUuOhUPRWVYONewr/CgyaO13FHtnI+nxlS0S
6WUbMaakwFMo5T/hfqM919Ak5JdBk+RiHbx4JBMRiF+pPIbk0IT5XxH5EKoo8rA9
Cd/o6EcjT9FjaOOu2xudOwoG7gHnralrZztjlw90xGylpPrRLLFcN1xesbPoPrZ0
BRWyTBd8wzVBpBgdOh1XcJWh9mJz9CcvCOJ2sA0z73uslnbZy7tcwwaZ+gpOXOEn
v65V8pgD9Y3X9BPddCj4ivTYZUALnNeKMfvFbRvGYiCV5S/iuVUii9AWDaxuOG3n
c006WU35SV3qHaDJVmg6nody5zen1CXwJe2F/Y3qNdKh7ZvRv0xyCPa4mFO/I00m
0pJvZsuv981nMfGyewM481SPkMA2oR6eFy3hd3GvDS5rhFlql6slX/E2hbsfaSW6
n9hTc+g04ENjyIygitSGQRADhdNSuh7gzphL/CzQFLPGPdJgnzcVv4kT9e2chqC1
qxwr9ggt64TO9hZNdj488teY1rNcLSBFlLNknAnIrT0y452SZoEPEkqJFpwi99IR
ISMo+93DJfLM7zNAW5HdEimZEWvFG0jwrkzao6klrbDlQJfrCCLFXcSnkg3AhhRI
WczosfdQd8DQZehD4kGuPNX5LnVnjziz8zIqGbD2yrc+m+XttlvPJ3PsJNWAG4r+
zABoODAutXIYZ1c3MYnPXr99xdbSLsS5eYhTZKHL56vLQb98ENoIp3CS771os2Ez
Rlrh0QmUbkPzM9yHhl+HyUeI05G8dSZqQaW1VZSnmORlvgyo8FVnfIJFEqjAedE0
d5cUHnI8F1YBJiGxKG6PtyeqinUX9m7rgPihDDXJH0pVYalMsjFfGDxAbBzBLJCK
Nmiin6qaXHAOKM6Ax75m0PIuajKswVtpJtLsQ/1TpbAvgklM2jfja3M1RBaeager
HAHzQnsCyjy9rUVAzVZ7hfw3kbsn66epCA1EWEMEwponiNTQrUzWet2/kJo+zmqX
FANmgHf7VNG0K7lxS9u0GBTsxAcFq1mHOWrPUUWQ+X8Hj9X4BzhaPGfI+R5LRMcq
8N/HktvxrCsmszag9FswmYHJpyeVrtFwKaKMjjGmUe+B6/Zpz8TQEViNE2o9fa/n
oJty2ZlZlIlZ8VYm5/hOZ9LC7je+Nc/0WbrNGUficFsvM7Uhb6NUPm1jy+N3Ot89
pNLApTUYH+iQxIS2a9zo6LuEynSpfWdNpUXuwP9PUTyfQrpLIFypUHXM9G7VioUV
IeXqTCBDxGur7qXzF63pPe9QTze1TzHzC+VCBl0d0zFUsqWbr1ONay1P3XuWLPsn
wBjpi4pQ/pnirXF51wIKALI5s/ePgdkZvIGy+gY+WfVt25fzcfmmGGYKczvlAhzY
81atO+o8vGs09SNoGqRiM/GRSGRH29o1p/bC/zWkrZ9X7V9pzWrIWNeFJCxfEa+r
2HooMSqxcQaYw26QXz10BkHoWRpPe1+5Gp6/6WwwS2+OiOtdBtd2k4U2o928busr
8Ta7kXDJve+5H8DF2lvX5zRKcnhS+SZQtVuoXnHCaccA1vo8zflHYLS7tp2tLUG2
A93oAlaV9hyjcn4G08BYp0k07UgQFfcNIvrHarplfT6bBQa1CbEOaiUBDF5L9cD8
OGUJ5oYCf1RYF0dCKv/enwdXlquWmuRYE6QPwIDJR4bsoPF1/eZQS8oVMBUBw2G/
DYMDle7uZFp182Le5IqsArMtQI1LPO1zA1fO/YoIjrSeQrCAX8OipN5qBCHWSZjo
uNEUuORzEYNjQjWRnUvLqja8YU/bd+VIs253r3lhaDnKtArx8j4gF9MEmVYBNwCF
JUZGPKkXibKDZcDmJf908U7qGypO+cDkW0+ICGM6SnAtjcuKKpXntk4/KyuRUwQl
pDJopPcOiUCr1oaFrSojgx+gepDdn4yWQLbCqGECfveFHM+MXsRbgUigTJXGrGy4
gtnC06StQKqz7W54snRgSxIekstywQaqwg3hxCTIW1HL21YJZOOIN9fzctPP6B9y
k72+lvNJaoHD1wdmMylopHyGDFjpRQPWDyBTTolwzB3rn1YRNYWrh1fiV3e1XfwV
BGu3mQOGSod/TG5sAXO0A3zHk9qQQYqNsUHKMDz1GWuJsDmazmfsFmdVjD3M6XZh
N/PzohFLre3V/Tu5IcvKFRJYmp4byy4k8VCFe6S4J7X76ZrwfPfhtiE/1u/JVvxl
JewbkuKdS7Lql5g5h2oZV7LJBY5VHMfFia5HkPFmHuC7LXGfBmUlDqal7Z2eJcD2
Zb484Dl2/BXc0XKExUC9/9QQd69/RDCltSvzKM2ae8h8UUWtzcPKpdpzhRSFiFG+
seHbXu9YOFKrA26KUXktCc6nLDsO+AKd5rneqtwFLhBBw23rMwCExQUVz9yrUYh2
DKG7rYlAxGDViR867NOH3OG3VP9cthcThTCOQjzlO896ulD7uAYpkngJfCjQU6ix
JM9FJ2mAMq1yoxKJWbF09SLL4MxISoSVqJ9wl2/KPcsUo4dOC3dkDfrtNwTc0KJX
rjncPdLLGJMrtcPvtHUUkJ0sfW/zHhw/ZQ7tirCXorLEBhydkC8Ir3FQ1M/Y5YAd
UT3iC9ju7mj+9hG6XxAT6+zygLM0pnHUmKZufB8dhUQC1KcSX/d5b3MQzyZl370u
MbtHhcZYfVXvloizN9N9TDBTUtVbPsCEIBIBhKL9kq3QLWXpq+ymAL2ZGB1tA40L
UssSSxXUGc4p98x8/qHLwYtxEA2zD7jG7IfbTzQq3cPGiosec6+kFKCNW4kvl00C
uk2FxdbVJ75+idIeYLJ1Jozpetyd3CwESgS8hyqZ6g7DMv4zVeSfZkTz2EFjhjQw
zh8sPC2/h890Em7k+JvDOag/zS7RieOwKB/WB7tLzYOeAxt01NsIhBDO4wVeEiM9
fOXZ24NtGlVz3L0J/oBQG5LJoz75V2AgWjm4aWTjtPqBx3M6L2IAXQKbg+Z8BXek
cQZmBUR4H8JU06bKMLgHDstAQ01Xjt/32K6LEa0wrxg5t4x47IhxTomMxDe6Teuk
dobeRVgT6c/8GPBdq49lfaPGYwbXY5wWxHsqnOcHUDG+lv/adv0BeYYoxBctPyAr
HWy+LFdQkGiKqdS1VtYs2jmiRoAOMHaqaL1sz0hyVM1YgYPu1PvuvL+IU6ZXt7Xd
S0j+DCFHHas6yHIyMEUaJ08WGwKR79qahKrKTMXx93MnSWMFGNN9vYrvef5hJQ7Q
hAiDVG+1oNQlWOz6ggKEdZ3AMh8m8ylIYSKpcao+vedN8ocnJUQavRmt9lHVpJtg
yVshKJbhh5Z8Y0gAmR+V+xCwXW/4G7/fgEKHvyA/sQQ6H3HSgxfkZRWreONKEi6W
7eR2BOWOipLiWIlEyQH0nE1IAkw974MY/qRhlbsXthQhn3rIjdjK64RCfXAOLGNv
O2IviRc0kdVPqOH7aSyli8VcFwUOp0Df/wmoVz7Gc9LoR7tk52k69IVO8n8bj+a2
qcR3D0uGxsf3i4J8EDrQnpiaMjsbKAJGmAix00oSGJ2jU4dTV8qFTxOoBTqYFY7r
4EqFBEUa8bsg4oGPSxEjXkosaMnOMnOio/zmAnSFgLN5Qk8JQoNfCEP7268QesYv
x61FtyVrHJv9DGuTfaYZx3HezrAGzHSCkAJprNvCS5ZYS0rEcn7RRwu4K4BU5K1v
Fc7ZHynKPrRBPa8Wzu1f7Ujh20Ma8c1IuGgcHb4CNQhx3GprQGKUJGhd6kTfItcL
Vz5JmCE5mTfcYfklGK/rkb279VRAwrT+/Ywb30i178Cl3MkjDdtqQqxwplR1dYOf
cmZumGpxpBaf2MC+q0UVwhZBXhiL/U+44XprEKUGIyK1aqnv9He+s6XibpKvx5L8
NVBq/HHIQIqzie5oltMUKX+BbSOgD5FpkUsaVAXQpQINYLPRCSxtz0O7AuPlCuBf
LM5Wv7sSjavp7SVDN5PsaPgiCULIibEcNR+v5IkqRhpSPh7G/y17DFKxdZozD/Nf
PN95HoV4z2PpPfjuCzdq6JCsMCG6GT/R2CYSAsIhqBZIfUYTuiwERZs/ZIjDFdSF
WgtEbdIyTrHDIliP5DdQ/QNE2KK5S3L6Gdru13Npnvhg1PYovj650pmdmdVktTAw
CCpci0kTK+uLpDiNG3+N5izWCBn6uN+GxTJmcPJSt2mwDqL1SCDnAXTKkiLDNwYT
E6G9FWXuksI+1/3Ho7fNrqodiKMhpjx76+A4axqk/sClfrtEpaa7IpWKvqZyeCic
pC2xt0cPStwPReV0Tc1VoJo3qBdVpAbjMF+1pQKzu92HXs1J2xRZtTIzo4y7v4uw
Hc07jYRamtig8aKJLPyI83wCVWkEQf/erO9DBgx+UpR4OBdZexrmUqAyIvbMpgDa
Vf7MqqwY4GJVq63hAvqCTgmj5tGtvpmsUfFcrJ0++IKjEgJsIwT8NFStT38M/nVl
VJNDczYLIQy69JJM8M6u5APOAKc4FQ0rdG++uGLgrVVn4gWnFRMoyBnB2UZPhjyj
CqO3WSbl0HwEjChv0Kmx5NVaBwFD9Snc9Dr1BuiLM0+/dLvkVHHCfbThRN13jmjw
2pB9YGoaKub70KGKgElL87yJYdW/WKKYAjaLyWgoSQn3s9WuvuR8qkmml6yPI/A6
TqU1qgl8WdmEmT4z9df6MjRKiVENyLTxXS5Y6nc8MmCcaW6Hydtb6EcczbvzV2mZ
mGQmK1PqeudVtBAkpKIk0R87lKP7i2aW1xNufSaJ1pdkGbeaj7o6GyCoG3+g1GCE
4BTbtN3nCgneC+QwLM0d658geWGrhoUgQgXDj9+rahZlWzwTHXJvETnQU9fbnzmr
UMNfGwYeb6dSxkNGqzHPtsG18XfqfIvNNKQIEste1JLKqFs+7qnLUlf0b8nXuV8N
qExeWOnBpY3c/VdTDhGHjDJ8+8zJWfNS7doeuRJuyxJjB48fMmdBC726BiutZLhN
04Yy/PXWS8+RxvFZsGWjQJgPDc3TCyFXAZd82JUu6v3oa6VE7TwbcoBgXbAjwyQ7
IwpvV/GMgoMlgB0slNM3xkDJDoxwmNstmFP03hbkFVn5nhXUy2KgdR0/mZhKAJfB
y+JsPlUEkdX7AAneoyrX/jnef8FIYP8KI66mm37ic4eV9syG62eTR/dTXvpWeuH4
TTXrQyGKaEPWBvno9bf5UOGJjJHf2ZJ4Hm2mEsggSe2z8U+Khoo7DR/24E6DTaN/
rhTNyaveEhmZnGyTkPCjAwKnRu6cpB/ksRCVMVzhpKBWtKd4OwOoYVxay9CfWVxv
wAdSDJjw/C4cX9MtpquyxA/SZc+nVf178bfgfR/t/0VcoyxhbmsXUsf3d0MJg5jf
Gdf6wY+6JCmq2azWiCDNK6JdthsKB+MnkZtNYNOGHBs1vaIXqciV6HybT13uxL41
aTJz6Svkv/I6PeBe1f6skrswVl5y48x4FTUrO/7Wx1eg99iOw0Tux/VlfyTG+JyA
+wqDHHUlZMZ6gONbL1pZMjRrrE/9KMaehEOhipdsatqvJcqpegnN7Z3XNmrf8X+s
X1KtH7SUlwuIQWJufuQkmcCFJzhDURKn7Ev3IFRhuecU6hfIEqdOcGv0DJDnoTF+
w8sJ6jecjk7r9+TqTKrfgJVoce/KSac9nJnQEEPOEti0QwkofprJN/7N7CHf+fwE
wL3/ofcJcBXW3LUMAaQKxlrhJBS3y0tUg4tp7FSrymot5TJ3YG6pEULAOFxJCUie
20BYO8ChB0gSSF/SDQQrnsEn85SGBGOYIXiG0FTpvjqqPhCspSFJdZt6JuUepz4f
lWykMhJjcomD82yg10p8SZohbTDrhIO1e3OOIVgqjHHzLLtE0KKx0ClLcQzXvaIO
8lfmCxmSIiRGVB8DBFYf27XkM7GHAD6kTq+Ucfey0uHiNXyeHFeY8lXNJekienop
/fYk6+oz7QelQP2DtGq+knWinqjeyvjl7iTTiLrWyEI0f58afx7eNUM7+yomkyRW
q+p2eu6Ex6FN0egf9yjVduJwQ38k9pmch9UmBLAaF0LQ0wXBKlJX2ytIeEFbPPL2
qqX2FIgxQaxQY1yHiYCHsiJUlnARZ9AOo6jVgnuVqzERMN7DYI5wRxNM5kAa6KW1
XNPrTVFoueJJwQ7FQdGZOOYHsi1fCw/6eDJBpubSdsk2UY/cim5JJrXKEYALcnWP
z84hNGy8vwBEiyBi8HcVfEOukxUVqEofcYO53ah6flAN9KjoORZJ6NMMIDo5jZEk
8oJkQlUsqBB4GKZGtcMjWsx/ZTOgnO2boGFd/i96v7UZ2MxSxC5J+EO/el6LfKaK
F1lzG7rzzYjhFhCsWdcEMrr4ymaZxv0/OwPElO4qEf0fUlpEd+Vwxh9LlJHJEPUF
f5E8eYSnhABEJPIh4Wv+yCsM3y5o5xkHe6i5kwH08iR7rT5VyYz+WOMWqNAhWgP6
spJ9paN72Jp859Vkwb8Apdcmm8kTX5GfkbW5K55h5HVQyj57OyzILa/lyUEjOJOW
zABZv/piiHwGKnGTuywzI+Pptd2S6IDsvVg80E625Cw++BA4xDRCrUoWMTXAum9G
kEVDA+VUALEGvLRPNbzmmtdlI69U57iYB/Uli58f89WSw6j1VRQZS/gzIQS+WwpO
ufQ/XzXdgb7Tg1ild3Kyk0NmesLP7cbp8W1Pq/dRLdwwvA17DmeQFYgeTbQZ/O/D
0t3ulALQ9IHvNhK8Q7V9UBrR0RKb2ijrROIXqdSHJ3gr1NSE4BzcovOdGhlcOsus
cnXRtX23Actm6c+piUkIDX0Bw8Qb50R3kRh56mnlPH+/Rv48vqgcFLrS+UCDU8Fn
UhyszzqLjeHbjk8j5bcSGzmui4l9/UIEAwiqp+vy939na0QBhkYIbZaq8a5zJh4A
yvTsa7MsakqW9bVMMScIKFRasOLsli5GZFewT1Vu64EKBKZt5NkNqHzb4AhH0vqS
0gDk2T6MrpERqegQ+QmVcyESOoGMiKCBi9W06Q4j3vO/XpMh3ZrO0XjFKkx3RFeM
JQ5SJs3Zi/wyLGtxQ3goIMDa7up8FjVpU0Eq3CqxCsCbjrqHJoDWxMUonAohgwhV
N+qod2HM7m/qvd+XT0JK8Wuco7vExR8CJReXrErwXXlpFkGpE8TU7qqDoRgf9Dd/
a2/wglPBpX6Qhc4kiouszfyEKvAJxyi3W0qLwFxYs2OSSVufhFElpQEyBom2ECfL
MWmDZOZUjHQo51is7dhX3cuYAS4vmOo7N/QCEoJs4KiiKoh+Wg6prGqT3zBOVwD9
Va7GVQyHFs9Aa17H4GUCR0RY7DOgmTOIPFF0ey7Wy4luOoCvmOpjM5lAJxAGbSAX
JLZPFEZN3XmUbLXqOpgX+D1M7n10+8gOP06lbIlBDayFM7Ve14GzQi3VpvTh8yXg
/Mfu98qglTJcdnsJw9qXuzjYjNSsON5/CU/jx1XVeXFkQzATSMIgWZHT0/IM/5V6
Ba28WwuEJxQkhpi48V9DkoyUERyeNPrDGb9KBhUT41611msUioSIDzf8jHka1mLA
fDqZTJ7KG52TIo5V+sk1AXH3ow070eYDunlV2/1yyCmiVuqjRZgC39StoJUcWudr
y1RlKsQkUCLetXAJqlglSz+kj4ekWU5zswAIOtSvgxpPF028bLNfcTeDDNICl7bM
C/NvW/0NDWLO9yYE+fUn0gcV9tryXNTvj0NgKn0pbOEoHCAmd/H/87BSSgkYLHcF
iNREryD9Z65wMsb7BIUclOQ4WjTaNfpzYxhIX+10pTsZVxFVbPnnj0dQeshS1emL
Y/iSuDWE5TOIDrrB6MEAK3PJADvIgs6QhUho0Esce7OiRrOrYE4sPKWxTDEjvEdc
s2L7JJXG+C75dalN4bpubT2mIaNMc57Ixc5Yzjwxgjin24blmrT47Q7qraZA98pC
vKpB/vPhqj0B6/nU/KbT2Bq+/7aQulUNpZbjLr/g2oZ572qF/lx/z/5tQ5clug00
WyiI+DUXb5Ht9aXcmjqYswv7ZxjH6YTkW1O+CVBxkKx/Lvept6kp/bJ8bhFCACPD
Q4JrWFv4biG8pCzkMiZUM6B2J0i7/PbP1VAKi+T4BBOeS2WYijTiEuO8FA7ThlkW
sS9rs4WJpvkvCgZXYYt2TWtx02FmJhRcrQZq6uLkyYlrlybAp9Z/B+fljlpGufqp
zVZkicZvSjvlHczKV/ML8/NYwwukX1Aq9RyGkaJDzhkMBsaFyU9SttpHIXYgpw53
UwpR8M/R+xQhOSMdjkye5hTdCt1Tk7n8PQXw/AXM39bZZlA+mJ42T65PScbSlRE5
4PxBjM4YQ1aI8bDzyvs/WlfynLxCkzDHZlE88odPChwQUACK9ZT3/vor1ATLSU1l
LUtfQTQks1mhzkv6rYtFslU86m8WxYBlFGjFDR8SqtG34B2FvSGBHZavY9V/SR1x
D8idaKNS0c/FlTbJTzRTgMoh/M7BmiuWWmzYjCyI621WD+xXm2t1x57T6dwxwx8c
ztkHvGEH6aUYptDQ8OXDH0cqUv9S8hpZAo6SeeU+XGuw5LfqxdZKPpDfRjU19D/g
GmKIRTJtvFhO2Uymbk5DWcWrLAKc/kmkK2zSjPvtHPwNlwy1ZvkVKyRX+dx5SKQW
oQoTcOSxtOK2Wd3q/PhfyyMGgBJjBdkNiH+c9vVM3UezPHhI95wyWIvcBkQ3FN3O
mTPzackky+loCuSEz3KbD0PgIyMnpwYVlbcx3vAfjQhOhDCLj0a5v4G2zNH9mG7Z
X7CqRyHnMpkV3xGnUfqDOD283NgwoMHY6mjfjRQxmzp9xRnhJdEHTiGaAruenDZ5
hYM190nqElPWRUjHB2pCd3Drqn6+HnZAYrzfxzV8sm76XFH44AAEO6eo3kCT8zOU
DhY1qG2CHR+pNtmQh5n8SU1rUXNNxuk66gmhnB9pUSP94hUh6DPKIA68hmzEbmV3
rajHW5hEZww6ukhM4sXgE0P/5QdNfq6QMtEuJ2+QTWPYR+jX6AzYpNlLnWJHZqgm
+IcG3jsaGbarVQkRBxQH1HkBWDwe6AGXWJ4hc7fw0Y4wPkwkzU5mVSU/tTDLk2HK
MAGcS7c5GfyUhvYNn/A6HVn0BdHx5daXBbdd9YSlxz6y03RHXrJ7C6LQrwKGPyLV
L5Xeo3G6HvwcJAKjKnDx93/cf9zt2J9/YH4sD2nfFrad/KUA6aXvim7XTfacl3T/
Wgv7RlNL4tHmxjfGQxaGIWWG3GMNTYGjr0tBU7dxPj+EXcOZZKhLvDN0a7D4JDhf
/oWcpdoSQTar0M0OoLjmxLa72RiQNzpWFmAA8bSUu62SWDsg9oL0UhvtY4i1x+PN
b5oBLWPnVu7E0/Ac96wIWfWmgWAMd9sRoGmo/kW+3fZyJRVpB3hcwGJlV5+3TSIc
2ADlJBbwxKle/c2hJ/5Sr6qxR0JWBGl5/u6YmfcaxIHb1c+VuXie1703T5xZQ0l8
wetu45nW/F3i+T/1jgef6+GTaRDJgkliGIgK5pp3pD0DZvYwEAeHNZwdiSiMgl9e
26pelctRmFf4XC82wAJgyPLxshgtp3H5pA10tMoY/ByLLCi6aqIqcR8CV4S1Fo5e
WVOsA7SlLllrGErNVoOGcMOE1a5EqhZerCSOzFR/Ia+29GENum95lUr6cT7Lx3R6
8zlz/u8e38PS5oops8qLs/rF88mu3Er2jDV13MYD0V6v/AFerfITkiaxNtf7jWdY
1PuLnLczAw0dhy+SW6PLYERv72QpKeWPaWTweti+4rZqgQqI9AgMria4DkfhnbL7
WpX2uzfSoRmwA80QXsfBxHK/AvVNEXVHtgcGilIThTXcf8982sv5GplRzr6f0lbu
34/5qsXaNBQCJyFCK/YbN7haqkk5DhaUZeMdg+uf92NpIsQua4K2O/3ichliWG/N
oaCyXvBp95M9k8RMQ3VoHJqvSQL+aBtn07wPKV1cDw5r8IL0bt15RLmuadL4Wk04
kgW0kIc4vDZfOQOJjsK1iqOVseMbsKtcjdqE1AmjVLvY8aYRifJyhHYy/8+JRWs9
3zQOYVxJSfpO69lioM4hYpPOeffEhtUI4YcfnR0USSPcfToPcpQo4Zt447/dZ+6J
z1piGd/JT2EnuxYNxglYtunprVhoGTqp5xiw/1y5DnXBfBYZJDgyN+brAOjhJVJ7
UQQ/jNLyCXbFRG5kX/eImwPguKt28mfTyN3Wt8OeCNYXDRiHsnpUog/++XzjO+3s
8VrN7HJubSUYSpNzm4JYyQSsjIHq4wsMcy5gwLEMnHbRQjjxLNgQc8VfCDqHwoIV
xGzjWnNw8dYOfvQbJ10MmL8yUvOuuPwMQPX1qOOS2svFlCUgctRU4sDrOYtkueZf
g7Ig34tO689B4/AFymTu6GfqqCYUZguBPUexXwd+adWrDo56uhko3ARKglHDhVtI
68wesLdce6Br9YAufP9EUMZijlJ3CSoQZKIAw7LHevvs+nnU0OWU5QduXPPTICTU
KMqnlgafy7Qw5g4KKz6dQTdeTHNT4su8d7KSO+klQP5UzKcRDeaFjg6LfJC3sygZ
H32kH4mgmcIf2lvK+uQFvWg6XFEvkHaIexTqeuxF0Tgnc7RNWL/MObXi3sVhDZIx
aXetTgM/WQ0ViN6OOiyaoIb+KIb2acivWQZ6Cb9HrhfHxQpEn0zLwVn73xe1P/DE
AZyvbLGJTSbtpLobgQCQvYW5B8eb2e+CQc6MIOg6m7ZihCUA6akI2sQQ24qIpReY
YY+N+CY7it2PckEaICKxcr8C9mrMTtVghQJy4t/QNOW3VqzOduaKVEmIOosSeVKm
ZwO/W8ex4eBoC5W7DJNedzfjkg4P+fJBeSSym+Y9g/nRIov7DZlpt/57hKQEiXIP
uz6zcO7Ju8LtSsLyTaRbk6D2Q8ck40B/djBA2O0rwoJIMarKvmWMCVtDTTjuSVBM
llVO4/4FQkaN8R9JUupqUMdZt9fNfhOuuUGxNKxcib1N19UH1/x3n/ZjYVyTVIg1
n5PUqs/wYdRvbB+fks0OgYZux/6WN7hz3hGvWN7HLz1rlqZRfoJ9JG6GlBg8hkjS
m2NC2XblJ+rMeQuCXeMbR6xrQxNRsRwcjqnZQ5MlQDBT4POZmXQUHhdBzUer/rGm
KUOiBCY+PBXjtgA5vpkGjyVSYEObVqqBMV9E0jgXo3hFLcZI8n6Ap87pfhgi9uY0
YfRqDaW0tgsET9P1/is6kxR/uXtrcWg144koyYc+3brEUDV6y0RYpEw6UYn+RuAg
dKDvkiGACGoTQe9K+9lt2TuBucCD9JGgkHaVDKRja1RxrjI/WkKE1s1DE9vLcuAG
Bpinh6W4BOmyKVEYq1HE4UMBshHDSn6hQUNyJi0hAeoHtJRDN9Im5Atym0PkvMsx
PWiQ0UkT3MJvvu011jm8NZZ5YqJFcKobGH/gBVV6ZXKlSxwgsXXmMaBPyQxK18lz
tQ7IJBEvxmnFU++G6Y1e340sz8+jzTqch4n9CXsSONVcR1lIbItMyV7DawW2cllB
TJy6w/OEwwCWSlmDiGHGqAubDNTCYZR+J32B2LSv49gLDsSaDTEaoUG1IUJZALR4
y3x1ENztmN+zye35sr2GGa1rkIjsoJbY6eteiBV78moHIH6/meRm3hEk7YhxSj4w
2HbSy1icpslXEID6gPE+JDLiE3QJtQkU+jk7+Pau1gFHOKJV2XVNkgZb5Ls2L9p5
rRijHxd/Va3H6H1RKdCfidXg6sSVXmSYLpQ6uwxycIFkBzokfejO+zSPT7myQ8jK
88PXQFKGBowg7yo5ta/iq7+WKrLjSHoBcNLtXPAu6bmQ5uDqK9p/+TdddfapvDtI
CQVLiRtTbaKwr+52/9/OArLZfJzmY4p5Ijch6PaGXXGZJIcXr5sCYVoP7WRtQkz0
4TxD3ngZHDcMSFkyso1CUm8+LE7sbUEOwgV5ZDsSS7sN92X5kKj26B/ZjPylu4QY
rkDZaR4w6A1hqIu6BSyXkEMtXRTSBeRLqNa538abny0ZgIMGOPhXESaibSB/G2dD
qI9jB1L9IGtlm+7TFKm93nR9Hfw40IjPxx11gNe6f1wxLE+yHcbkgW8ETMMnIXbx
r7NkJLUQO2X6Zd373sfiTwh98PE1VUye1s1aHdUXhiZPSKj4KfUEVkLPfmqdF+6h
cfoAhCr/hgweD4VAvbaeHRkXT3AtnEgUhxlE/QiSEwaZCkBGnPITbMQpDRHHhZmZ
C8qFk3ieVbX7uRaE5EUo8Nb7DfQj86RtGhR+b3KLpeu0Bbl71y/FIk/sVVZWvQyd
J1TXYziAt++C2rXZDb+TpQPZnz6SZBFPn7FtGuUi/Zo70t/ty3uayI5zlRKprUgQ
TvUic6JstBq4LjfIo5t5T3gd9bOZXjuusA0XGJciLwTYIgNSkDXxTJP//c/iaWr/
jNrV5k/GHdz4KFJSx8sD9B52ARkCdpshAGj6lyL5Yi0xC/jdGzzM1G/I152p/vME
vdL1TivfHEca3QnIRdfs0iCa3mf8r/Mv+v4/l04mEuaNSYv/wDjN38bASa+SqbU6
XQyfUMLPREa1KNCvn7dKmrFKYY0Hzr/LG3CaW9LRZA+XomWWRNmddAMo+BePQrtI
y52LogdUCdgn7knGI1gy1xgVeFUvR4MAR+eE6Q2jJDfUhSqq81vSmS92cuciO3HR
8LtXVleEuoiIfEbBMxzt+9Ose3Kzc9FJc0D7jVZPMiIBS8wAFZKxvD/Q/3rHbiyw
YbEVcIXo/Tgxz1ksfIWHFq3ABNIqvUyudTYBHdggMfCpAKGtw9ztqvcOqw/rvGEF
iWAr6k+kIhMfOd0kugvDvzTrfIDFDstu/VfMVhZ1lN6B3ckuNWavhmLcmEc7p1XB
Q/QfIlGxacR+fDJwP4J19paZp4CO2AEzoh9CTtZ2KPvzPJeLMSZNgMv7QXuiNEgR
kdiir+Msxp8hD8ceDhaT7zMLLlF3xWrCudYdgQr3x8mOVzddGqxulyHdTJSRawJ9
ZF6k8jUZfL+iwsXoD1n+xVy1pcZt9+RdnG+qOC7TsBhjkGyzEOJ6HjkvS1mTC/qn
kuw5+5YwhF6bnmOChKwIzQHzi1c4ORqhSm+60LR4Q31hYKDk4bhgUPi0qBUCmLZB
e5Odrh+53+P5fO5f8s5iwxj4D9gKHTTNfKcbRaBTHpmYTYziQLtmzfezG9WBbhtd
5hOyoBDD3RLT7+TW6zoOgD+4B/zUV3gwRg7NEogdVaAr1BkB3vvenP55pYGFLyM6
CQIaoxF4Jzf2321DsvMtxWGjcxu7N6gR7x9/IFgT2qvzDnB4L7/lmHbPjnCmj2WC
d4Kke4O6gdFQ/tEp+1I9d2tRoGjMFASTtwJqcW5s8mqH90LkOkd+Tw4nW4ndyk6F
r6MiWVXn0JjghXZOV2XBwKRrxBBn3gXLeCP6apTknd5Se7WIc1NMSqbXP04EkCM6
bIpcv8W44a/P/PejNiByMk8IeZmQVLlYEomNqUgedJVTb+wiHQsmnX37d+gV5ufb
A4TMl4E9jXY3Ytrk0tdq7B4A1cKCEjwy+MveBVVJCKHPv2NuXk9FFgbSlDJJgES4
OMLQPmXUoNd6iRLR4QoBJ88OZBzdam5HoJdPAY0jvaZIG8XvnPFEzlC1RLLfJCQT
0z+S8EwymRZPXUKPpi3YfwvaEDi+AXr8RLThQIlN3GDk0a9Eg0wjRgDJV4+Kazfd
HqyCLq7cDH0tR+MOnPenAIIU29rUb/HDR4QtiwxJqOXZV3I4o6SVUQ2ms5qrn6Kw
uz3AhRG/kiCIDmrfmj953eTBRUylYVT2QNXGeabN0cbCrVGmT3djMy601s6iza6/
k9UTxFqOOcFlhR38IvYy+7Lj9vokTo2eRdlo5Qay9FjGGe0S7mMEe7iwod07vgQo
7jKDr9jV9srRORhZHDo4U1cPN71uZby7E2DIIy33rtz/BslmZMD5m+rauWYDVayG
X6fYbVn8JAVNy8ZnJHkL9jPzIafkqgf4t4mhDzpZvlxFfXVrBv031H8LHAac7rOe
tZBexZLIXTWUDOizhqshpVeJenOyFlZ3iyelc6cRtokeu6CQtgvth12ne01zUSFQ
tP64mWb9EKCuIPESV+ApiOL2u9gy/EyesuXCsqkvdfAbvTkZa+Qr+IGzHLWIuN9N
DR7rpTisNzRxMGpfZizLtLAO641vD2DPJPHoaKTjf5yxYblZCfDCICKIZram7++X
DcF1W9Lkesj8GEddSfEodUYGWNq+/B6yd2nRVRDIdGxcpdBh1FEZQqrlh6L40IqB
7si8OQdjehkoIc03Rvi7dXW4ql0p34u3k/pXTgffji9OhbzVgc7pXEU2bhzIWRC4
Aj8D94rNdMgQNSPxzUYgWs/sM3rSFywklIzawhf0pLtzA8IAHfkTUd67M6ENfcnu
ul0CaWKJY8ZZ7d3TUklge5OpVb9LJiUR1v9LgfgW4iwyddGomdJfu7DNxQ87zJ+s
8wao/CsQvNymaNktvO2KCtfz34WvFwSTV6fdrx1GgeykK5OBmrm273Ie5Ixz3MX3
5u1/3bSwp/PnSG1oJy0Iqol2hy4WwM4s4h301Q4qISSYd5VKhVFdxNqqIkOMaKoh
vbSmethRghtMyDp30iTe5C6XG4uiPUxaVTorEWeib6ZE4HlxtKdb1d7h6LNv4f3A
B0sbVbtW1/s36Koh0sfuVTlmwv4oZX3ymYN1aIWCZ9lsR9WO2waZ0b6K6Iu6BN/B
txQq/BqAbHBjL8WIAmPduWZc3H3WG/yXi1co63wA8REtl/swmruR3s5/YBf48jcu
3wFTy8s454pjWGlDP1qAm2tTdMEWxfqM1JZiLtIZNU2n+9GQN+empW/8kLrlVf+j
tiqS7auYevSq/m8K/b6yOkBBJh8b7RBXz+Ta2V5U9ACtkeyKfIQSK2QLFRrU5b6+
nLPpwkAkTquj7rtixXmQgHk3wc9CQm7jyQ0Ku6GZIwLswvMy3w+SFLTPmtrFLqRe
AgmL+LPe3hewmznNaFOOPv8pu4d9ufcLBUafXp2ebgAQdiwk0/sfJTcACQrq620N
MKcVQ1c7xni1qDNrkL4zb7glCnDGCLRotBDYg/jKCzwgzj5NjGfXxCwkdxSFFJVj
FezBwO+CBmzqkCszavF4XrrbdPzpo8EAL5uGgMBY0OtKq9ZVrgjFLRzOWnG0lKLN
Mq6ESF9TWxdsFJMuievoM2XAgt+DLgrRIXqcQnEvrinw1Vol+WBNK5yg45KqJpzV
qqb7sl6dYDef5FU0bfsL10a0jKeqr9SVxwnEA+KAXfsZ9A9LhSKZvKcz8HOFbCfr
061WOealWR266uMsZi00zRXqhDwpj67rWCeENc1WK23P4/K4Xf6O0DhkI4NWyG37
L+byg6AetiuOtPpaFgm3QjW9BYbFa4clo4/QG6krZYlqCcVaR0g2nvEoh9pNEJku
yIx8XoO/Cg5a51QbFE4rqGsrV2xvfVHGl5hT26qIBNQMeuiZ6+GGxKdb/ZKhmART
zdj/d33iMj91vv1FGlMm4+XbQp7FeDDYEQUXcfA1qjT0UIb5Swm/NMe71ST6liC+
RegFgAvb4n1vhuC9N/VHG6p5y9L1/6YMOp9ajUArjnPZpQtnmmIqVpQES/nPz5KB
kpJXyGVkw+gZa0WCFBB3A+q/0b6ada/84PPBuQyZCGv5pmBWPRIk26Cl7qOEjibc
gjjBcvzLinnTpK75bqlDTCvv144Y0ISj7XrJ+D5gXhExWDSqgT5rc/6DQSYfGJjA
D9gmK7Fb8IR9r/KJmR1IMGYbpG66xjHgg1sVhSX81mlkj2ObW+ZIImdEvFx0hMyD
LPIFgrMAhQ4fXgpHrw62GnIocOxgq+AZ7pTaRM0u9DdSoG1tMJmGREv7XwYXIIpF
X0FQJcLBBH80d7KaA90XK3XH68tdu6IgXX8QZUBDxqATW5hWureivTIYgrYjKgfK
9V0QvF9RtFBmZmNyHc6EuQ+S+wH7xfrFLNbkUQSoYOlvsE5W3/nhNx2YFKanpdXc
VhyN7wLt48n9U/YBTrLO8BOX06OBv6OlCtkgZAToeh7GPko6kxH+WI6D/QPwZwpw
csJXj1MpwnFPBxxu8sc1VvLYpoNLVHPfOOSy3FLr4A7nEZL3jF/5j67vyHINUFMB
qI/Lsbmmay0s0jUMT8ij2luFFsS3bw6L0JBKHEgYRl7Yibe3Ha0ghkIr1xFHQbfJ
IfFc0FeYz3g+/uD4SoXu4yQvc+mRqez7IyWGYDkM0ulyQoGFU2xb5H94dOpJcu03
TfGwRN104gr+bXWDw+C2VnmZrYKvaCo8OzmJNBuojqTBPtYZBPefQPUbPhIwQlpb
gCKGBCi0kc/EjU1Q3XUodrVE9XT2/FFZ7BWZMv1Azb+x+1Xt8xOp07S59vJzfYHn
/2zcNTsftdPLKjmUSiOkN/Xk5ESVXK7OLx6nDYnAjP9WilMmScZEOyOE7v6dFYwj
8RS7ebrpr/MxsTxbUQ1ISSLs6lVjjjcbZ5sRTcQUxU0DWbmEOSBD1z/w9A+C9TkT
dsBKYzFJugo82v4inupDATIx5OAlLIo7g2yw3k0XGnguMEB+/kPQSCk7NEmccbAu
JzZfFWzZ4IPpzpSMs5KnOS4TN/ddUX/+zdjzOA4LE5Zx/e/fPgfRdk4LH0X5X3Kw
G5/iZsaCeC58tZQWguI72C72aKI/QszR5Io12zIN6BF4wy3rCq8bkHGRxQ960uJV
EdhgKTEdobfn10qY/l9e7oWYkORQDpnLdDnQc+w6EwPOi/oTiQbc3X8b8yRoTjIe
CHRMWPodX66N8OHJafdiwi+L7NOnw4WQgN3HR+FJzVb7LzE9QKMN0pGhljST8f1J
f6HaaURmKv6oTG2n1IZ8Yab/TCkUT4me/4ECg532iZM3cSVQD+oKFZZrWt52rOsD
nb/JyW0YVhTQFfuvTDF8TYoeGcSeMYYfTLG4HkcxWouY3OGDXdg1pfZp6GDrdo7b
2Js3DZxN38a9+QGGboklDOfd2Jb4PeyoyUP1NctbLt1kVL7AfAP3bp9ARZMyWHdE
BB/pAwWGgqty15WlF3ZFV2RSjg04RVzBSZTw045dxjoW0GQoEvCCtk3mQM+tUBWo
uyEbi/eYuxX0muDq36WCVrGUkmQPjZU60ggXm/+yuiv2jeNj2+Xj+UAeRmbKds+K
30ojts7KhpsZyc8RtySfJxQScN1aNNNIynCWE2RrcPcUh533Y1Uf2JkbgpvBMrHZ
mq5kwqDTYi6Pj2f2EeqSOp73CyTbE/s//ge7EIeUGDTU3obKmfMFb73CG4MwZphz
Oe0Iba8rrvlt/hWpx1W/3ij3xTLbaSl7osxb2BuO5p9SKeSHg7JwzSLHbMWVwkzV
17WaPWu2N4CV4987oNPn+tw/JzWcBmhS6LqTQIJyJBbcbxZZ1xB0LMoz2EUxN3by
xRWgYCX+okRyHc3pYic/UvPuHfEZrWExllePo95JwNeh/GQs6sObtnHWdLA5KanZ
uORf39TdViFqjm2p0jlgjnFJcxkbq3bIQur6nM4o5w+6VzVTKdr1aLwr2puBJ7iN
2C1G5m2tcOo776kt+Qkf8EMvczw1lp9+qduwqtKXE/jDpM6eE5IYJYUvN5Ee2MT1
vBv/h3+hWJD1HEWi7XlCKhBAi61kxcT6WPzEEyI1PYG1/Ss6UwfIUAvXaTpaxzUG
BNheB06fjne4aBmbrCDH6yy3as0PfMQQuC72nNEJc4iGh2DAEHkf2Tauzs0ZZKOo
dYMVXa7Z2beaQPX6Qla9Z3+yTUPlQq2EwqGIA3g5gfaUUwUPB+1uQ4XpBKdRgdGD
vS3wfwn8sLqdFz/lwIrRLiozmlilYqzXoKXX9lHHLHXIIea0Zb8XoAQqiGlx0RRg
tyhffhAq/nM8MWwwfb5lpfrq+kDQccTxGbgXmT6LbXChyvfpagp/ff4v7cckXYgI
OL83MrD3RRkXpV4Kck+GHQSmgjxH3k40+mqoVoUYyYCCJUrQ+S/wF5RVbvtTroxe
Sd9hjLBgKSfwMRIKgNhxy9CION0TRRJYlvjVzIXHWMM7VeSErCDRi+z7Q3+CE8m9
ivXwSMqqxuTo3qdUrgobVFSl0tOsUMMwKvsYUmZELMB2OVz+wj4T+/eGGGhoFdSK
OjDn6Dgx5n4UlT5QqOsNPA56wzyVqEzYG/jkFmi4icKxOQMLzFzXIGxEPJmQu3uy
Bl9v/1jciZ1m/9aeLdmwRWbsqsrcAbrPpbal+PN8XWubVCbCJZ4bVZKOaivBu1Qx
OYMmdpokOLUHUkGpCuxgKM4vDeBO7+G3X46iIOWnzOv3ecLtznrQslaeAmLLqjYs
M91YstQ1n7EqCeGfKKrfJIDptX1s4QpI2EnnOz/EBTDaOrhatfBE2n2oeAs8skiG
Jqd8DdrPeFIlaK37GaRHgZyytNkuxyvGqcffQRE57dGfwVfre+ip+FBe23nYo3II
Zup2q/Ttt/ogICBe8HBrKb2RWTZyQfP0OnesAvej1xq3zi6OKvMgAgJEFk42t3oc
Ylk0S+e0Gv7hQd2HRU//WA5pYqIVlMP9CQHm1cy/P9GN7QeXMeGNg6KcgwVUzjNY
ZK6487WYKjeNCtaUJZq/jxQBW0wYuFiZNBvQh8+WM5EWGS0gcCZnjNA53NZoihpo
UnNevfBn9POm0iHIO9+JdWgiTpDLeK3HK9xuWg2TSbh24tStOn83/VDAa4d51j3+
dM+3ppBquTa54jwXbuWi46/2nI0di9I6P9W7Spg+rWCn2Z/+WiKBlDqR0jWyWmwa
bne6fX9U1Z0P1yLOU44nlbuAQX39T+/pN3rXX5urPT15Wm5RFW2fF4ZrmUdOFE7O
aEv3yTd/7LkEhEu+OkWLyKSXyzPJ1mmsRhl9pASWAsQJqyNJz3I2iVa0DZFaGOQ2
4fd1k0L04n1UXLVvuViU5BnpxyNxYVnfzVSa5xi+ySxkytXhrk+zkzIZO7Zob7zG
s9l55yuoMEgTR4UOsIKpwBRkDXpGUFRiJsEwOHB+DidT0T9QtmY3tNuRim2xyT/d
1mNvuOnnfcDGrM60NyZPcWiLJHG8mP9Z3j9ylA9xgrhRIYfdr8SY9yXH80W7+/Ns
wk+QhdBtuMg3tRzHdPlgO/KDQtGprc+3NrJZvUlUk/8TQMwxVBVmVadTIDPhelPN
4bSWTf0rgImShRb4zxMzHpLCJcJ7YN3oJ2F2IwLN5j2bSVSbVyK/vo432C3+93SC
qWynTGBrbMUa5is+0+eaCZf55Pb9AIEs1pQ1HaYw3b4Mns7TJF1xtvYDx5T93lxL
tctVSz0nw1nMynIqhYK6rxMKG79qB8mr6knn9Ti29/6tJB2woo2aGzILgVQhgs06
ipPoOf+q7EPbkCT1hjdyH7+jzFgbeeWP273GyLt6KA02n3cGHicLbOnNaEbttIQt
OBFRXoF6dWEQAFF25WMO1dG17AxoIGbyzaLKtA0JfoPtVtcL8CVgcJ30JO6JAX6j
yAEvVZIRMsDfi8V3Bal1Mb88y6OrXfTWHQujxHe7hT6vs4YGEsegUNfXsguf5cnw
uv3swi0Y8H6jn9jgzguixJnSaPdDj40GuBo9VjEQ6nWN+19cARXNydn2mXEcYLl0
s3FDspPiT91GeI7zckUkyJcls3zqbDQtazREsw6mUPW+IemOhSD9wfE0XFRLhquU
XIotf3Uq+JLCXGd+cZpFlPk9I0uZ+Q7w6nIiQG77RE+u6NtCpmhiCavw3rvYSTG/
Vv0X2cxkaCtQ1p9QmzsLtYlFDsufRCmNgUNmBqC+SgpobN//0eVAqqkn2+2954cE
3vJHanzLqnNvkOSXg99tBzuJQF4NBBvRmJzEddy0TGeAH88hBBKk2rgpOCouV0dq
KPQHCvajXeB3DqcO2jE2JjXuIO8Ov8S52fhmz570+J0qb+8o0zlPt8XdYVid4WmO
QWdG50d8qj971Uoc0CAIYPyUUs0VGK72vfssQvchg6gm6gnYyJYaYumjKfTNr6iW
+uOrYASDU/vn6kBtJN1JWoO4zv9A/xyAZD+vQRxYIPvkpMb9vabbfeAowzUvp5hk
SU9WnKLDM+PtxwzTrV5LQaHP2pze5gn7yx8z6mUqqAJE8LQKiYVKfsGVjNZdoBXL
NmbODu5h9Y06DS1nn94D/ojIniWecT01EqSkY38atiDeclDxHyezu5c1UOhs6WFf
T8rvuRlYB4ksdSKiBWc1epjvjk2PlDBt1Kew0bkhKHD/6r+g+/QMOqwo1hNozNKy
9jzQCG6BG+BhwDbguFcLnIthALKfmeojszd+zwCu0cBXSwYbzNPzSBP2ihPZiv1U
thAqumGxhyxAZZLJ8QbxokbnZ1ZBToCXzMGsWTTQSbPZJuUkcYdOivzseGjfflHe
ZnvVcQ7j/E2nci9uxN3tFHkzR6XFg0TxaTo3g61QYK2v/lM4Iew/SmHMdwhREwWL
TrvSzdljud/0bemYrDFdHKUm0G3CwvZY5Zh1zmI7MLacFPCBj4m9iX3vuwsyNbxX
5TFFuP6LD/wrvSsXZfabgrh55vYXygW6Yk2xUcZwCRnB+uf3cqL1XJX5Z86RPbrw
mz6fH4fbK3MiwnvjEELX+CDLGsxNJMiZ8KIhUGr8dgHziNQZPYiRNRjo1J/3ei9F
JY4VUYrTD67sD8ud5q3pfylEUla04oGZOH3YcyTuqMZW1LudVq2MZyfos8THEC0Z
h+zqWF/AVI3zZofhhpdzVrlnaRBXdwQ4HCjyEaLx6yKBbe22T1pkIMBDII/UjmlB
bCBZ2hmE3+GZ29hXB7U9qsIA46zPFHjaWOQspVvHjIgKDk9L9Htyicds8gbWgIX/
hdG/c//uy9se+qGGUgnIkWV3tOgXzGM11pRG17MONzcsH+3c68lgV0qEkX/NAmgr
3sM1PGwro3kprgYp72+WfnlbksI65SgyDePbZIxk6hN94jzaux1QurNx1W2Kpedb
oVS3IVZYdZ2s+kU7x9984aac9lYIHZaHnguZFFbaiu4y8kZLlcVj7BXPGg8XtDpu
8Ccm5OL3UnzuK3KnLdslXQOFHaqNZKm7pNE72ZvEzUzG96JWiUzeg84V63SoAdOG
vIX48WULjxjgBB2pfzSMK2EznIw1wZCBTmqZUM5bzAIodMMa+eNYYsfK370ReF1n
crJvwVvcWuZhTjizDk5KNKF9wwcPhImLzdMKFgsXTBdZGVqi9rR89lWLGolwdK39
RcRBlP65E8WMX5fDDs0Ahw/zC2mV2I286tJ83K6YcbA6PSXCRb06kbUFH95RAawv
gYo+xkL9em16ovSLEWzDyIukZzqyBFI+8TCGL2n+yYTXOa2+IUqigKqhiRkfXk1T
/afZEdMc6tBaFnDKo4HTif+TK1M+0xz4VappfRPyluPACZ+oQLeJOn8mg4XOqnMY
91Z6uyM0djrtUvwpOVeEMarxIWdXxyfs9va89PRyOGqwqVr74fUbNeNyUuzpxH1K
auHKgzEmR+vOKMWc9K9RTi9ZhEifch95ol7EP32bIaFtqj6nCE1DkwJpVzyXiCHk
8K3sLWyrpJu+g70bLBMBjypPCKCUstKoZeasJOXswcCv4Xanr5Dph046lD+Z5Tj1
YCgLWfbXxSYqp0oIX45/35z9tqRI/RlCM8KAZXSvPrO6suAfcPM7F603d+ZuPHIw
fHGxDcRGuEkNVMDSUh/BcmpbPotrK6fzpC9ZgPOFDW6rd/MbULM1lqY01Dx0BoE3
70aIDLgtDLnmzPErxMkuHsiFOh+gg++LWaaBzBb+v3OrR232j5wc/IynFDHFEl6l
3JDP+FDs0mtXoGiqBvQZt+U0I4FZMB8tXSM8eGq9XNJOxEhqR9VeyfXoalp9rRPb
EUI7bv4Ul4gk0CVjKsq3cuzcUdenHjzOMpYpDQCOK3IS8oku8on2xuHnF/pWbckF
MZAIc0Iq6tbMdJHExXmBdYrjZ6PuHcVkH2owrS5pJUBamtr4J3tgPifp5qN4heyG
n1whKchtFj58z6cwJNOJXUVXfslvxGJ7g656Hydiu/Q5q3Emhfs431A+OMNY8kG1
G04pL/Dp369atTb4EOX8lyXWBUS4Ezn1b2tqW498YJG/xpexDPCr3Dt7TqZgSATH
VdC/HdK4sSkmmQ4tQUgNUlPSHBdop4HBd428HNEUhSW16m4QddRRw7es9dV5lXI9
pX6ud4QW1+AGHtoQgqp4BwG6Q3n0wyR3tdyOzxrFlqr/GB3OhjOjGgmYh9hqq3nJ
AOrARn+LopjGXk+PtszMgRFd81E0EfYxwVSdAsqELUkIWelJ3/tYBKDhe8lMLdPT
g75XNTE4IeL0xAQp3zrOKxwIT6S7o5u5LZgF4b+pFoPoW7OkzruBFBEukm4QnVuY
qUX5gC0mmS+IrOo3xEsEB8SboJ9d/3bFmm23jHqagrTPeaIQJ8/m8L7nOqe7W9sr
mF7A1Nns3BhUcOUPoOusUos9sOTlF8wHdwOLBl9Wt6RuZclM7AHE/UejmCByF6T1
/I+ZV1bi+hR/qr7VTJgyTHwA4otMQjWJmI3WolwDJwVFxhcNaj+XjkHuatIpdciB
YQmN4wkBHIxpyCfUeWvefjnlTtsH8bYrDh0Ahu47N9d0gCqf+MvuLhGIOycze2Xn
cEZEfKyJPkx8askobTAseNiEW6hBxJdaePvS3iBktgUs30jrkGrdDP1OX7vTQMG1
/88LjhTZ9zWNrNbFNJowI2IGar3Du1I25dB40oHaRcvzzX3V05OMXgch+StxSVm2
U2N9z82dQQBz/lSHZBZ2SEpPDyHe6LZHjM3Pv8sGpugjl89z/tqHgzGf9pISJvPv
/Hqyb+gi/8BxIEtcnhh1RvdK46yaC/zJXmVxf+w8BfU9dbJpSEUyTW4Wi6b3gneb
al7kvABSXkRZYjHnMghywS9HGZtTtMQkLVJR2SDnJQTtufxBIIL4ash6NUSilLHx
+LTuC8mFiJ7PgNDmh9Iz0kxnhDpK5LnoiC3F+bvLP5/d2Ng2utaOqHjyI0dz3d2k
n4uWxz39pF6dZCczUK2COStTw28MDzCghxzVBivrRjgRrSOMiLM/CbfaSSpGG5Ko
WhbPbSRXBeb/Q4bU8kIvikWUjVIjDsS4E0pRsQYctRPN0oFiHDjR7kbqqz4mMtSy
ibCvga38kRundFWTkYPg+ze1ZsRyuvlCPPwgErxAtgYHVXivYBrJ+ht3nnYywtn2
pvbptXw/YeMHZr4lYrblsjplAceCEBuU69iugcq2xdriY0BYoH3lbkbdOZpLfqIS
MxaHBINE8yoe3a08l+dfwEOS4MtD756OqOHj2uOJXO/1cVo+aa36wXsDIvpg+B4+
dL+1zTnwYIxdHJpNCnLeOKwXK971UJRRtY8jgmV2ZigqMp5vnDW3SHjs9JNTRXY5
6mRaRP6eTyMFWc4rHQuRWUNA/uvB8YPnFYPuDiVbmHqcD3DWuMmvAZPCPon0fxM4
JLAhKT8SpZX38UieGDlHuFGU0VJEYNOFg7g/l/3yKA5YTvOJevrIPDQTAcZ3BmK2
8SVrCjDYqtw5sK5lDR/B3ZYLOpUXpqBPv/zt2j9NKzm5V0l1cvTiWiXl9j8/vJg9
chJh7hGK6nDtEJKGFvjVNsqoG8ePANMdOJnF3nBbHICzkGaAjiMVNflgztyY+dqC
Gtv+WJ6i3mVscuix+ZrxrXpGAxaWHr83dNxLOSsCI7rNiAf4AQQ+ZUd2A4X0e8lK
QbYQ7sxlfAdb3/qvy5DJKh8xRJAefFpuj3ivZ7YV153f8b3/BMg2IpkiZh6T/vGq
+DrxyEx01bEU9vK//fnu58u/2UwejaoNtCkxxoKnrhD63f3Nxa9z48fWpEGfxOsA
uV5647Vgj8WF1Zmzber8CWjuDz+Uwn7FYL25yFojkcwzMMbDRsA7kgEfSsGAn1Yh
hbwqk+eT0//HSCWIBx1uxICmShbPE2USuRWahdoP/E9W2X5kkizolAiXmpNf0C2x
1ZEjOKXS8nwhmkPEI58hzs+yn7InCJZt4MhNKLZyV1w8uS6V+V45LRDceh6IoF+w
tcViK3hFV+dUdXJh+rWGudh3eUfZhjRq5sJWtecr3SLy6Dv++8YqT4WiNd57K5Yj
8kRTkDBSGS8y49O6UcPv35DUnBW/Tb3m7avI3VS61DlUZXariX9HIl2VA8Xne0Kp
4rYqHZiB57NwIqqgwTcdzdunI7bO87pL17/K3et++MNG80ggbvKLMZQ9UTDT9IdJ
hD4VuszqN1v75UAQ8G3q3q8jB8nKqDq1PDK8u8NmzH6sZF9MXIg0q7zlYmzgWHxY
qsaRGTQLhgErpz5XcUob0fO4KtDC7vfcmpG3DMKp1yWf457IoHp7k6Ku94fm4SYq
Dt2wChzkEV2yPbxMR5AI6wS/UxGL5EZZjdI+XweeVssJifZli0g30Jy+4ViojeGB
K9Lb6sqZOWj+gOHFS1I3A1iLfIciX3Kf5s9vWU7CxyCvEjca7Hzr0K3p27Lly2D7
pOSqoDQDfTJFktERJnKy63H+YVzvqP4a2NzpLzPRPmFJl9cg4SFjtDK9aDxDGLbf
rgeGyy3DUP8OCy8u/Glc5Sr+3oZy+UtxR2lAfbPxYbXEpxCxKlo2RouHtAWn/Iej
OQCmSSyNHD1RmkoU7FW5aCVDqaAhFqH3uHs7qgqVzwKjpahoy4cLgnAd+NwvpBa1
X6X36qpu8l3xn2y/4XCCgWqU/SnfidyhI6o33e+yiyM/0YMGeAXqwcH4Snuhp4ko
3ZfEY0iVWL3HXneqq6xamOINV8e+qSxav8+hMUyyjzYveTRuOTjeS4vFN/BSvyRB
zABxHgc/oMTEhU9Qya9m4wJ40xwMahpRTmwyzOsY8wEFUDePZIELsQvzMsjE5j3f
HJ4BHudG2Ea1co+RL64sCZJQEq9oL9v/xcE/bPb0Q0HBTC+hdRWWSJPUcyFNCSkh
5A9celijKgJQVBTo4XUE+Sj3/XBr0cnOYIqaz7Q2mUgvS9HXyAFikbe3ke/bTj0P
1rkIBoul8PyYYLsE2bi1tam6SqQr8kPnE0KXuqWumXKtmhOkNu13uhkSVYik4V6X
pYtLmbpMcAAlZBJ9pUnW8o1QlRlBhkRJe0pz347zy75eEnX9x9M51mdaMviocE+4
m+uauZVarxS6rAOr/tHypvo0HRSWwjxqIp3A8NmewVTAQEugRk5p9/aVMD7348xd
c/g4/KoN0J1AHKY+96aWTjOdmvGX/U8B4ByxvEwoTaGpC17zC3yPCcwx47HLad68
ri3UoqsvTvcA++0UEYK/g2D5hRX0RHVAoxT1uSrtHcfl989sJT3GT9nxdaYh4IR0
P51fWkg6KbKGOcB6RR9MqfakSxTXKW9sDFBKzSuR8Ga9xpxIEpihFDkCC19XQ9G1
KnZauGxSBjUWh+4+XpOTEnCWQrRegwbNrlYvlUA6yBw4C/pGn3l/E6ktFnrFlKxn
IoguwxDS8CSpS19jMtKf5RistpdbycZh2Q6kDpVyQwTAKfTFmNlANvi4ZzT1Z+V7
PIbXjmLp+YuG2mLmimaDf8qMQ2G9c4VIIzXsvwiS7oE4CmkYst2kUZvtJxLGALKi
wFLXEjNLHbY8p33xx6b56a7qS7xgqQnONMGb+fClNhVzrp1Iro85dSODWtVdazWy
laHbS2c/mRXzOKDAWkhrWYrvNOTfw5OHn9UeRziHWMjXnIJTozNpft2Z1xhnOB3S
OIl7Y0JZnFBPR9Cnb94VoC+vVJ9EwWSmr041Zb3sXZk66JzS5/O/b1sn4nzj9pW4
+lGHF9Om57FkJ6dF8VYW9KvrXzL8bVZie44+eSQ1GAvfytqHvgh/dmZdb0sWEeHd
0clN6nzjTkc+0Uqz8z3izwOqHx2qj5XJlYbkmSHPlLrdruc7ZGsbMK56nU7n+uz3
mHGhaeYjJhzv0MvtoG+sR/LpAibNw2uACnahcssy0cOV5161lg0I5C178Sg3RQF/
IFb9RlC6RYFkdC3QP28j90oJcD4/IoHVtRoCqH4Rx94/ICd7KDsodIeFgvBP8U+2
o6DAN4Rtr+tlAm1xJP85xNheYBA520w7FlqDjxUfJoYsXgEMAC39Nox9fFuthx7x
/vSyg0DLvtiZr1CR7FDpapva/hwBCOsuieq69b2eBFU+f5Z/ko6hQrdzRaMDM4gQ
eoGHRcEe8aojp7ORKVNsAOAiHJRk3fuSD0uP+jIpRKk5SKTDJqI7AsG5TBUdhDpx
cQyYxdBvwhWHESKCQ6PkQAoMmVcjNkwgtTdOOS3og6Y7NtbfFMUp0Wws4mo2qK3Z
5LaJONjZbdOpkk/01ZhtCuTJrjFSTfXqNOFJV2QcMwqtCeda7csIwCiuWC9w9KFS
ksPL38rstQka5h1ILJdOdFl8e6bEBb35JFA0zQqF5yFRWE5u+fCYamvI5ghFOyZS
RzS+FUGYDQwZFv+lx060a46xo8M+OFNd0VitH0GfNUZkKq+u78LXsV1/pASWB7ok
0glKQ/tEg5v0GcCYA3mtuEcpzOODIq3RuLecP3bX3nP+qEqVKPuVymEwHCXftMoz
GFfxamJuJMad47PNFt/AGnoV0IoUpHYlfex50byfIJV+Z14rvzGEMJb5ADgDOHCr
bqFLqZIppIpCjPbU0JeVXfuba4wcyob2pvw+zUN9Q2tKbab9mHbD/Zoo3kTj+Qq2
ulx/mM+NdJUDDxb734bRoihx7NqhuorQZE0WQJQHq9ttrERw8NGB6QRDNN9ItN3V
QUUKzkDxyF6hT68TQABzsFo6+SYbpcapXfpvJHMdIN41gRq6LguV569Sdg4w8/qP
eCKAl4eXoXBkq9yO+lITWsuIV8g1M4lC5wXNSziInaMTpidj/YrVc9sQQBdrd+Gb
gyI4gxR6cVBLihZ63RkJgXx+cOUrqrQZ62HTO5MEVqNBUWfXfKd+sPkJofdMF08A
UMSt+glSHKXkzUuuGzc9j40s7aAXHTGdoR1Ftn2/cSd3eKil1IbxPQcx6I+cuj1L
BJRjxzt74cHQ72g/3daqufU9YpqAbjhjXzZz8K303eZl6iUDz7dUDAspkUAUdQLu
PRYPIXI9IAsD7KZXNELPLW+F2U8G4JSder/224jUW6sbO3Mx9lFxoSFsq+wAA+71
+VEGYkysz7BB1idmuwllL3Ig+qV824XNhqIimzcyn/Kfv0i1MV8YV0MU3de7KhpE
7iWoVAascxFrOa57oXQFucGhcV9sMx96XrfZ3+Fy0baGmZ5rhXYsb3pSbtNxyCR+
E8OllcbRBO3FdaBxiLmTkZeHFP18GX5ysU9UbQn8jEk4AUFgVRGcYZyzUFDsi1DD
NhuYGEl8t84ID91ERiBLmjfUgFiEZdZseYLEDV51XMY5DJAUbocg2BIF9aF0iYlF
XkF5z9lawA96sFHiyHLtU+Lx26hQeGefDPCFQvRPjIa9A4VJKGJUZDh4+8OwqZW0
HLL74VJwHldKE3r1hXWOSK7zpyZF7oClONNVrTAWmYiRYDxZJvbu+VRKlDZU70Qo
CYMcxoBs3YxV+Lcd447RjuLB45ggM/ia0EIrHu8zAz8Roy+SMSm1l5AXOuj0ukCS
Wh1eOE1JpJk8dGlQUWDNM9fxuhw6jHubI5TzBKQCeBfqy5w+BDAFR/kaQyOqqswm
dD/2TeqOQAnThuyN8f4Xy7KxO6pyZzd0dhkQ6nWl3IAsS6HwU/VdqwYvmmCodvH9
EGmRelTbb4+FiSHV8sv8bgeytWAlLe84kDd/SnE/AKpaH7engJMtvMWCFiOL+2/n
PNf3Ib/pSwPTlqXykMVvmt5SeMR569+CdgWXD9d61ziIRCWDM3KNuwL4fYdtluFc
nzH0yxLroOO9nVBAlC7IWcmYkdqiWmXgEIzeFhWqdXIkU1RTyMIvGJDv+9g/HKAL
XpBz+sjVOfQE3kfIhtLR1ypXy43yM2D+8JnRuMo/hb7Ig0NsK8ipzYFoJgCzmqc1
rWx++ymyooK6RE429tQAKqGsOGozq32ma4QrVyAH/fCpdByw1BQBzTlmP6qzk6g5
wApX8d3q5wEYi7zJPY8PJ9mpwNuMinakROmj9sy1lLaDblcWG4GRbv+XJYazcex4
DQtRspAAnMqFy5MhQEwRbY7f0kiD0/KJU3KhGPyVv3x2Uacr/5VgqDGSaf6lWK73
eW6FVXBoDRm28WlTunjB/g5IPlWQvsYPAUQG87pncA/WOHrSYjLSJKvSo1HW2B3u
rmf6Jdqix+Y66UoPSIDEwXWtLjYqbTvcG8ej9tAkHNlPmRDrM5DqHW9ociAjlHLB
dwBJNsTsYidyW7CGnz42r67EW543Lua+3+o3RcaLTG/9VICCAi0MogNjvXf1j2Mq
SKHw+pvcQ3terlUP532tEzyr/Ow3hI3hg9tHWdFV/wVvP3aF6zabPnsKX4Vd3HbL
0gvs+sDVTwborDLirGOrA7vuxvquttDqiqgND9FC95icHFg0aaTLzpqnwQhrnJPK
2jUmhsqpD60/2g7sbooKG0ZnatoKbqx6zJdqN0PZYlJejiHlfDSBBEdBZ0ojRgY0
oqpXq3AjPhb+BqAwiQM/GPUUfVBH4cAEgw9ZGrWxKQ4DkL3D3Ij4aoalCTp5Q4So
rVRtyhIEWBG8c8bARJOGpAEpYsF+2skOFPg0Bv80eRVKYVIxvcl8lOTX89PEJ1hu
l1/uygBcrP/VFvfxcapuKLV0U5r/78tV2FkqfUOUiOkvLY+yVsAOTCDbjKwZ6zOA
oKbSHOaAu8RdGMTmkWsyq0xvdU3abMALAj7CQ4e1Nx9F+Ah5CBtTrzbqv5wGOc+I
LpnAaz4I5e41T6u431yt+O4UWBcXvf2eRdB8/u4xMIVYaADvjwysK5kIoGMh7QzI
2Y5K274i3+vj3rFzqEvcRuMtco5Uh1cMUvAZZfgS29Z0fAspFCZ9b5jNNh1BOSdm
DGWCNFo6ZbLGIuhIyhCmF8lqn+CMTy757+Ir3AfVxCdkztRW2Vk8mmPEPtrci1MD
5yP0y/cPKkAIc6v/orYSaNPin7CCJXCXJgZkdlKrdsiDZjtwesK4pI1585XGzIpz
xGZzEKOThifwTsX2nWf4jM9OnGqt7BQ1GPrUsYEzM8OcKeO9LAKCEYSg/lBlN07q
ZJEjFluTwbHJKKcsabz2vO/rhGdasAVvHq/ypxJAbKURrpyln2NpzDBRzQGa4ibJ
Ei3KoD++3xTWlBoXFxDSI1QGQOquXPe7ck7i+8KyWv24GzQVAQf6kLT/RAXy/h7H
eWP/fPzCRess5/ArY2sE5vl3pWBKqgrwU+Sb7+z5tVjfroMSTi34sxuAdaOMfNTu
BDGyWegAxASWW8G3IH7JoELKi5aRSeH4n9AH75D8W12S+4vDWCvGHPxXt8oU4/Uj
ylGokqEvyhHaISikaYQ5bxeGCEzUWsttEoap2eTcYl+vS/BlJxLgAppvb8tvsrjQ
cVtUA5Odx8e50wC6MHn39hCdgaLZh2c+DaAennOJtX/sOT+/3aFtHZYBOENLOQ+4
NoiOesR0fmci9YWt+XJWk075NKc79VcH1ApqYy27dYjfpbnO7weESz1zmGwwAXWs
/Fj5d4A8A8t7SExU/wjM7Ts3TcQK+h7PDOMJM7YhFa0O5OZKq7jE81St++NfWJnW
uayom53joKwbpkqjynK7o00iL8knt+7fPZ5TAcWB4MCM4PlFm2Pj68KqqP42NbU2
6Nil3lKARGZtG3pyJH9Ji0tGfbPVypg5asoUXhgue37RnlT3TG/A2Bw1x9bnrPo/
2opXZCbAop4+4yTiDx+sBXjWpcHlYN5T2KPd8fJgzcCEvBc09Y1kiHxF+MeVrZW/
T14MByDqB42fqaHLG5r+LBX7OIQrsUSLv7QiIsh6bH12NPbQLb6xx76MY0OEnIR0
8d9dfP41EWVX81G5hIVBqkTeefDkh2CyRmLaWUMpxtwFlaj4FWh+nkj6BXHY1lwJ
5YxF5002yZWoMKBzFvQnUnjbYveEF+cx6AGZxVGoAxeVbQB/RsW3B3HTE3QiuD69
NzYOoGqnyzKVvu254iOwprcHmfrlUHy0I2wMvALVNh71uZn6Kii8mH5/IJU2y8SM
yjolHFa3K2JyyKU1QONF9tPIVdinuTookhve5pMTM8UAnnrhWIkbGAQflcvNx2O2
fhld4HXLevA0Q5t9Mzw83Knvia4dOnVaaNbCoBrjIP+xiP/CSvh5zkDmXJpCwkcb
Fgg2aNIwi8+DnXyWBu5/YC9seEdqT2Eb5c+/mN5phjQBpaAb2dgA+VIt6fKQbTWk
0QUtXkcgN84NWTg3rT2Bk9a6mv4kMAcw+V8EC5taJNuOiGL35wlsmkAJneDoyuxr
xqpB51MprvxrK0dcD5FzLR7r0KGvGesb0+tH9Lec5aEd6rarZwzrxiC3S6U6mPW0
QtdMxECP/p069kNHtcxSgN/ZjMMlX4IfN8Ptdek84PvVVhHaUB/QVlQmr7jIp07a
51plV/svbVscMYBGosCHcPhqbURPZdv+jdSMZ2qoDZhWcBNPNI4foGMvz3c8qjDC
2lmIGYWTzxbFcoA1jlUbOJ0es5ofk9ikkSObWQJF1XmuZP7IEpk7nNtztZqdPH9n
HkCHFPvt0bS++PSwvuH2BCZRJxADNcqC8H904+VvANNidnkLpVEhaASdINIZZsEK
2h4jh2hll6FFk8TWce8vXKkwKaYV/MJcxRhKyoWWBWsYZ1ZdBZHTj4hKg2Bb9y8O
lbfGmpx3FhvCftGUweN63ySpmjDBb7DgGZGuFSmdIQ5o97OuWud8oUhh1CiVpM/m
tZmUECQU4Ho1cP64xnj3M0bIEqDnECfygntr/Ax8HyiWocRrZnuY+eUx3Rh0sn82
26WGmyVp6lTUl/5ED3uuj25z8GizC4t75BxX1k/uOaHvlePGvt8QwP39kvwGQC+j
MvqDzjqlTVh6KoG+kNQb15VvJARKz7TLdr6UuNzGTcX+/w/e7KLWRjXgex6SeCLk
bhfjp1KzDSms+FNa5XmZrw9wP8+ENwFxs87jAbbbH01CTllYpEORx1dlstuWu/vP
P2gvJr3iDx5kdWNbvvJtQRtYI0mu+o5XoatwhwJu3+uGCFyng36uYqESgY+k1AdQ
DoQMmV8Vi01Mqy/rhAY5Z8QTNoVB7P1UDtGU+bFFA6+THAtgW4XiZOIx8qu9WmjA
0hC/x3WgYOVB9rYjDbzG1EKQi7HfsXAvpFG9z9XjxANEjjIv7C9SmfBjgIUbPyuX
C6O3mx+hrD/PpUoajR1/++ecgNNNAcZdkSCp50x+qeLX4Po2AQg/xRaY+En9sqEk
/WUJ606YiH4rIpXC4GVxSo8kQMkRLVWCLi3WUTXfCIrsEyct1x5UnDbPkmqWDtOF
x1ssHSyY8zil0uMmXOButt4Sc1Nd+KcQIYoldIyvP0eDmG7wsLZxJwrPAs2DmLk2
eCRwtFOOk8eXmdi6/0FIbYQ4pKWhoHrG4w9DlV2oSyy0QJ+wDo/+fN+KdR8hCedV
0NNVHJflVM8c4ejXhmdoYMrLzMHiasOuv448khUGbb46NhgQ4CEukpojE6Ha3rHP
Getr+xHC/+EDvuig3mbL+7LQFFbYT+dph8QbL/phbqKU20wOwlYHgiXS8DvBViHW
d7DRfEBPxKI9Owp/CUKB6T7B+UP/EzsgixwCfq99qumZgWgN+zfJfIgVNtHM8dcD
Y26Pt1y0b4U2w9AhxoExu7LY4bFr8XlhcX8IHOasSR47dzKuxFqgBTQkNBLbHHrb
eeCLijuK1tnOqTdmFwSog4InHN+UX9e9PC0kfC/8dwhfRcVgSNJUAUv26Jl/+jlx
QzjwHyOa4fANbwPQIxzLjHZuaMkWcQaTHQ9NHkLDLpwneGpROaGAVEPavM3MPK2i
m5JRS4xhen+5IaCBR+TQLoP8OxTB0VCzjByUk9drTTuqNw8CGtor+YIbuw1Nw9pU
W/+XdXmZZrj5qxhmMSEGPYIwqtkwTsmENNOYmwz9ZTrAJs04Uh2RlRF4xxFNfdXH
QGD/4mauKdTXMYZZgwZ+Q+CZdiXSRxKetPxkqDkEUNgiTBlsKxc0kyGn9HQ6+UwW
PcrvsdosUx+ypFn/1/B9Mh8aC3qzTBQTjjblXCz4aQcQOh4Q2E2qOWq9NIiPkAaL
eSei5GN1ow9S+R1VSGLz3yOCPfNUpeSndwcAWjW0ntIu3IGiTVh30QO6Cwj9F88B
SCYhPvlIwgNtLA6eFJgoLKxPGxQ+lqQMRAwvobX0b9qL7l1jG68FLpRUJj/4ZB1H
1IDm6W+GLf+J9UmIBBERgqolUMd+ZX4PzGeIQHYulZHzW1wWSMG1n305myfogYiY
jvSoUqi4B+tFG/9cskr5MTNqO/fpA5Y/6sui8DpRMvqNJQ6hcTBxPckM/w1WQS1D
Em8xaMk951bqMaQkBBQR36MgA0DfWN+yDeWPCSmeEIm0TUtGGKGJ4c3Xjozq1tua
71U191chHZVJm9UzBoJnEQcRcJXZZynPbVhdbU10ueB1HQ+WcI1EoIyrNTlSxC1P
VaVBSU0+OepU6Ky7Btvi1xyH4u9sJqelLdgEHHydPZceG3PpONRzeQQF9Qx5khsn
hCOeIQ8O6LMJ1O38cXinVxHs79OiZ7ybkcPLJ1zeX8LsQRsF677VO46nmZmsX1LM
j1Ow6ER9avanlqPYRgbjqhGMV85KIf3Yvwu1LhM+ZKjNXvr2pdImrETQaG74/qzJ
p5biq0fOOpsef6pnNc1+nfp0Fpye9C812Zvl+IWCkbuwvfJd/Xr9So1UgjMioaGw
bJfb687p6f43w8+OX8LZvcnWig1Uu8oaEcAeS211/DJO0+LYG7FrUhNuEx1LfoTm
hxfx7F/vq67ir8e8yjUe9RopwwRSwchL+jYyamXpAYYafCgObVzFbvBzizUUF4+y
gW5iptuUj6r7pHoRrDbaP8P4h8aRncJrncyfhxTKdqhEyIXDabc6KQdolRbxrRbJ
sVtkf3L0OcLrnciXm9DdiDTanESwcBwwhZYOpK+lhqa16bUr0FW39Izs5+hNk0Oi
LzIIgznEakZQRAuwa+Ub88VU/o7TSNfiRztuyYEOF/lcfjjOIH9h3W2MenH1TYyA
MNPXRGpRermookE9ND4PmGCzOk9LCu7lgV6a1CUQVbJ4jMkTSQ5Zazv/ewR3qakh
AEvsN/tYnC5lTiq9uyBDz9Wh8cPSBPl3WDnbZQB71PhIkF3mBxW4q83PKQIwLV5t
PQ1XAw5r0hXpvlnYbGqlVyikSdEPnd9xrVU49vLTuE+NPHsc6E93fP5zaCg3t08N
IG4ylm9BPWurNTfjU8UKFcD4QYYi43rHoNmuI0YcVEqE40zujzyRuwOSaMeMyfuN
sdfyOB7vtkoDdsK/g5tYwezGB7HiFm9z8HFpdX6/kynlGMyzZ4rKhegyOFaT/kMX
KbLoTjOxQYdK+/NfYPf3nqbug4mpzgUjSpYoIVQax0VAQvCx7fg3M6aFhQR595sR
NMhELUlDHzy2MIIWyClpCRmvI26aGdkQkstes5A/Ofo7iifhTd/3LrNpALp2j5qm
akZteFKA9rM57quQdpOOcHraRH5f5yNWZdpzYHZShgnJkhUClmBsoD//GEE3WKnC
e92FnYicnNugArB38PTEazv0gJ8szI69EEHWf8pcetuYUB3o/7mkVNbCv9u4n466
+47t1Xvfd3mUdyKHv2xmGH3UMJX+kYXyZ4NugqL+MD6Mo5TYlD71MkzcAfxmU107
+n3DIxMLcXUYi2cnkSZN8sgx3IYDKVlFkVGR1oUkC+9QRgyGuCHOeMbGhTvBZ4zr
UzkHYUQdTxvD2ISVTxnG2YYmUVr98n4PNOhudZVuIYa8RA+a0KhkxkUPqULoHa81
CKY4ZGF4Zh5ZDo4j3X18mAJBqByGnnT5u7cSgqxYmsOnmVEgPS5RNsY+HLTnq6TG
Iay6+8jFHvvKLQjetq/lVWxs4bfuvqHEcexwM6irdwkuI6MyRKiB9IkMeBim25Jy
tEz3f/7l54jHb/M9VAqBlYT/Zy37aCeND0Zc0m1N4dYbHZKkw61h83ai2OQFeHBs
iHTXoUe75Rnxucg9OoGCSzIvKwdB4UY2qWpyYlxBkdPVcne/5u/egke4fALVjzE4
Abe5p545bJbh7V0kxwrQR9eJy3igKfYtNtTvbEXBkthMYMmxRC2pagMt4DjuarR3
UFT/DgzukQhQhnni9Wa6ZLOAKAVDe6FI6XyhXFi2H6iR+BVodNjwtllb9KXhbiV5
IcUZg+S3XgTYUrvB5QusBS3BCZ6HWmLdCjMB4ELa9xtEnqI6C54DRdUg5ltnVSpk
rxcQs6SqeodgVc65t2ZdUvkmythCxSk2W4ctKvocO9sp8ut4TH5dAhEiOJtvHWKb
jbhVK6V7NqjA40xtRpUfw0Fw7Rd8w4ZqgsEKFuy03EGIRzCGtpIzV8x3LxD041NJ
8Mp1jjko2hDWPXGpMYYutvFsJ0Hv6poskOHSMAqnEblsX1UQPJVyKmuxTm5AZThg
eUdtxiubdZ8gTljUCDjCZkfJ3HUhmSemQsIlBL5pgXk5Tch3CFprNe8UePK1AdxI
AWlSfoSFqS+LSJNkUaEvrYTCevDIaoHesSx28wWHKJMZFiUKZZklbNX5R9FUKJi6
g62+0fmAJ2dnANaoV7tYnjWotIjSCE0IiDUyVSb2hOswgazLf9yTS2UJVF9fbB99
NhQrllLb/tn6upRWwBrsCSGq1ihTu2PKbP7d/CWioeb5OBP+c+wPICwj6UjyMKII
jCOQAJw9IakLNpaQl9KFsnkA+pEOvx87QPjkyPo4zWKKI1UJBEuwAWkPU2p02DWI
paqOqE+guof5TNA1vjUMuma7ZFRqj6/MjqMsH/0778rgssTEqCUYurxyQj2QKclh
VLm2do/MttbQxKwPQ9P0MgafVB0Ozj4CLxrV8+6e1g/JkFB6D5vRE8WRN0aCQ6FN
jYz2ygYbe6ljXfTLE4ldzlTIgG0pv/3tDEDHi5ruM6ZPEXeOMrtVCnJ9+F0jr/Cc
8EW2FVUDEfWvrPACYqHlWB34gyP2HjSHWyImB1o14pcLqT3MNF7UYRRiXlXzKnKh
/EM3KJanEDJcmaefzCpd3S/HkW398jFViyOYdef6DjOWzQITzZzzb6iYy0XIzWll
yrjF3vQ55aDLV/vHq8qwMav9Uwslswr7DwIAsidziI2pF0caK5HoyAjmN3h+8OMt
9Od3uUImkTJDhRh/WqN8JZEJ1Y0xZn6YNIrNQsn2ruLaJXr7537ntR9HEZqZYjQp
LSIBtmupmHn8iV0PnO4vsXP8kp5TVE9ALTB80lueRtXRaGHlhkiVmxH1qY+5Zhns
d6fgoAJYcoLOK7yzRg0vM/yjvg93ohTPPY7+JunWCX7FdkNdrAgW9Hi3k/TrJMhG
1RxpkqMxN/KsPLHrb2Cb8XkLeIcWvo3ywHAATj9hqqeeIBuSjMo4CaLlsMGtlBIq
7qdyuEFeUf/E+VR+Mhpg1AoDwkOXAnigQfuwHh1Uty0bFCwylBpQtN61jKnqG+me
rUhuZ0Xzded00XJgRuE2hTSZIE8HFRZZ8cs4TSTnmkuktzeXjs6PTmFeKF5vxlJe
2pUmUXanOozGkij/qlWXzlPJHnlGoByDPrqDnHorq1AOm4zewztutpwJzCbxy2ZN
tqo3Fq/pRxM6qv2EvYrdisWHL+y0VOl3WzKOTVADZKlKGRCftFdt7wnbUMEEWkEP
ttgwc7HBHoDiqUGV7vGRAROlalXN8YbmXR+0vBetsrPjEkjbxlTm6pQoUoyJO9er
4fxxm5LKUYiYqU8RD7GAVr5JDFOZyGNR4nC6r002wnvMohyF6zZiIP7tlHpVlaWt
qHfF3PQd0HDzfFEyuEt/B6fRxWocv3W9WAlRspMchAnuQvPnSoWUM6YRSXqWHJUn
VzdSAHOgzfEAEO0ku1fOYsGrpnhXtST8oqPDUWi8QuoMMLHsueL4KpyXj0Ghz5t4
GMlyVN6PUesvRAkrD9qlEZECx2VRkYlpFzv5kbvW5Y8aH/uqAUqwYAccBk9p/omg
jvwUeJSiVOsTiis8gsY2Qqo5/4f6+mAeZJ/KgfJbogyH76TXmEEVUQxoAxykper8
d2N+tL9FCfdWfjgv/PMMvHqwlWcBjOZWXGVEQGh4rYVHUxaodKXRwYN1pwNfbbew
MYHJ8ut7lvW2B3QanU0VnqgkupavV7R00KDb5lHfRlzt0d+W58iXYR5GXBSwzpQ5
A6UVWvBIJGtYC9cP9gCB4aHLYnndQ40nmDjD4yWFugv5ay4EnHEniaiYJ7t4RQV6
AdzFVsYCMbA08UVSYf1N2DXFAqcm8BkkDYSGo8Db5S+mX8ib/ZSi3vq+G93RKK24
TcjwoewQSUomCB3VjOcbNfpX9f2EAF+ORHi0g9OaSc9KUUe2jCbP2TmJ3UC19biH
paKpaytO508qNxjIT6O+3riHsFA5PjY6I3pZqQxpO8Mp3uWb4svWWyUFoHyss8t2
PCSjp5kUEAtF0360mAFDFpj1+zhreH+XSFMM07CLQurHXEkeup193qfz/UkMOuUg
rjqQcrpX5wwCRMPgcND7cTH80XZ/MI/McUuujOxOneYP0OUWnGJQwVnT4IAm7FzE
2eh9kZ6Mrf7k+0/Ponc0nIRXatEqLHaY5chQSbCSyEjJBy/0b0TwRtNKQtKSt2HT
GtoYllxYTsHg0whS3bALjWXXG/jQk1iLFENg+eFuB+J43Ql06Nz5+Zh2TTowcw2b
4k3Q6/pyZAl1o9jJg7lVZAWRwPkRmEwAP84Zx1Pn9WgFUBYuCfzQluitUviQ5yet
+jzwQp1cpxt0MFkAfiNOq+EMN6wphLtRXBltac+h1TQGYRE/Xw9073Skt0Hur8Mb
0y0wzuSwYRGHAlgfr+bMDoc4jMRxoZdQk0O2FAimaJ4c9vUWmx6byWmkOcGjCzuJ
I8IoZfffBxDisp2OUdS75AZOscWLizlW5s+etYv9nDAH/6iqWzlqTxr9DWZj4XV/
giAqG2pVTkEg7Zc67Lw8iZhPZjO2Y1JbKZazGj2oZURMaXo1a1f1RJmXQ5VRDJs0
gBWWytlxxhGv/00RSmlBSi+8Qc6mD92Uqx3JobPegU/ISWPyqRP5dLe9WGtdLyvW
fmhf6w4uNlcJCoM7l/9MY5BVF5H+ZxvGkEBs6TmxoVBf51Tswv8odaNQgWmxDkhR
a+GM0cQbzUNLBXzCHLLF3De6PzY84JaYtO/kdxvmTanlRi2Cy33xf+oqen7VwyS7
sqFs1Rg2xjyAsliZX5CP1NBCccO7iKhI/5+CtcnI94rzCc/HW1534gB0m7QxiGca
uVxlTsIz4wr5jvTnUpVJXiKqoybNFf+4A7chHdI/DuaWf4+2yHFuOT9h0Ycc07Bd
2amzNB4/MToZsyGZtOCZtMQGG0trHdHQtYOXTKKmkeIGzXJh5bd+s4fEsEGT8zct
C2DKEFspfBdYBpfrBjyf3FQwLQL+eK6mr4KAqOEEQthRuvhvuv4FqXyBqo3yrxUm
UdAz6HNyUBJC6fU+3gXApkH+suqSs68DpJY3WTgbZkAVTHT8mqN1YPXm19WS6KIx
aziZg+XX4RVgwJ5hUrn6mvqpn1jvhcC+mwTdn1rznW1UveMz3A7nRzmBWS1tNvT6
8fmLjj4JWfqJ2eVhjM5fF4J1foFM5Kurpw4FJjCHzdyInJsxAuDlwbVe/q3Ziq34
gOgHdzGPuLOtY7WrHMkHLPMohCw792CJ0CgvbamhW7x4opjqf1JZRmAntKlm4UAF
d669Cmmre/p8C6z9WntMDxHA8jXuCEm/kKa0uzMDsXLS7efqGJsXkATFlhtOQgl8
+vjvtp+ODFQfQw+eBTnXL9KuaBRM79UFTYNTzz4aHnfhgGWA9M3tS0TxiO2apX/Q
BR55dc30IcRSgC4OgnV9jqeSOB1I8JNhO9c885YtQ0/gdonevgnxfpEuy2OJYxis
FYFs0B1M13rmLXyxCqwdLmTbCovQb0CSMmAn8Z84yetI3Szve2HIxy1JpR58w7vJ
yi17As6vlFbwL7pO41d4YW8GnvZtYrvpq02WRFQzYjlstpRQh3O7SAKMh5b9mBzm
+DAK6YNp1YFN5xit6smUlHZFiFVxCVlD7Jt+vDbm4vuQt8diav7bB9krUQbfbLTW
o+O53ZQQcK4eBRMicINaHrCtYcT5gvQ76i0917Dinzw/Y24oK+61GGOw1FvHa/gy
3b5jeCJXoLtK/7lprwopTVHtb09JtE9NAmCIw7WE0Usg/ezyu7uRaSjdhgq9daQ/
V7pUCrhx5A7t0VPsj9kjOzmsRfOnyzzqB9c16FF9e4+eVr692ho8icL0nSbwClBq
sXqrD8jawGO65ON5I4rxB/JTHtiDH/xPvMYhB2gR9xcNaYuvx/SvLOR/h9ryzdfG
zjXm6N5nD0koYkuhaXvuhiMMV9ug4Qyecc06SMs4Sxc4d+o8Xl3OhhzPNeorPB+X
zigIg5o5/LYlwxCeICquiZkASAMn2gzbxkk+z/k/JFIqKCWfznItbSKq381PH+cT
0nyuYdv144yPVfGTfhdndyN/Lj0Cqm+byPRqni4DJFb1Cy7pmycIl/R4aqqhAqij
GzPXoDsfrVvQVUwh1LHTQ6FEhOJanEOHnk00XpPORfCU8YcuVqW0qj28EBqaQVuQ
y2Qo0EavGDs7+ayApO/Hgxk36jMSi9y8e+mAwq3ulH4xqLoBCVl8gPQVJlaXKGwo
XdhWUOEFmY8TL8nV8ojW0XLni3K4fKuU6YNr1A0srpa0//tjbMi2lvZxKL5qdxEr
VCYc3HGf5PI+fJBGkmJB6KDiIwv4cxAceopIc6hYgN0BXe0HsuKrsR3BKMNAVFPk
iWnSNaneW0/GlJdkshl0DLsw6RSjpi9/iu6yNqtIw07hfKmdJm1BL47DX/0zE4R6
NpJ2abSvr9wjF1yuwFwvnII+UTIYmGZgCDpxduUSPuqxvWcIF7nTpy/Z3fIjKs6p
rq+HLgM9Iq8G1SSxBS7FLnhsHSv/cmG9L06zn8dzrCM4/6YBhxZwNWLKoZiTH2mf
VTEurfdLqfFK8W40PI87bdwINGbWBTPtPm+96ErNA1GuFXsTzaQD/FyPSKdEZ5Ra
1/iIRiKSjWHYMbr0Sbdd5CW46RVCEydfp8+/tv6ybei9qkYL3XggGz4Cs+DZC2Yf
i6Ou7KjBOpgQoFhGqKi4zO4527TqGjPFY2Ag7vojeM8TbQQ7PxsiA1Ttba1U5GUH
OzTcVtImqSLoYaJl4kIqt6eJ4I9oIZxThViQqfzEA/yL8AmbVIpt543XcB09u88o
GrQ19YvU6LA+EqLe0kZXb6Ad7jhUJQ/KmSbcox1woSG7mZmKX3PQ9/nam8mgvJfO
ZKeprFIub4PIMG6iWxoD33IUKkKnu1j4aw3Ntrx3PB1Jjo4L7w3ZWsn4e+C9oZpG
IOeMgRvxibMzngxSdLOvDsITjPmAWwvz/HE7PhTlHlqrvWiWpaEDmMah78sOR/nz
C6kF3gqlgfHezII8eaiEh4mCAyGYZW6dZ73X1PsfNPpSuMvnaYW4glUx2F37U8rH
GZ6fOUc65c53CDGe5oiQ6H4I8P7LqvMrTghzZ8ODEzbrBL2aqT0UdOm6GKpnly2k
DgPdgVX3HmU8RhaNMCtkIX5bZsYvZg+a9xv/olOJr7s07kOr1p0qDSKzxsDCODke
wAvz4DoQO17UwBaKRPk4fVjQqb3mt66fGDWrHlvBMpMiTlHdK/2KmpQJMbTgWhUn
J0zYS6r2pSwuC4CXFIZbB7tVk16GZoKAEIvTMOBJZ/KKGs78jeIl342bGuNvgIdt
9f2p8JbCK28/8/zjSdiCcxX+0W4ImrdOOsBjVZ7V/94+81fFO8iZcckYe25wvSdC
aSmiiUdkDQBdLn/+/Rh0WD0cEOEOsIcWQxtpYSMD/ZICtSqrQ41RHokhRjPfF9QL
2C6FG8ZS28SD6s/XW3easwfK0/iLExOwln9pMxoud8YZ+CKGmRJJPVWnf3PWh+N2
rVYuoq84wBJH0Hw/f0oGBWb26gk8w7J6DG3y/2JtTREuZzlGblPMRjy3bmXkl3nE
I5Z1WLQNNo9TxSLRJ1pqfmL+T9y4OqcOp9XBcwJ96HWiJ6xOayKPeEY+qsdjqq6t
e8MRunIj7+rbx7HMH9FivZJLM1sW66PCch2fOE2xzcfiZm6ErOpkSJPnEvJouRy3
VAJrOcJbaifKpqGAtA8InJzENbocX1ckqj9Hl/sQFsM84Jup3+1Pb1bkpsOQ2Gat
00YSgAztASCf+6cTD76YgpD2br/Fff4+G/lW92l5xEcVMBOUfnQ0RqISzGCALmXd
DhD2CArdy9mAlhhuFDHS527N4nGKAoz6FtW9AhxKcgWB91etyAhb71tki+ps8OUM
5G+JPIYx/6qQU5iSwfsrX8Y91Qrk83+pkF0h+p5tX7Fxhj1Nfvc+WH9IZ0xBfMt+
YNS3plM+JXawZurPkB+ONQA4l5u0YNDcAr0zTY95h9F0bHgESgQni15Uo6Rv+wnn
odIixQUfzz+8jD/No5kqoeU6Iwpds571dDH00WdPDM42PQt/BpL9laBALngZnQ2i
KaM0JEB2WnHI6ogKWn/bN4uPH1gijZ1Yjb8JNNzeJ06/HdG2IfcJOnaCl+ckYfCJ
TqDCNP23MlmZ52cGMfHRBt45bfZw/gXTA2q36sz2aTAPPf0Rgz20WhsHQyXbbJqb
iHD2C6GIulbcysDbTxm7yhNPPlFtvLW+UgAImUFnuTexNi4OI9el2pQGwUO98N0o
3e42YsJCYoRtei/CDY9F5GI9hYxnR2M80GGNThTRSviq0QxLsgSDkm7MXEPfzjqc
8UULUsbtwRt2rxYbEXrtpS2uEBx4yO0HN1WM54ixPeiQcrbb6BOfgcnn/ZBFHhSH
VGVvmuyEyOmyGhWoCFHwGSeaKMuoAuDFAk9mlu3F3FTqm+CQxZH4uDNGUISI6aHV
Cp3sT9ScyFlAtqFoluQ4PvelaPhttb7B13y+zcxoP7FBqdwRARGEqGpVHdigdDa2
ZNUjIKR8YLT3eFGV/qly87TosBcBabfrs0UIMjcdl0kZ5zuJmoLJgS7K3sUXdu7Q
z2I9Ti8DrxQrlrPOIr5mbnSFtoJ3/spvr8ZeIJq4JIUpVVatQntvT56VtB4HO64+
9buIidNkg9Jpc/gQR/TSIYhFUWqnR1PjzNc1s44D/KzdA0koGWvk1IjOLcWBbjA8
bKdpdnvgL4HQ56MkJ2ldd+eIJ1VBphiB4ISvjq87bSvov4m9T/C6OOH0vBzXnS9k
gKR635H8FAaUgENAiGsFPZLAWXe07lvScQYXNTIdcr9914JylLKDVtOY5v7jin5F
GL9bQ6aYYpnjxpSn2lh8qDv8PL2x8s+juf+wEIYvIqUrB7vQiYGJYRh10yBErcEI
LL/G4CeI1Eah7dWfyonBnaGnaS32vXXPaOWCuaztUzi08KoNvNF313hGAtxOb1+o
evhcDmKzWnOmDF6IXROFFRjBAUJzoZE2JQQYlcgqlBnsVs24ilHqXX+782qR3ZqW
b8zGBkW99Y/mZPX93ThShsgZ9IUfSuaJf91tw2aTvySoO1CM7F5DIcwmCasJkEl4
wXM5GqmH48n3EnYSVeWIQRNZBwlCGuBGsibX3e7EvHWGBp5dTc4FgxBcmGn3YXcK
g32e4+/yVTCzJpY/dOgDafVTEmrJZhAgPmVMWZrFQZZljC/hdwSjfCmWpKVrLk0K
h0hcbEiCea1rlJeegu/H4w+x1gOBr9CCm/xKqUNl1SYLYSlSHgNCqIwwL+0Sk3vq
NnSaCfgISG9vM8XtaafRFzKsRLDS21iy43i5eueMsKOGR9+yT8UIq5HalEfSnC/k
v5b0bMCxqZMuzsu3qVIoPMc9k9ORQWQxYGze8Z/yx3/pDcjxVVvWbcVGWX2CyAX5
MG/JxZF+4sviHsS0/VknV2LlAtCEpwX7MvUSgijRE4XR+Q+qyqE8pV/zISdDom/W
CiwCL3Y1wbYGNPuASx6YLLOgAwMgeAa5G3goxBb1q3EsnrW74O6NI5MCCUK606Y5
eiRWnzrZzvq+6lqV25gKpfsoFCYQqW09ZtG23iaYHZrheCQUvnuEBvYqrTGALw9D
Iy/EgD874M1qUg9PGA/qfwrM6FGh9RdCsA4eU4XeVobyWhBzy7W9wXhDNNa464xX
0nDBL05fBb/4CM4HQdPGcPpl0VsKkPH9WjDKiSphVPxhXO3S0ZV9Rqk6ek8Gk9uP
tINc5Sv0VM5EtWDJGwLoPf+bsYbQrRcDyM5/4qKpUn3OIm3yZIMA9bw/xUwb22k9
ZA/bvNBGH/95Ptjk2N/XR9F4sd7J7nZiN556NGbPXrq5pIaAfgRPDmLG99mixY+B
LQGSxLXPlF7hgMZzklj+ze08moL8v7eonQQCV4vBxwkxhjuSSnnSecV4do8W5ki7
lIi+nFXpif8INKc+wGsdKLIN7GKF1uJHNtuys1GziqmXM0P84eb3TiRLnMrQGnW0
9YMtJu4zLx3cSjPmR9ayFaICMgRJiF9kbCLZUXQg709Lj8mLli0kIejXuO2sJt2O
HxftJv6PRu0QoJHGqEZUXD4aWxF3+Wi9lvc4Q8Q0hL2T1AxYw7zIUA1MT1OPdq9Y
YzxJsKNS5g2nL5Q/Si/DlZhiZGguqaVk8ZvWhJXSnGPyuN5cdjt2BfhILODFANIV
BgBShRtAUNjfPaO29H8ffGL1PolUi6EfeDjyhaNyV7FNF6QWOeEt1xpWSLiT/izE
8HhrZ0KK/xSPIEOBBsExg82pOG5SO23TFWV4ya3FiXs7Dg8HO4CyDCmVDiI0x1Rb
rAT8ohGpoVlS6ikAA1ghKIzaHWdwiuHiNZeX4JXJfLutemyqlITqGwX2cnGAsQhT
odYMiG/dxSs/fTeohhcfnnDkLW6r6Ip/QPYB5xVQ8sGB+VJIxH0b6lrYxcjgtbkK
ELtdt+YvXjCAdvDpBTxhOleaqV82RIKbD+ZM/LELLaa/xpt5MLmkh+/nRedorsn9
+B/9UIxUPR31ULUuko4o9pgadJN+3PWCCGAVMXSQ7FUeJtMnMpVXjXPe8cHms8Xz
zCSj3QUToY3Z74mFASqLu7BbsGV78aba+HK4sElIZ0HToqYLzZn7plt0+eOE6XxF
GJy2E64Pb1nevzrqY2zc9C3ngC8d7GUx76GfpjmuH40XWgIi4PWLtYWeUga3VTom
1//q2w8aAGUCPCmUN/aPd3wclG9ODQRskimv3X/xvTFbEn12WBQDll1a5QAYikuA
JRoUrbdikdh9vIQQ+Jw4Pk+RPxiyWJ2TcukVO237M4VPbKASTOPYncmREZK5HCvS
+tARC0t2nO6fwb4qXopwmrVhrLwyZrozYdtp2hK4PdJ7YGAZHVGhEkmwpPFS9lSo
IJ4F9Ix0sqiO9N8aHRIT90XU1z5lmCxGZcrwaDY4eeT+co8tSb90SF43+QxdFN7s
1v1JKQ43Oo3L3iFlSNd1L0JQXNhIlfxnqT8aLcLOSHQsFwILdqg4dz+/oW8xlZ80
Jp73fZoJC5n8cNltUUMGnkt195eGvnnpCZGvoHvyN8uuCNCmj++YgDicOTHVHwEv
5Jyr3RE0P+YGS9288gGYtR6g6amJr7XT3h9qNwFuOl+DD2ih4njMisy1E9jaPa6M
W1ABtj8wCISpnIs1A1ZfmAILRFmDNJ7TOxujykR41IkjGJXimwJbUSQLdomk1aAu
wEwvYcW1LUS+dthmBSU7qL2hw1clv6QdDIAUd42/ETyFRQ7CVT/gNJRpHcVxAQ4i
mMx5hLVZVbQrKkNIsKqcp43rqmygUixZ+xEypbmJdes1Mwa0A3fH6QOy470T7PPL
19nBznEsRX8jK2spMUBDzKdQGM+SM26dH7mLtxBH8kTjFzIhV/LFHRqfEnHEBqBY
JbekpdyRO2zWrE+ENbJk5nE1kHonyVD7GvfFMqEbB6PFXEl4gBS347PyLdU6cgLI
2p5Hsb7KWrg24ifKRnu3lJdredrOHpXSq05oLQ6WYUdPcE/tOt+e8HgwsYLGxQWX
RNEZkX7OUFrHr7iGpwk2rMcf40LLKkjwJSVkckAgdl12tfzYfmC62qEfDoel/2Vk
JjOGHJJfAa9CxGE6a0MWp4zTYyzICc8AS9jnwqppVSgRCNi3Js9lzlX3SGtQ+rr8
DfqpTQ5lbUbvrxdXsaKw7VR9PRfyNaxMSG6KhfcfbvdDLDULOQaVFkr9j+SfN1BW
erHaUxd7xh5m65uvTQTp9Z9513FHVulYSAUQMXlO8SNgX7YBnVGYLnixUHQvQtf9
/VMl2NDnM01U9ApnP+Rrc+JCzBKrY57Jwz2Xk0gIB/0jHeguCVvgKJ1vzg9AS+9j
D2U9tUE7Is7TAu97weyleZ6j1zL8r6afim5EnpKgPmur+bINK/DZ1AgTZfGiZzcR
obOv0RLbjIOMAfLHL/9OKyQ34B++BSDgDjGnT6W0Xh0t0GAPhbuMZ9IqXehp8SzR
081cNLEXnjEiUbWtVJFeHJH+z5uzg0e0nYK8567jsAPQIqktgKhFfxxxcHSrX4ED
AsjfNHzse3fG3EsVzu7qXcsa6HJ9OVwnaeVEcf9R2ET1bNxxylzFD+m6JrquT4QV
QDMgTNXApfPz/urJB91AZ1lnDH0xQY6+0Od8KAnV/fFTDZM6XAfbtj+8nLleSM6/
LjndymbbMxGLItlA56NB92+zQSwXVICma/qqiCuW7gTbgqM/94IjmwQ2NsUZSOw8
wu7qfy8fm3J4tf1Gs1VDCy7mCj/+jYu/AzpFrWUIm24ekLmfVpjFfu99eESPE4ls
1+kR4lKy6iEfXtOYtuDMa1CSm1rIIEjVVFWJPD7rgjWS7Mo76Gx2I3Zh6WQNPTwA
LNM0318r/n2+3ySY4Rn8ycbYIEsd/wLOLBGy5Q3KhAa9IEGz5QlLj+6YH85Kszft
wns8tkv2vJHXlNhPkbCPLz1bD9jUpGfokthRIuLq8xkBUnitxjTfIQ2vikGtNyMD
8XQVy9J+7HEtmr5XycL90LzA5faItczEgywmrrH4cEoyijNkjIYF0GddhKdU/jbj
L/tZhopRXET8KY+4ICiclegAz/7IcV9vg3JQLYHh1cTvXkBKMg79LrwSe3mqw6H5
3iPeI1/o+hv0OrkAWozXeiXV2CGddgBr4mDVyXt82811rnUK0b5ohre1Gxvv4/cg
bo/3r69K0oy4ljWoyjPtO3CB+ySwzPVZEgoRcs4RJeR87sPIRVv1LDS+vRfXsJzc
h3p1onJY32fUlpoVniMmTP8G5vdxBRccfsIQ0pripQDx5f7nKy+y7bhD4bwM0OPf
BHynU7wKiNhQPQddXkRmHX2+4MBBnRYzhgDN3Dz1PZinAwzXCPLttwnCuuWljdm9
hSCyarJCntrFGQdgiA6kp2kXkSXPQxik3NJJfsrWW7ngU4LjJpbiZi/yjv0OVC9M
0bSBMuvBI5TmS5wiIs8RVHVVjns0hAEeaok68h40rJnx8k8opb2opjMopdGPYDcE
n2F425oX7L7SKIV5A78M/+dsn5o/gMbgmozXMfTIck/YHjjndv5q40LL+L2IquBw
EzHiTw84xrZIlRPB9FEjXSFyn10/yok2jF8sLintvU4S4CB/udu+UEkEpfvNnmmR
lTX+4c9uxHkKL+Xj8/4Cmgr4Z0a/fzWXUCy+DgRhoKKY08PY8JvQzYM9/sA5Zvo4
Aj9SoykhvGYkVAN78mbLRinGve365iEXWO+/JOdgK6MuEjJ9eXSg8N2eghteoIlK
6VnyJxlnYP38+/5p25ybMXGOJls1wQdNcbG45GBQvEADl7TJ5GBBOlR8C3gvlWWW
U6ZeN1nb01/Nsvo2t8O3bAE/uCPLEsj+wzvBV61en7UQpVHv0qDJDa0jpLEReBfx
iZOaaQZEpIn9f+g+wcudVC4NMllIJJKjnTGSJBqxy2LZkPHMvwK8KYhE4vBsZpoe
+sc18zyROZkxEUy7yRgHmYN14HN4zlo2rQUU7edgNeOcJ/M1t/w3nrSogWx3uL3R
AuI+KGVQRIOxkqrY9CHvcmxiilNUzNQ/fI0wV2EmIZJPmx+DsRlomTTgpxwJZFn5
fsNh29E8EGm56qMY+1xuLtPzfA/2YwhFKIInGHbUtS2s5soxF7UgzdA/7AbhZtSQ
lUTjLoL8upkWpkBvma9zxhfh+vtxgsfdUwq+7qutcLRNYccDfpDAqFYFkF/ky1Et
paZ7Aqv6Eq8T5SFItt3tSPrcWJ8kAAMINaLQcYL3f/rnWPKYz828h630+jZned52
s+wJ/DERoGPT3YHhUjPajzdey2FcyEi2PmT9InbbqnRWWCGmkLBdVDaQCxtvff3a
WFOsAGycsiklIKkH/ctJ7i+ir2n/Ts0khjLQSrZI06sC6vwHRpuuUn/2IP25WwO7
9UEzVRA7YhBW24IGQiAt+3UWBUHK8CUh3LWjyt+IdCiEhmzdRHjLBdDtMaVW2Uf9
GP2ZE4595Z/pYlsBH5Jj31bHyNXe+YvzawXDdEBSf0zlhJQc68StAY7zocM7gBOp
VWlGl2XpakafGvjrtjBvlhBxU7aPahJiyQAkTTgCDknGpMzAmVPPseqfR9rDJ+/K
Xc2MOfApYvNTnpCWdvb0AGShO8Lk5LnXgn5ZjFanV6QCHvkj6FqiAZESuhcXgHOF
/oA/+s4qMkPI7KCeXxPGR+WJ6YzkmFblbUm536naKsLU+Hq4fhh6sR984Mp35vkx
MbRjTSC5O0Ve64xUugV3RA5LyWmea5w5haANpo000lzltslpPLvTsRWAjcqdIINq
Cu/lSgm3v5ZOwKmqjAsN2548i+aBPZLQV3XTtTfO44rY5N1v4CYJ5ht9WXMCZrdz
wdgVU2MEC87isZXI/lROK2CmxvWZJDgeeHu3uf3WYH2nXAv4jmNOAHzvnKpuI1sr
/KdDGqJqIsk7lUbSRRCdMrxeVfTQN6NHoV9wc90wijd7E0DJiXTCRsZmUZpZozW4
Dj8nAnkC962RAN08/yJMP+CN9CODe7VyB38S45gU8BtjIO2LyfUP8pvUVVaUT1t0
OfU9jZaJZ55uwrEt0cWGovidhzOKX+caxkq7n/vzam8Q4nAUkNPZ5gCLaUMqwy0E
MqwXSaKj0RJuqDiD2wa3cOuKVsEOimXuAprxFZ63vQWgCLV5Q+JPpFBRuuGiZza2
e9Ag6Cxd/eLoJ6ocV42g0+E79w6AQ9oPLmb60/qPpdn0jQI1l/pV+35HVpOhQG8O
ObFaHXlFitTNWcCAc9a7xbC7s9/kuJ2zYmSbPvPLmcFANKXPY1HiUOHRC1rExsYp
aNlkqRR/mc590ROf62a2Fi1MgDgrkAgUl/FEUF2YTko2Yy65Blu7R7rIs6dp1bAm
w/NxUX6PlHIqCn5A22D5KDUeCsIT8On8pw/43SohPxyguGwmpi1Ozj8wcfyuMX8B
9AZvV+m2F7EwyauYx37gZoVNRQaRn8Hru1Azcc/QOn+YwTU2z5q2nLAQPpVzzFea
wU7AxbZWTuEz7H2B/JHQ78f8xgWrxxkzEW4Yrazy4WU3vBt32U2gAc8sN29x3Fw6
N0rTk56gQSE6Ifn1kzxEnkk+kz8pQHObjYyGxR8SxKt1QHtkeUhACMIP99tmxMB8
w5QrYWr963sV7Sg9euCo2odHo5QPcChJalyyNVlBVXi+4gygn+fPJsRfkLB3ovzy
68zdEX7BwVqzYBEcalqgxgYCNjqhEjbqg8JwkONER6pV5ZAxy+Lr5Z9N9bWQw75/
SVcpZ2Jw68IDvrroM0jzcgMiwllf5soWj1rLy832ch8s9llqqfnV0MwxfMIKCpnt
I3bxacqsbjOlmTcmau4stmqKitSKUOsF4Z+FR4D8Z7ToicPpcCvsgmROPEFmZGxd
SToI/kG06mEjfQ+e57ABbsQ1aj1ThrzEysenNPCS0tbWyRETT9McON7B2zUvJmvL
Ztq3Szn2YoyHT5OHPA020Z7DolGNLyHMwDrMwoT7xUjTF71efWEOBuKJOTIPdy6R
OCwTAPGApCg4ClpuvsF9PTyJhkDbaAXSyZ5QPIELR2y3NUKHPdTrhjG14vqP4ybE
Jx4NbRKg5MWKi7f1OvhgoPXNTbOmLwMmjFLr4YnCBQmfjDR3b7j9dc5vKqtL7l27
fCuoAYlft/zxteFPAgz7hvXJDst89fuOoIFAQ/cKVZxVn+Pa+CKuQ7izddIKIJXJ
5ICq4doQr2CZk7EOfXUCbyvE9I4fERa92+CStZysreQAZ910ygnC4RMaKx0qBiVJ
OCmvUVWcncp0tTEPXTsRtSR+ftiyu6bHlK4ZH0WCAvjAYFfsPRZDejTklkos3w5O
gP6eWrcw4xb/YlAioDoWWbof5Ge4rEw9gegzm5FR+aY7+unsX6gGW3uUJmpYDeCp
UzWgMvOA/KETtPMdvHj0+P3F3FSZdvVC0MYAK/Gl7UnJLcys8GOd+fs1PxVc12LR
jhHb7ZvVSXIDaHIoFH2e6DwmOrNTuJeBojNqFZn3ZULsrSI2LkVEiODJpvZxnlnD
1rLH2n2bNdrNmVfj2SSDyHn2e/dTduKFfch3ND/CVyGQ7w2NSvP8maFIlymjDCCq
BmDtWPghKTdsITcDw8a1pHoPuWVwkrqkrj+UNP3cAIrEAZrWTjMVlSuMPvFAd76C
blJeQ3K5LWoevwf/g9fODvtxGommvJ6qUkImtTKeR1s5jNDSY1FhTKgNos4IHuTl
Ea8AoJ2Waek6BbF6UH1x05DsMn7QpAd/o1YEmYA2/MpW9m43HuItAno+wO0f5EAt
D+YK0PaqalaRarKC9MN+49atID2XWZpY7pOEiNfdiER071nSFZfRoKN6uY94FeUm
W//b6WcwjqK3wGeLzWpMkRYQCtD+UPsTclP4jVuRZV9AmGEk5NFdRn8V39zAJEC0
YDUp6/19AWr8IlUvmDhJGh1q4XdzqH1yCX73V9cifWODlX3zd62ZpsM1/5kD3Ywn
pUaPCsmMQit2Nijnelao6Hq8Jdq0O+m0yPmpwax2pRETLWkyDUrFNpypMfi8pprx
OEY65sFC/xXXApplXky6AlR6xNfty/cQRDpTnpcl/aXa+q+y/THZ5lavycmnxqAG
LRLorBtGw7yRM5A8U+W/v/Uw28+sBSdARnBcjNn7j5wy9R7wr9t4GUtD41PQCTmM
HlcFNIDDuqaRkZhDZnHgez7PtbKqSAKHJEtnElg6TuWe8ihjFm38of1nz1bEqvL8
ckhFrFVMDJ1uElu2OlW4Y/4DIlxd6Hp2M9g7ddoxf/r4yHFInxXH0V/R+o01GmDv
bxM7+1bx+IfCHGznqV0gdo6389a1i34dIgmvrQ0d6xKGtb+VhidXXrtagHYwprDM
j6AXVFOWoMdGaFsEdJFCNL0KeMlXtLGzGuPzB/Yl/6bD/9TeYp/SCs331RZhwMvz
+LYPGsqFcHnPak8+MtXdBY2uIkaYLYT1m3mxIN+gOqmVIC72CIreID2kZAdSAidq
hA5m8HHlT2eBzHnv90s4TQKMlflFPFtnMiKak20kjhoBsJ6lhK84HfMG6qig81rC
VSQsFMhLy26WKYM8zXa0JQpuA4GBz5CXb+HEM+fxqeMo/GaGAONx1rKgk4YrIPt8
k+4cudjaAmqYgt/Uti9edwbTQE4ZXGqxVSLx9rnelJrR6an4OqR2mYCqY15xz6c7
V6E/9MgFVyW5c79EjmLvJEZdpBO3EuqxgCUeNkY7O+KoSoT8sDxrz7O/mF7l/Etn
FUK6Tc2ka4I9hU/ysP84oO8jWu6VDhpu0VufmvLPGNGswash/++WvQztiUM9IX5T
3XLIqdLQzBygRBTdWnFVbj5SAvePJyNn05zPTVzjnOEOgQBKDCWtxD7ubd3odYo8
XBfqANgK7WFBxaFA+D2m6KNchiz6UlqkrvI5WqL4bzbIvzHEFBIwEQm+PDdKuqAb
VCMbYrnpccRC3ZwHPVVe7XNx5Opp+x0bbFcxZfyohh2YkE9Bigo6pKhybRNLlf36
jpcaIQkiYIyiFkr6ECKWwqG1X846cNTg1AggrayzNCsSgTWeESab+ocVQH/NvLa6
Ui4XKVdHd9bMaVw0Vp0S4XzPj43Urahq/CQn4RqWT4/+bFnA+UXo3cQn2awIxlUF
cycWQPNcy1zxdj1y1YoGGV5yScB1/d4TNwG5Fbq5E2H10lsuBI/m2j8tTLXHikJb
zoGmJPRDp0VNpGDyafYVXfSj6rScLcYAC6KZTBlZkJ3utK4dS+96RBsS2oSp84pM
ImflkIp+Wik0D1zyq/EqHpli7qOZJgWHlsIfnDj9Ahz1j3es85L4sGZXe0HZksp2
SMdxXwm+VRjh/yuOKM/W9/7gotvbq8U6k6ZB31hfno+Q7zrUotInf38du3UjAdsw
57+W2fewXH3vj9h56j/KKPM5dYAsMqjdsbjF8z12HXciQHDaMQLb8HgMPwJsiNoy
fEG0hgRiB1rbEK8oO1okE8WqI8Hudei6DQtkj3tj+KpxNxUCe8EYrgckRdUoDSxN
YO/6CjdP/RPQUhu+PDcmBqDjCENqas1StkyfKNmvyvjhqS50rFuabN0uwe4X7oWs
M5UDI227m+4V6lYpcJnguVwh51u/avokdxkvwpr8q+/ntFya8ebxx6LMD7YDqBof
vqlQ5+PAEHr4OjAFdD86T/77Aga4WzFZ4g8YUcXTnK/o4QWD2EH7cMjXdWjUw/0w
4iXgSK4eOGLzZcumcYsHP/9OgeOuSONWUgC91EAe8/ychGvsACv/tbqZdec2PBFY
ZXiyf0nJwe+z4tEnyldLLREPX3eW1VVBPc7XOV6AVUnGKSodLYSmndTYlGpPiSVO
eL08Z81zdntJ7+KkOirRDm+pUg7L9JtVzRLf51Tx27GQN/eJSe3uXCd8kc6Z3Ft0
KeNvGgpvoUHHFC3x5QkQMlneU0er/mbNo+ILk7fXlFvkwbIqWFqjS/ZEJEqu1Vs+
5qBTfxCrzzeMw6OVRHbCL33W32k8ipzalKzQVvRMupj/oqIbm5YM7++tsgpja6wY
vVT6cXV6fd6mwf9X8404hGMak3/JsBxaXa6iomEYGVIwLldnSU5y0kWJ3Yd0IZGL
KN8GCwntxXerYe0fNe0M5Cm6HfXKTZ7TszEHiMBEohwhlZF3g/dRJ4lcxqqvykZv
0HaREBGGaPzH/sblZNYwj+vwo0CCUUGnW57GycVbMVKnLyUmYNjpDZFLdlYComPq
cop8NOgIczb72QzvWDvRerxXcOVKgaOlWhbQTmrZ8ER5BlDZOQ1ru+pQP8CJh7Um
PmKGTJMbhCwPMVt1nzJlyQt6+O2aO5py2KvfQeEvQ/EkxgaFu4rIfnCrj8jNMs32
6pXyooW2h8DsBTbV7Zex1gtEZyq+hNXULWzEIVVcWGW9v3em1zGomW/LD4eirdpc
n1VZ0EfLJLB6iSA8RHUAcVvatV58HataHIOPXx1ASWPKGlNJunNedVbE2d2yEtwf
rzVjXzhn64l0e8SiiFwWjXKmY4aGGGFy3d8DHNaWOlU/uxsZnOQp+pHzC59XKJFt
v1B0mA0WUzFDD6iNcvikStNgmuIgWxbb4mLTnMMiHKgA/ol5AKpbHUDG0mhIEaYC
SUaaW14EWuSFz3/Y5KJUBpZrBWzGMMv7liOM4yXNXFTsZNeiCxwaZkh/JgTCkU+s
Z78T4GY9rmGUeVeRf6zFJekoyBALmueNxK2aIWUws4MlZvsnDC0hQVugkHAyXgxR
LO0lawfVOanLZHOz6+Q9FoFRGV/+ROBrvh1NMOmMto7KON2I/Qsbs7HIQ2BEo8t+
hHW1Fk8B4ciIX6hA1wSmITyUsDlJPjKWN9U3WDpEJzRZdG/Oyv4YnkpKZlGiIMET
gFCB6QALJnKQZluHQ43bFpYQauFZ+32KfonP6xOvBTEmDFWDMxgjB4oAUpwFIN8l
Q6YXgDM2CqAL1PV8zOyVww3ch79NShvITz0eLntKmBS1Th5U44CMOTbl/fFPzrFA
45WTnUUYRhG6gfNmiDzreGo2DAnbl5XZZH1DSrs5D8VoUBbQKXUyJpNatfu6VATq
HAk2RTBpVTC0AK1er33zfzYBPSKEnbtd5MlbQn9VUjmfRvFlQnEl9lUV0MfVUag4
DVKU2KA4pZN0KzOMJbmOaeLTlhliXfK5DHRhij7Ds0lw7+z8qYFmq3lOSrBNZT+g
vIDMiOk1UgLfNfzpwCIqWxLbT1o7dgwfHmMdyDKVswTAzxsR6j09j331Qkg3CGy8
fhhv0srB2VU1oZF8D6q7/yilEizYrvrjZPlN+S5PozMI9hW00F/iGCYQhNpVB06Y
ZSapGTljOKC5VEUMLbkbJrGZfd4M0kPHjVU2b/H6n/LixQCa6JzGyCNxq1zMbbKI
kEeVG0qzYqxzRs2Cy03xF/0kYBdb342PRHXufie/F+YbrLStiz+i3GpUIVRd4b0z
mMQoFjTVCWQTX9B367K3n+pYCyiZNx8RDa20qN0BCQ7qK/DPZcZQMfctmnOP34/2
Xsbsypi37NCIu1sknLxijZe4pW5IC9OT6CDe1ZqTfL+aSXocK/c8HtfGOYwfRXCR
o3eCQpoky7tm5avunyia0lN2uLBGlfHVLmrzn1ZqWWO2PpP9ZOR7jNTX/SPlpQ/1
7VwrlOXp3jpgbyqZhVwa88P7Hzn4JhqUmiMElrzvSQXAHPtKjzYlyTrbeF7IbVt1
ni3K5ddI16a8F0rSJHlhOaSBMCZPiUwQZuhlt7vjZhzMIsREYy7WeMJOm7vGbo46
cPaZu9qo6ak+t9o6PiM/7F1grtSp/uqSLPjUks/HNwb90itz+viNpoDatmRa5NsP
il5rRAhtIPQtpIFcxyT0XuqTS0cRko1AYYq4uYs9fpVrhWbGIoCxeXxsgd3eDWvh
1BANOwaKmF0q9PI06I+S8QF+7IevSDZTcvF5HI1SjSmXAh0fxx/SAPEp0AnznMOP
ZjgVJbSHnJ0o+k2soaJPdh8OvOoSoECEW1xv7rEhtjJPoiHc8//S/V9CD1OMrzJl
OZXQ2q2ZE3FZgAZ47tkxtv/litHN8inhcSbRqA9k8P6ldr56mDfH4qDy31Sf3dnt
AbBPB/8gnG5aq9Myck+C2vgRONVuFIL91ieRHo7nkhKkmFBM+2pSiva3rzIIkX6o
MhWGGjxub2/Z77lfvNGfGuG9up/XpzIb6YMxyi32KEkm75B+xopn9yn/Cjg40a3d
eunxSxKuz9DmtrpfHkj9wH3fpqeDsIA4TAphEbeZOW0Jdiomgyg2vRozg+/uhtCl
Zs0dsSWmay9vfOcWyOnzUfZwEpL0ZkjupE9vthagVQ3h6vAL1/hwdy/w4N3ntc+S
xAy+toyIDzHVVAYPnb4Hl4zg/UXNUWHjRef1BcXblYiCSBmvqE8E7L1HBmwbNpOM
Lr3Aw1NhgyGjMvnK4+ApP6ZSB7CvruLUuvul0tcJx3ghv97IcAJPrKkt+Z2TtxaY
gy6TsjvRsEvGgBDaX1JxLk08e4B/PiCeQjrvCfbvGYnHLFCyPqwKXdVL3CJD60Dr
HSjfHj5lEaAHYAZRHV6FBdo6l0SAy7otxgrPoLTOHPLmIe/XiuZGliSMXniunv4S
NxgxLm2FjsZDGrixV2jLiXObNkTVJVEs2XpQKr3RxViod+JAJibDaVFizKaQtqJj
SwrOEhslRvqA+8dX4AwSC4B2dqGLlOXtrRH5JXiQHyyOli8vVDOLuU+HtGepmdnE
18e+PtDUaLlSluQHeqU7kKf8a587zKhEHye7kUEJcyhtLGATJVVc6ZX8YHIxVi0u
S4nnPkFJbXIBeh87eebHPHpKUa8SvFNI6kv4gN50qIS4J+Lvwui1aFlo5AQnCJvb
Oh1KgovTJCl4gkZxb1PQlE56jySZlimEtjgRpDqPgJEPEfIixGIbsNjVpIjd6GwX
rdwckdnuCOigIB7MgO0W+m2zxi8+GYGjWNiH6iDqrhaox2dbudxSraqy+Ds6dOxp
0Eq6h7IrmCDFiosksaWh6CMGNoX9HP6M+7e7ltGaw4CTW2uVpacQPp+VRwpTexTL
hNXQelmsZpOgofHWNBhVauSM7/EqRi4NV9CuSST4usBvAiTuBasnVNoZuJKQWtf/
r8RLqrLCaY/CCvTLtwU1jKoFzBz5PG4pgb0h7F2smhzSDa7jse0LGXAJKmu5Xwtx
H1AAokFqdUJHovyP2kQlrnpGiXipmT+nBs6QMJRCw/o2LGpC3c1wwcoRZTPFAb+q
fOBxfSmp6J6c7KNwMncqzvCkMfPPW0NwKc8jIlkVSCs8nC4Q2IhCaySrgS/hbSCn
YYv+sKUL5M5S3VWkT3S78KXY2S5KFcR+EIC92kPuz3o+1Cp9uAwhjMCPwk5xPTO5
IiNXdzzTNERfocB7ACbvSuCpbc5k0WCP6PlHCKelG97dy29U2i8RaaeNfBeoRugA
jvgHVJMCivC1se+9nCwiRoS6BnFqlZkRTdWPLez8XKSAgr0ftZ+h7/L5GQ+P/u5V
BTbh92TcxKRaI7Kxfca4kQ1itawjK46tvFtjgQMMktSbCmH2fp495OGun18Bm3z3
ZZ8gWYbes3D0ei8cxpJbE+1+yQUxzBVblz5cbsOtn3RdJpSOmdCFW+ffjMmUBZIg
3O21KJ+mlFdYPxzl/+YsAjKFjw2ZjtyOiYqDIu1FIdAkOo6lo7WfSZqewMe8d/S3
7Qi7YhpqAknHifIcnKtPi5wctWM4+q0OMEYdE1hDICmi27wxmK6vnMwg/Nx2W8xC
8nRs0e2gmHaVIFfwT8+HnQXHQIqPdr2TZ6as3w7i0S3eFluiCVDORyEqOhhMgVax
J1Igdokq97BKbwTq7mY9hKIjeJioSygwjwF4HfoQ217xmT3xk7GWFn3R0R7hNbRV
8D4XOM0JCikhmHS16DOE7sllj3MjjctQvIdds73zQllGvZgcy9oqit2Dh0b/XnhG
+CyAAKGMnnU6mmNz3ki5MSLgCda3bMqfIbCoM1/z72fx10yULn1WhkMSqIonG/rm
V7/Xfk0WIHb6oyVqkdOAF4u65Vs2eVqbyU+rbJMkjbXyxx1f3a/+gZEqceCG+52E
W+E0FXCJBRjffcmRap0P4bVsuGGcdSvFuVU/S8Ot63mDqguFa0l4YUASsO7u2ZAw
k9wbh+30ks6jtief3pAZ30l/vPY7RyU2JOw3qEBnBBSWnozJtCibNzilYjmNmBAW
47hPq3mnKngQYSYA37ygB9x4Hh5LPeBaZCKIGuYXAWNGF0wWBW4Lwj4LTB1f0WuI
olbYJEjLVNyKx2L0gvuaVzDZvOJWruO25sQhkzsApZL+t5Jk2+x2XKBEpPic2WpP
KcknsSZeNUREG3D+z7UQ09DBRlu+ri7NqQySMhE5MNK7Y1h31e4vtwCGAiiP59eV
KMtVo/+u02UdU7o3VKM6csXloIOtquE4BYOor5xpBSM6qWBLinecFUGfQk6hqix9
ftetiQDmDQVaqTMcknG09rcnbFrWBNoYxsj5U+AtPtNvmlNLrAIuxdsgT93GPSjv
hmnjq3z6oNTOLX8/jaBxCpyStrhuISy5nZm/crYXK/TtW6UV1sXdhXivaNzJ4Mzd
BepnIonhsK4nRAP7S09mPLQeQl2R3nvMVzZvthPWmZ3ENesSyIeqRAblJwtGSY+S
5GGbo+ieYPklDRKGEaeKu7fVwsOEtyZapKto/OOJIU42lyJbCDrA8y+IZgkfOrTJ
xcJlN5AodcFR1P2IDWVV97UjmyEj2fz+Wj8+qULfNR39bsIjdcrzEb+HipYsF6OL
n5M0u/4dxDe/FP0Qhjuli0WDeFadEXfPeabKxr+vFjjJa9tn8uAEpQHNT1iiGlIF
FpN2xFcq1ClzaBT6uV/tuc6k0xI4kSCXgC0WBC/itzzretn0qce0uHRxiFgJfgC5
dBtdFf35Mq1ZHv+byD8zPxe6FPiEfAIpNXeQKMTcILbivW51V8nJ4atB7uErDQy7
Mgxan+XCLiqx+5eI1nPSr+RFnRb8wK5ncfpJJtjOBuimOshVIni+s6xoQCVRLqEV
ixUK9XQU3i8W7QGByE3Wdv4iqgwTnVoyzdYe55xFgGR/zaTtfx9G0Wl63UNc8mmJ
MkF6bxx8LBMsD7JHP9qhc06NgnsuF2Yh4dt5YqvSzPKosL1Ewmw84M1PqIkyvF+q
6rqshn4Ek/dTJlDp8yVSEs4BWTyDI35OlfGBldIMpNyjN3L1rlPOpBN0SayAkBPI
FEFiZ/xz07Mrk2X3A8ykdc0+60qjtE1EJZ9arMjCgefLLnb3Y03rxi7pY84Q/Ax2
Nm6JHL2g+vsEjmQuI1Ivs9IecuhppaWkY5/cgD+bdYj1V+II/MxoPbA1b6T+X9rQ
on2x4LUH9oOGXP80bwQKHzLWIPqFccGh807zZtHQjJnrx000FJXtvUdLdJ3kItBa
Lsl2o+oKjtUzPb9wqaFdhoFKD/VzweeeMA3gmmF8w9GJkSvuRA2RO3NwwxE9l5NS
uRukmNtOKO592Yl5DxKSG11f9UjbKgIsBGOhJv9zDmmJ9ZOsEIgMEa8HHh7m0ml7
ga0rgwv0w30VuqXa5Sn8tRwVvuyxCeH5YjJyfVcHj6N5R91LD1nx8+L2qQ/qfBh7
xsXdu1GTm3ZB2KOE/7PZrC/6mSMRGm+RhPxKQ0QryVXaemNyDacCJsn7iqOMfVFP
ppYlf2Yh/7UFlAmZOoISZF7redkU2BM2F+uBTySdWPSCCjxTnVz1Cy+4qu8lLYcO
L7f3ZAUt2Ammsq5tT9noDBpqw3Xq60aLgrFtu9vI5F5bvn1ZlYIL03aqEye2xvba
6DYsluB7JiixLZkdEeKCnC4ep7UoOWIn9UD6FQmB2q7rej3YpaxpAL3hslbQYvHQ
B84ZfEKjEBmEhUwiGTFLeXcq87njwhCsyBQOVYoAbf46bRVxfnSROwFlGGjn7trO
Ezu7lNUjkrlwj38z3mY5ifwNJtg/ZQrGiWhzeP85hsk2kzl4+Kw1o7SGGME0b72x
oDjWH3m6V2ssZQrWXGoZDVybscbdq1DDQXyJKhPBtHl0byalPIZEBznHeJeqWerO
yzncGDh8PLA30Wl9MrwgLCILV73N2oHR7Qm6s2OEpobw92LNfttNXzT2LRwruWl9
0SLPOZCzxIwxaxjC5g3fJnB3D0uOQm3x+IC2HlCt3pHldbNiy9h2yPeXCs9MdIIt
l2IXx+0r5pN2De1x8GRNtBeM27NN8rooKLLQT0o+5QtROIIXYaAwFBzXE2/tV6iO
mqkROkVJkJrh5EKodijfT47A316IbMeeVeQcZ6k8g4M9li1welMntLxbs9ywzsvb
AnQwe9oGIoAOH8KyhUCDMPqIwj2MamT1LRY+tQVFisxCwsBf2veBQOBD0imWXIud
4Ewj9s3mbocAjRuVatEZbgZAPjbUgQs5P3MVwwl6zufN0cBf+X1iYkHvgFxfAQGW
MUmlf4Jm38TBT1eRI9up+yJNAAeDGwVL5P2z7s5nN5PV5+Zejz7JvoTE6qwnWvVf
l2A0EYEKL/PpkgI4XrveYzHptpgei9vRxcCAvhhCuxXZlxBQu5vig0UmKfaJOUVE
pprdWCfhM7zSXp50wJIZTKkhmrKSoEVHdbai6csAw5hiPT38zNwAED7CzqDCN9Uv
5DIuwHuZ6IpfrXeooMhPTcmV5Xsow4liwNFx9ho/XHjNjL59a5fJpt+pfaj0KrMP
brv1m/OVSVEcrzQxIhgT30bdHgrIIGu1rbD3bKS4ygt1fIrLfnnBWLDRQV9js77F
Qwtcq5UL2coQgE3lRhL38/hi09gznYPELgsWibpqJs3A8SHujpRXIB7hYtJCKi7u
wK9zwQaSNw9+O0l+kYkD6QIID4lrdC4e0fpDicgdW40xJY/225hefrS5Om6Zhi+k
l1LCFUhvjlMmM3JzPSbN6pGyekJAXjQ/gz+y9GkPVyi6IgpV6g3JveDKyokC5SA1
CcPtk7NRuooKqEGL0w9ZM/xaHQEw/AUynyhLT9Ztoh01vCUMDaxIzI9BRWteMzeO
zOx0WC7sW4qoI7HUyPcfGHAcaB0xg2K6CZQj7TVyCY433Oszlw1rKmBUzVYRi2ip
FiQLCYirbZkoO4gcWqCU4GUd2zVXqOVrmcERfxF0OKGtVl1Tfs4rIySxfq/W2HnA
vl3IJE2a3BUfBqMydQ6W8uLbOwg/HjX3RWlyss7YCQLoqVyZre6t1cKrZi04HBdb
yevSdCi+ezcC71jpzFgxv3PehCNN3UE7sZ43Br6Xv0Cz/PowRWGZtPhT24gjmMFI
2jZMUpH2WyitUl0Bno93sXpErUH4pHoerNMrr46iU0f3Pij6A8uDT7Uhwj0MHBto
TI20yoP5XqAcM1+CSDaye5pIpFN3mw6qh2B9aKf5JVWwiZDGnPD3xIpsaEsdsr8e
ZJS2e2DZUjrvOSQiPErQlBb66dOSRwQ/CX51akm+3BJbprg95TOpQonSaeH4cN8l
qru1RMyUoIVgsO/ChVxmuw6Yam4pQWZZcKujBRxJVrvO3ZgFTsHDhg1v2lEOM9LN
wtTi+ft+UKo6Bn7ZO0+aZaafvJP1h3GOZxhAtwrf1PMc8A45ClCqS5U0nRuTPNEY
sjYv/rQPL9ya86FgQPiEYrXQdSmRIRbdwV6STTENW+XdkXjs478RW4lWttJvXxfK
2/factG1eb3v740FUXJRNeASEH8cnGks7cH9AzbCE66gox0lJqUkLgNi6DY4c1X2
LFK9g0RMRGL7H0xe+AhIFf0wSspYVuxy+njwESPU6YP/PcE96JXb6YzxN8Td1cHM
dp6aQ5eyJ9mIsRFzu0csR4U61bOaZQcke/qLFbEM+QDa/k1BPrkSyXbmTY0VAjvh
mQip4dRkPJWL1ecgFunjjmGV4LV+HpqMaWjHLCNjtlUFtrllkloBmcy/29fMkWv5
wGpzJkuX4UyJQamYoubKXKmB2A0PKqivZw++e4QjgJ/CQbtfC4CzhQx35Q9t8A5u
gT1d0vfDU64ojOSqArLAxrbEildZMyAPMisdsSJO8Rv+y9Qvn/7zMaPIN1zoO6HT
OeDgCQsqLR+8PWB4XxrkZQD/lLOpgkZRFWirtRbjI0DEqk+I8BrZ4kkroRctobuD
ESSlhUyY6Q1j7zNGzfOr/Gk5Tiwt8Uk8ciKt/2rb1xBXD1Wz4IKoaV+5rpqo/PbC
xHuWNK7s/pnLefBu/tZOODc+MMZpXFr+earKV1Rmk2JzxKCQVeo5fs+rnZ1F6al4
DqvDlstKStfsOalPNimmUpYixhCC3LQSmWrAj2DLki7xBwHO8ktXheJZaFopFCft
1fyMhmOdLHJUNG8zA8IKz578PiiG8vAQpXljZr0BtndOxJMFyuTgn8E/+Dru5dL+
B7nblDc6rq+qeM8d8Cj7aWOKrav8xwokrRtupADl5xPkEDXyBiBMrxYOWylTb2tk
G8Wxc5XXfX8fLrNP4Z9vnGsOd8Z/V8ggiJ3ephCjB97M+mexVOqbdQqGHSbEENp5
FL6TvbIZHI7u8Kn2tsCxyljM+oR0rwfSgKw/zfzvJ6y6mTsdCQeFSBqmLtbcHuwD
vRWu4Yd1e2s6WTZ7WibyXgd0qOGozinPE9QyE0Z/eKBovIStxhWwy6gUUWCQu8PR
nZIlXkR7CcLUMHbfzYRs+b1FgLmmMsWXxzw9EdXIkLjd4EuWO/f768Bir/xGD6h9
bOu3neLfFcS+7vDMyscvDYO/cAwnOgXfiWxVf7H59urIFBtXS3Y1VIuz47NNDeR7
SIPrAsGT+fkmc4kksIPiLRUwIqN8vvzkA4hDXRwPpkD8UftmD6R8GCjU4dZXqmt1
tbGEqcNSzYyTA89ou5H2HG0C3WMCZfE33f+7zcucqb1ZxJo+xcDk7MExAGOljJyr
hiMe7/XjIvEq6qT9CJ9GSEeXsE4IcrpW3eczq3z9P4vfjASTlxQKHJp/KXmAzoiY
16bZpFHvfbpKkMjQAkWDop836njGPgvCClsZdI+hVFy++iyn/TcC6xEP3xPmThp7
jHFtt10w0ZGGfUmw3iuDFCaI/ScBns+dIfBTkWy4GFzbqnIBN5BxPyg/lttBoU51
Mz+psrfLZhbeK7wuhaQZwTupxEM7X8on21gbdnh+tzOCgSuaNx/vz9K4IcFL8cMr
MHiP1cHocwj8K1obmlo20dDBI9Z/DfOX5C6cH7bTwBVal6bVSDIEe3AmEzidZl7b
DyDk6hIqar1tmGOZWmu+t41yKei8QBtmWCIXC1GNrnvgMZSgedKMZNkE+b93EYxN
5O8rUMMaVRUu4Nwt86pkqAefuwcayawEHS60xZDpYYykX01ZgdEHTI4IL52LgSxl
FPB9/VsYvZPIAOvRoiyVeD5PHehBkZOjMCGcgyVf7wx+lSuw9Xaj4K+D4+NAumM4
K1sKM1l2TrTEE5RZ/osman5zJhWpeONZTfHoSa0DfU1ZGRszciLqp0rjhu6/usLb
6B63v59mkXku+MJVOdMytEY3nb2vrP/s8tHNUw8e6ip1ry9IxYbZUIgp92QrAP5o
ZfDLe3P0NXlznHbHFybOuI9fECU4EDIbAlf829eVj4sYxHz1oiqNY5uYZqxHzt29
1/pJLGUBLxDkXdRjIaybYQ0hhEOYyhbkVIDuDHh7RXeutCfAXbeVX3HEUloW+RL8
BpEJYkHSGjftmgnM0U6nvSLtrybnpp6KIJbNUv9rkb+y4lm5kqLqmnYga8mDFNfi
ah1FfqQFCTH2mndSXNRNDHGlp07R6La2ta5FJPupxFrbwS6IgOb0VQergjxxZf/g
u/0eUrP5++xcrnugpEcTJVS9k1uFyD6BhHMvcbn5kJ4z4NSfE+4LasSsyGGFTuBH
Bdj052I1YQAH7+4agDLTwMagee/QfnzBVGcW41P9SNhezPtdI2/V0v2ZMxq7aEqn
A4PlS5Ut4jZzNXcGLWWD6EKi+X+h8SS7i3FNGOXN74AZlp8cyJL7SV8I25LDN9nT
83o2mJT31bS2e/ohlu5D7+OR3CUoTmTZOTaGYmx3zQVksKllrcZKeMgICaITorMq
Dm63pfsMEl+By58uKxHemFSlj2P1gYxE8f2FIkrzic3rLn0e+sKSwzXKFgUzMTaR
jIQVDLroT9VmpiWWDFSQvir4mXL0ppE0nfL7XpyNMGpfeXXgSK/JCGWY0jdvDEOH
xzXr1HQORQftXN1MghIiY7UFkrFhNvlhckajDYt6qDkKf7d9o/Lcg7i8Nikg6ESr
B7AH9GFcfUbjlw2e1OsDLMRZ079VXGVjFrJCXAGLBrZz8tffis2iPAOJlkNG1LYj
kB/sFTfmExeD6IxFSyP5C7D1VWY7XRf3BXD3Zh+p0kZ3Ttl9YAqEnBjpE7qaA6Ef
k94fXSs9gzlUO7nxDC5LhmH+DkTLRd9w4eY8to+rL+RgFttzMtj/xKzIpNduYSuB
KNDyViVxxZ7WYGmScutSVsDoHHECuHo2zd34eo18xN0ENZTJEknB+oa9JbWEVdWx
VNF6w9va8NZJ/lW5NOlDMJi+18PsdIM3Wo9q+MAWlhWDvMg82zkTrUkr1XEJziTX
CkrV6Oto50xazGy+AnYdvzFnji3wuUBjj/01bXKN0r4wRDMiJoKK7aI5D5fUd4zE
KevAWBV/M0B3tTVd1xUj/wG0VXkzGbMnmMfi8xBun1fnKK2X/kHgOWN/2u7LBMNB
pLKVlin49TxbgxCNsgloVBrRpcMbEnMPHHPxHnFD6HW6bhlQdBAt79vY8hnHHztl
Mi8Xf3HBnXuNfZ4IBLOnvFZiWW6rdTjN1XldjW4AD2Chciu/jDPVAHCaVJ8GgZeo
E1thHr9Y5vxwZSaTg6In9HVUK8aA5s1/XpkZkM8Ehtmyu0HOku1M8ZSkvYIrqft1
KK2O8l7pWAMh/nvP1QV4OHc+3yOEgQFOi7K0MbN3ZE+h6WvnvfiID2unc986KYoV
ErQwmqgkdqbepoGkrMiQbuPIEVH8NzbselQCu8PCBznfWdFGIa8UOTDgMhtW1H2K
IFMXv53OU7bqZSJk5czpVae6q3Es8klJn9Y2/111Wz6cFxcwdewPzeQh8MtO7TIb
HgahkF8aEgeAiZ/l2qwSlesSVlXaLQmfh8klv8WWVrrDWL61JSzFxUjawLMOwcjM
wORXqLt4zQv+UwuDvJuyPTBbv38FiZjBIcj/K/yhitbESDmVpdN9mzkVjgUEYWyq
Q9tvjk2y70hqMjmk0Lle1YFQGM7iyutZ1c59KINRVGe2x9GwBPCSmdnHmJ6aibHk
i1Kat9Vw8KuxbMMLRmQfI0V7T8lroD8GPudyydNLFajZ/JVOxLNW8DClUNtpCaRL
0iMeRh1YRPhxVyf1WWBYBcQX+7O1KnV/lY8LEP1sAPL6W5+y0G6BGkbo2gs0D2t3
bdIkMzLBdotQKLl+vQ6qpJ6c67NwgnWKN5/3q9L5Ov3WxCfZe1gv+Hh+Lw/CKP0n
AxpujgRgfGcnNjR/pWz2SOTVTyW32+uMcKhGvIdb/wdIWDfsVZJO+qSwqCSwVcZU
i3/wHQnb+OMSNmXtsFxuQUn51OVIq65kRc6f+R90ozA7rNWbYs3Yw4AZU04/xEKR
5CIpxUafe8aGPHipK3Rpaz3kpV+/BkOZ6PgpUGeU6v9UG11YUPzVT1+32bxuqMcY
Lx0nRZz61ZTtfjbnmn5Vg11HCP2iBi1zbHNsZDHF4lD0PWB3u5+jz+f+lHgoFQYi
bTn0l+JxZbvUo0EryZmogWF+CAHAe1uOmtk5w8sJjVBBNcTJOpql/G3pg/MSRz9P
uC889C0Basy1As9x1yfbglVMN9WZUxJSii0w9hVxeQSa6KAjo/RON5ADlQNKfDjj
bmRnJJbIEte0oabNi7vfE2bEk6nhDqttsqO4cvD4mGnU6SBpwdAjjhKtTnt5iL9/
TrDrrmCInJJ4iT//8BfyxggPFHywYA8fQd5g37qkdhJ7O59PdoPwNtm362ZuxhWY
mJBrI8OWiTiltyQnoY1+TrUzicIraFzuSA8ddYWLC9srm6pWn6KRhw5FUC9yyO+k
i8kURmRjezzKiYLQlHTSkFkd5uBrIlZkn99R2nVwjpw6csaL/YYmHjmgYR3fwGv/
hsmcyEcs5P49ilKBmd099TxFEaiHgqwFLEtUCkYodIiszhHCdIzHk3Kf0ofizbs4
rj5xcmafP9KVs/Ze+SP+Gwd8ZhvxtFTAC6vgEx7b6DDvpsscbQac0rS322KCTnwf
hAQvch3EBB7t/5a/8HRS/5wDX4G6qWRnkPvUXP5QF/hF1F6Xul6t2dLEU5bfoJSq
rmpOQ7Mov1f6izpb9qwuZV1xEQYll2HWVTifpIz6EDWm4YTyEPMI77ZBBjSyPRbn
4/Ml2MULX8o0OxBDRHJ3CzS/gzCpVtBSSas7Ke74PEyLzBdngwWGZBu6joDwThFn
R7zy2ueCIvpaXcZXhlQuiw+/d2WqSVmj9vhkIXN+DVWjx9DmzDs01WIQG4G/4oeI
V0sv2llzibZqaIPWsxEGfpIsHkTJ0DvIA8Wv5lTkNO/XBwh7Tx8CseFR3GCKjkxI
hA7iwdaHFI8lefEMURUzsI9CIJJkTqq0EezxJFF/MfTKckM2d/TRUpAgTv7ocBr5
KL9EdLuUhk0q+WBFK9D+pMs3UXsbjr6eDmwt2UOALOnYPZ1E++EKw40un20IQVYm
j2jSw60vgvyJUZsGYx6bjXz7pc/sXvL1LSvpcUwKtJIbnll3ITwZG8D3I2PBY9eG
v5TtDtztPU9ocrwa/V6NlOWnCJD2Z02G9xGEDJwl8nu1CERgUhaGeM5uvAcmcor9
7ZOMLcKwIHNdaRBthGLnMIyKnjLtUfLuSEE7icI/OgThuQ9ek9HT3F3MhSvY8+PR
CN8gGKC9V2wNLZFlbujwTsFjfiEX+3PwuHWkJ6naY27FnGjk5BIToZN9u7agBqwy
xN560doq2/rql8u0y7+4O3sMvQlZJEE8g08AOe+sxDZqGngAheK5Z+BOBg9cl4R4
5dnCoaFFSwnHrjM/im6QOTmAV+ROAbx1FbfHPhm6Gcekqg5JN7rFxI+U6xc5J1gr
76zu7tPi2qKZEc9DKbi3V0aDLWqeeLzbWOptp7g2UIR7+Po6gmNkCEQNc+KDjzFt
0/VZunfkON9Rk0ldpznEgE2c1QOOvcWzcFVyudHo6Rd+MkSCzIhe7bbateJwnWTL
NQChcwGZLwZQ9sUwTFIIluIQzLh3mYsgp+hMaYjDVRXOaz8rRMpG3wHqqXQ+0ROk
Sg3MRJ4iO0P3J3mhwM+89hdzmsSYNjXTS/05GNLdCKE6ZPzdYBcHIpVbhC8Yvwh0
taJND59DBxaabAd+yj7lUSUZWP+B4kjaxwm5y5+oPSMctTkTScLXBW/dwIquzEDv
XC0YWy0tNq7ygAOLDkTsoenGzpqX7pUjaejKfK/iLEsU4x85fnZMHO5skCjPvUg/
N2tllm6ilfdUM6q3tbkHB84CO+heZN0uMRTArCigW+E+lGOC9Z1jE1VLaYr7ZnR8
5wRK6jvpdSl0uUtTytcZVaT+xUk7DwyBxRSoRbh3GjD5ApnEqwarHRplblQ9RIx9
IoHWL2Hg/p/MTKh/o0OxU5P/hQ1Htjdmc57z2Rq/904VhQHmbbj05kurOtKP1Yik
aFABunn/v6ZEYYV2nx1tXZ2eZpuhdeIfX3nrzqRSmRMU7eg/OIdy3vCYg7Aj4wqw
9QSTN7o/teib0JFntjrnVUWQ/grxnA+Ev8v7xK5YqFFQhw/1irmYN5NPCxSnuMHe
LeylCpe7rbAlK5QOPdFsuFDaXxgZZh+llvF3RdhJVX1hVyoz8IWDNKYpffczY08I
11clLNKZ2w6JFrbTBA8Kwpy70HurveldYYPVXcM9f/5ES8b9WkO0NYOjH+agKNfo
pid2zYA+3pWA0Mn/tT6m/EPg5Q80GpNpt5QTFHeZqW0LBddrNL5kqA5bO9eZkVUs
XBZ7/4mznkBvJ6aTYKHrYrzBUVLoxxUXPUh9brj2XA+n4fPwCs448FAw+ILCw0fe
vqZvpGmF6w+eqCU+dPj8lnDDollQffOlhm0WzaoX1nPZqmxj0Irq+fIpvSc4GQXj
AiZogNIDycSlsymjDlycwDs58wKZOXTPKZsbNFwd3iynmGLHxxgbGoka+ZQzQpfW
kQSARH81/gwcfcx8f9ubW4XsnzKj5lXlk9aPU9cpDAzqsLBUJvi0B/SGPqaYtBtE
ogsv3D12P0lgBXL943QJQ7CtsbPKmhtBlU2SMPwvz5izMcn9M1hztbyUhkQkP5lX
/mIKUCtjU/sCA0LLD5AMjZ2gaJhAx/gjmZgLF6HOo8jm/J9EoTEUjh+/j3uxPbYy
L1Bs+0xJH264A8GoW1ZuS7Je/p/mQ6i/5UaqFGvDmZ1+TBQbjbSI+MwR712qV4zY
q3bG/f+P6hPS5rboPbAKDpZXOhLRjZXuykXvp44PessdWxHpwA1KTn5FefpUzLor
hTA/pa0HkkqY0HJ04Cbk9ymWbdnVR7QtV1ndVXwJOpn56VkTZjtnlse0ksJL+Tye
BszyKuQiGBcFUrFLSIe811oUJ332Msxg1+t5ZYzGTWaiv6Sqko95ZlOEzxNGlLsP
EmfvWRyHM2uGxyPUtb1xCefAAiMcrp8+960qwu2Wuv9nhfr4y23X5Lib//JmgZqs
QguPPqAxRviCcEUchHB4vrDoUj1XENaAjdY8VKbkAKom3bpAJbAtyBluH5l66kfC
Rt2+cYGRZlBS/J75EX47r8zFzJCgCe66xvj0A0+6fFhdu10VSpZnGWxBZ5Rf1oPG
b9HbXDfBqmFXF2O7vfMDgRYRnjHyS/bvZNHb+0FGPIhh0bmKMSgdDWikL6Bzu1Gp
htQs3UPh+wsjbi1YBVVXLH9820XO/Y1wISVnD/F3IT9uvk7O+IfxgvKIG5KA5to3
SPn9XX0xflSXh70yH/zR6iaDkFetsREtwTaRXPwCNAn713t+f7lN2mQYHMzW3nwe
pjhaK2LbQdu45yQKBuyieo/V6g04P2/vW8K7LOiYi8ognoylWMtYndatrGg/D6kx
s1lepPNdhcIfFU96+2zrC5iOzJmAVg0rSXK+IN5XGCgRJEGVESHAPxTUIf+FZtJ6
RTYAJAbQ9q46PhK3w+9kcx9WYyIX2CO7fEAJuT6HCzSh/6yvNCCDmAdp9lG0t/lS
fUT9j95E6/XZ74LUeAIZSS//X3mdCV8hatsoTLkwTxv0wb8H7I80aHj3NNRlInhK
a7ktaf/hM2WcxuutvADQZ7t2TkP77ts0JEocAZkR3zy/5Fk9xCTkvkF7avPXUnYW
0nyuau1DsIWyHziUkQdZYbCO6i+s95gaLml2LsTZy0GYgWeC0AKbaDdc3PPzgvp1
5GG+AdPStrDoD4GnivxhMZDDQ6IOWNYc1JXz9VGdZwr+j5fWwvmBvLYSTVLkQXtA
ORYD3VopHbG5qo8sqpT/Ba8AXXGEKcp7BB4bHq1cw85MdcEUeBYxk2b1OO5CJ995
EFwFWvgd5SfqCajCVsX1b5mfZTCvEajpVqQq0KAQBdFYHNBSucx4hoXw2s5ZnDTj
NwSsRV6Fxhoo4pePy9WMSUYAB+LHowjWa6OBqRZHcNpe5nj4WyCVyToaIzzk7n0l
ck9VYmbYKgiAZo91L0C1pnii1Cdp28zEatLesqbIqOV0bSRWIIso3y0ZdStrxYgA
l7OR/ggGz/LAY4VTP+qg2sODqnWW8tct9yXqF9ZF/+FTkTR5BqBwRy4e6qUEzFWS
tZvHFkoqglCOebWwZYSll1eXGVYMJmNRjLpGmbH3ue/3OLscp/qJOYjpwSlE6T02
KXtfpLcobG7l7ckMiew+6KJBMQij3hTH75nvycs815reVjX/5qs9m+AEfMQuMv/R
Vk6dK4opb9zSN951wB+hsgPSN00OSik+lhm2bUZwANPqTefp0u1ctShiAgiu+qxZ
M8i0JFvsAvJq3a7fFjSjgo/8zM5OjuiRFT4Lw1nSgMlIoXr9lnNQx3Io8XdOjnpP
RpXYECRoio07MTf6xFB2NJmKkFMxU+CckbB4r647eEWgzqUMkWQa5OvHVaHLVNQo
QNEr/jNPpAfJcfMTUmjOSwxDHq2Zczjy+yhiFIAYkL2P9BVNVD4VqNalSSPCSmR9
ULxvhknX/EUkDu4QF0UVbmFQo60tQIPFu7GcU2t5ReDon7NkeQVisje7jIk0TowF
xQk4XHY8Dby45YIGzC0oGPXKQJ0Zb/8vnt/3gOsy15lnegkkApN/vPQ/7GpnqmuC
agpWj8yJoXDKQ7kr1M0/0Rp4orJ1wlOPVTDlaMxfgrurWkd0p9dZSDAE2LEziHoZ
BQ44FtJ/POpyAAi0s0xfMXEsRCsu8fzGZYRTUCORSBKv7UHh27MmDcC5gDL9JEfQ
ttYXCMfxV1lWZ6/aHv3PwQ9b1IP6le0P7pjMk09qp7TeYYw7Bur+LpOw5OaXVG/V
VYlFZeFYgeTpscYluSWK/pqIlvfnexajjqNblq9Wh44j0RnhtFStMCOA2XmEo45G
Qr3UzbhaB8+xOCmuQvb+R9S8mNTX69PtgTomrTIA9s3LJprtFtWgjt2wSGiyhJ9Q
iuGTP64ITL0zCVZrsi87DmRIF7fma6rLItXzQUhg39wqksTKyzN/jGU3oq51q4Fj
eHOUU8uIskfpXJmtIjOhbPP1zgmlbfK/MQwIPtE9pw+KGlcF8iYqK+TjaYUuN8+p
7WQwKZ8wk5TZkJyp3jtJt3XPnqHYE+61pn6FOjR5VSzHKSEYucvGZlpat+QVgBpp
NUYGAmU8IZHZhfH56WeXEDgUPFxGUYahyL6fYZGrJcApeUmFYmXSd/ij7Sjqu4Nk
IXTA9RzDS7VSY3uiVCPUwqG+KGX2m/Rfi8grKnIdhlusuB+VRhdkb9XQ4HtrZlI1
Up2QybSA5Te8zbze0HBIjM6irDcN+LVkKh+J+nd/7uZzhK0Ah3cABhwR4hJphqWO
5eoYHMRp/uq6aiDbBEXBu+j+hHJC08WYdVU2odmPBPRArLBQGHZX5EHuENGkEqcB
4n9SdnX+kFrpQLu+0/InVSfjYu9mr1ABfMtULv/nFMc7gCyYmBik7gT5FzlIa916
xCEABlnLF0mz5GvBWGocnFly1O7ae+4ST5qelEJGkjOhv0jpS40owMo9bopYYXHQ
YGPPDZ1kF+qmzHBd+lA/vWj5Qn9uOqgUz0jENSLsDB+X2AlH9YSEWSvZ+oY55sy7
k3Y43763scyb1WVN2xHGprafiQbP5OjZq9/FQh/hEiUgYc8pA1l+dGKtfqhbK15n
2uDbtyPNfwnL2Nb93dy08a/ti6jlCBWBErAwkx1CIwWHRPLr8pIOUTmW7F5O+O/J
CUkzg/9AWM/rb4t3Nr3jQcaO2wSy3zX/Tmj1FGpcxS33P5c6tFaJ1sbRrU+f7hYq
xPXyH1vC8qrahTu+Wf3OY3s2Mw1/L1Bs/8iEzI86/uQz8OgFuuWKj3gnDx8JWnz7
KJ1G/FBxq3xhXhZ/sQ1EVt2S34Eff0sr92AXxiZmmAxiW9PicNsxfSVzXBO1KI+H
9M5+ULGMq9EWV++p+4zYapjiSFNHtj//h61oCZqyzlo5a+kccjG5npn1hzIeEl2r
0QSSYcKc5UGPm/HizI9L2eqJm0gbHOg8Zua4xUkJdbYU3BdChPtU4uGKe6UnFpvv
B06Dt7sBCty9G5uIX7BK7LSqhTF/W3Kev/taBE/kQkW8UBj0cmAIQ28dnP/7KWBb
JMpJvlrXE8I1SVz+t/KS/bQfb9+hYI1eBXDAdDOgguF0mnFs1ZShAkIdcKNAGxM+
nnU0QsbeIsKpYfSu78tAIPHeolsDZpM6MalJSpuVv+PSL/oo+uNKI8H+ef8pEYcL
PWaEEduf/dCjNZxjRbm+OI50FG8iOLuR++bTqX4qoy/NEXCzLyS+gXGmVBwo3RjL
tDWCX04ffHVMWdpTvwYOBS2ZENMreN/3vJRBoGv9fQGckauDZsFiG5MckRqq24UV
7Wp0odh4XTnCHydD30068XKu3LCCCqssU+8YvNr5eNIiNigjbHg59UJdzZFdNfwQ
CP83rhiaUcMhWP4cPdEeg8d/ekPmURIKJ41qo43OIQ5IUTJYG69gVnraypmrAOg3
HmDaPL041xbbO4T9q+7lrFoPfuRTGgTvZo1zrv1EwEHx7ms1SYvtj+6BGr/wXQxu
zU4PXG068X861mHfh+2ANFtHUAe8m8lp600wo1YgUNwXWmO+B9OBEi2Q5Lr5gk4z
c83lOKCPdqDIQx0bfn7j91eztOjY3FsctKROeYuG4W3Eae2MYqdTcERmugBc4xST
6gPuVzqO2AFxWMKKQy9EiizYWSdTMvNf8X88NV0PQ0TH6XP2RlwqDyyE/bzrzn9P
jRTaNNk7+1s8LK6AaC/vJmj4ZL5U+KEvVYO4GNjqe33ixsHTA26V93vNB/fR67xS
m8ABo6KRtiIgz/pxKEzql9nLkRk/pU01Pg9rKTJqZpqMwSXVkkyyrkr/esAna/im
QiCB7bQn/qA01QZZvtKqmJl65XROHq0tjAOfDEgzZESbaYsIYG0dpvtScsM8SQUm
PGrsNjDV7RwM82ALpE1gqVVoCR1TiEQ1pOcKWnt0qyA8TL1QuEpqkFPbJeJYZq8a
unvFzJYp7cAI15iOjAzAGyl6cVBZFnaYMpR/jxNGNjWQofiE7z6TDiBznZVFpKYV
OAoyotugphrnmnGj7uoI65nkc4Qy4zEfNgJmDRRE/EHLk0yTwEZ/5uvkNYHhntlq
p27gNvak1PTmPjk5s2zRs6g12nD3rcN9W0Sbmk95bdNPyD3qe13BDMmfscBV3pv+
E1V4t32zKGZhaG9KID5gOdDVXf6jEeHB+XrzYKCSOwLSMjdjWHXS+KcdGCuIrLrX
ZQvHDFelmNTRF4aNzHc5EmufxP0UqWLEWVnOriSWILDBRD/KNr4LMSoevvELlC6i
zDIevVpDTar/ERNBQ7rhQipWGPFQrpJmmdyLxk+nSBirKOJkLnvrHL3gPhY7eDmy
19CnKlBNkwm84bHCkWESASbofP3EpSSeQg0L8GbODk/BjpH8XlWaFQ6d2+LTATd4
7JWZYQkbRTJ5Q4hFMk32L2s5teoFOGyVg7GunhifcPRhxV1YHqA3xEGTEMSeAnUM
nPX8IsaSs3gHwe02B7z/xbMfyAWYkGTXk+mp4ha0qxI9cs7CBUJEaU3H84QGj+n8
GmBZmrowrUYEM1PwvV31M+YnsEU301aPeOHVifN9nf/Vx3WKF3r8MO4D7qjuzhPF
qwtq+NwI325xaNVyDGrRzH7SlAXWrrbciExrxzuvzevkvrfeFGjVw88SWLSIURc0
BnbtKTUKSSTu1+ODRVGN+yKjpfopgNUcfEVsugv4E6Rdh5ABShLCjq+b+uSCoOIK
yB6W7zyq5239hKTxGc887qRpZQpd8VReUcJCGLL0f29BJZj/Raaikj5PfYPksAU/
hMhes2DpzojeuALcdnFhcovb1OAFKlA73earJFtW9UC6MWTjxIw5NMC317X5XNMu
sY23nkPT+pVlNYmhGLcDl/bT9yrN12vAakfctbzyOsxlCfdG2kVs7Ag1No24BvOJ
8VDPFO3XZEIGlYJg2zgecQ9gB8VSb4AVxWspssE4yHtDRRZTFT7YsnRSgruZIiYC
1qt4PhX18u98ne9bklVqwNa8teqUSh0Q+izhUzI+lfKCzrxP0IzTCvZHVqODqvZb
eixBqNejf7eL3E/+OXUcTHN3XxElugjl09e7CNZ1wBJWcBUI2U2Rdt6Fvd2+aPXk
DgNgsOSZFMNJ6V+r6NtgXh20mfW8XlS8Mz9twjktfDPQI/D7LGqDLkMg7tZ2xg65
l+2GeDx5UKkUVeg0LMl9PDAtgo0JhEuRpSEOymq5w/nHTDZL7wN9pt58oSCdxPqK
v9/dhf6gmV6SnCr3YdvPohGna7gCUHjdfnrvW4grm2/07rbPr8ifu0wY3m1302h6
mFFMMQfD6//ZGYHP5XX/YpJky5rD59gLXiGma/lWTkh0nYEg2POlY8nBt1mbs55D
YdPqur/XFXUhaCCLPh5nHXl5rmyhtZA9NvdEGJ5JaZ8/+X3hpIDFSXttIY1Ry8f7
ZfCbYKdKFcVztFOhRtdOMY+mgkAByJuF27DMIFPZxq4lGO8TqGQLkCLi5cz7RGD/
8tjPED3V8BrBQy59kLyKzYSJ020zSSXL0HlrYVzeoy6jq3U7hY3eMCvveNWnjCGr
xaw9wcc8jQxbiOkKmNLgyDcXrJtXNYnikGsweCvPUTIrR9uL6U0rNlX8ymh+XHjq
iq3GVuYoEOObBDEiK2qtcbgYUpuaC6l6Ygywn2HO8MUCxupnGU815rLLImPxzGyc
WXACVG1DrGatF6AwIsWUJSWlS3f+B1DjBgzBisggADhC6Qvcz2q3C+43Y4JpAMcc
e1Qj+zmCszG28tBj14T3CHeO+MG13iqLGhyVr01XxKHgigqyMS4oCieOBo2j9gQo
Hlq9lj0ve/fL9vgyLDlhdCSwws8ei8C9LPebO7BCLv5sJCq1IZJEPbmmBANTtnUm
Vb7DebNlCgWHLg+AuReud22yCBAFJDr9UivtqYeNbu8DelKAzssnNKQZUq7Jd7B/
G/yeUr8lBMZBIo3IT8OSCB+2j7jhITIBHeq55SBnofZJqjHQrt3ZYhkHwA9/hGs8
9X8dIJ9wTSntcqKgc/Iutct+QEusEEKckfLeOJJAwV5Dj62k89yPvidvpdtInnO8
D+m2EoeLQxdVz2k+EtGjbCXdrczw+GcBS6T+FjtNpU6xjC6sQJLDRenzI5W2JG5Y
8A55KbnOPYc8JnbREH+HIOsZp0Xv9zKXZ17983FyxBhQnT2tfdP8I7ogQgR7SKQX
3BMVEjI10AbFc9Pdt3D2XFfLpkbU8VPL37zO7LYSjunLVRmCKpCEYjaOVEuOpAEY
8ARM4rFmKq85025M+noOHEng7dgwjZPtQLK4HQYXEALhbsmGC4uJqGF1JBLcwmVZ
SWrqzSte/chIW9WMm8DWfdDSdO2wuGXtWGDL7JRCAUNsiHkt8Ga6MmXYMde/fwNO
mQ4AHC/c5JQPc5zM+e5PuwnK73cSTvw/ypkZBEuhVcuYfjsDu7jtT0lFJ+eyTHZa
Gg3ZSOba879ZpzAwDnx4GA58uiqgZgEl70yuTQEfUar+c/DerGZQs1/hkeGa63bY
ZxbT/+epjlUtZqO8FHAZnCMQg1A2iUj3gkxEc61p7RTbKQ0xKFUCPCQPQTC4eRmg
PGsDHtoyMZAjZtqu23A3sbhHxkrMcvw2PmUJEKPWzBluw4wXse5qV0q3DNdtH9zK
Pkta9qBVqOIADQsz+5NIStnHT2zdUjzZWzbzMAyBkohmLwyyMS+FL7kakBdps6Ny
zCEMYsu8b93EQvuUVMWfKe4kVE6vhiaqn8MljP3Djro8d+agegl9NcqSquRKI7Mo
H04xcoVAS+GwRgM8xGjS0rqreqVH22KnFeEp8mMR30SpP4FdMWrU/lBv+r4E87of
rMUtXXPNlHQQkTbJ9AspnGdJo87f3kd9QFXCvoDzJAbmQPWMO4n6t75B3/G2j8WR
6xe6zbJvwC/CoDGSTEBChrjbujN6fGEUnITVrrotWXyoQA4fHDmvN+ymn9j7CTvx
eBUyLkAOlw/PUy1WaK/9a5k4OwMVAiBG4xVKlll+mgMpJ4W//rnwKeq+J+VRZOWt
tKzQO0lyRelEJ4k8ns/dVoy5BjlgEGMZN+xuhrrORnct7fDTmXddhzfDXkj8uOam
lMG8SBuDNayqyadn/0L1OmwSfMmbMaxoxqEtTFB1fbbE12XwDaatUHd5Fzxa99FB
WINACgNZIrJovYmBJc1luRTp7AH8iNvXzeLlNZTM411VE/u23c3U2odxDdHo2Vwi
QoX50T6JvSFFIRwngzSJy8XBvsQpQ6DbiZY6MDpk3EDhx9gzsEkFuQ87glPuVZ+R
u+cUGrdQ32oHce0Z4pOjAUq/2rryHoKHLK6m4swf6O2DkS4zCn8DjGdPoy0sSKRe
Z6qHXIM574CqQq+RbcszV8NdErMALS8UA0sgdouVk9bwcNUSCOXdu5aAdRzaAFrc
v38XiFDzYtMSSE6wRSBDXS9ZgpxGSM5VyxTwRLayQkXOE8Dr3//Ue3fWZKvWGIi3
dp0Gu0tcI63S0aQHscXEjDVDNEg7S+v1EixCJVxFiJQcctjB+xsdGqQJibg9/Ioj
q9JPdiK+GolYQFzAB+5XEJEPj3qg0ysHk3jzxDOQEEfXiR/FAYZz+Vd65b03kMX5
FDvM3M9qtW/aothNivok7ovoRGkYBFis/DvYAiH/PEje+p6ruDMHte7lVq4SE1w3
ku1ZeJjVmYd4QhH1HhBIvy23PU9LloaTHTJtaLzZbznBSosH7XGsxslEH36SEFrz
tULCVhKpQOKHio47QGeW/8v2DnBG0lprE3HEdUkG4Pa2bJqW31H7pyRGTBkFozEV
sTHZ/RfGGR08PNr7V9Siey1H+Leo0wfn6T809VcQxu5pzzbQKArTn1272YiSiHN/
MIy5FDnMhSYXoiVWYJi8LPc6JE9mvc7yNW192R3FU5UzHWjGnPhhCNINCQS3SM0k
j7edh/XWvyuM9hYEAqGvpzyTTceN+9mrK5jKwRtskhnfqUjks/9YGLjtVWGV2V7V
Kt/Zmz8Cg+TREpxOYDaGNFA6lyc1OUt2nFpci+Sgae3848rQ8wgma9tDr5iJtxYY
wYwWoka+BNYaJwD4Te8l38dOE8/3HCss0BzZcA1QBOKTNFuFmNLbg+8evGtYrpPR
95jkHH8ry/gMKYVfXbEJZYEChUKzu88sMj6JkpUcHvlkaeilMkcPOSbz71HglnuB
I6rTsuX2IB2ey79SOxpLjBS+W90PM8a4l9buQoTLgLaej83DgTlKpg6tcnKW64/f
5HyMiunw54OVoReKkKXUaq0cjpYiM0dlZ5iuWMe72uyg1VHuxkwpNyHQ4tSYKzcD
wZb/iqUJn52+EiKahOvAm+2ximM3xYAXsKgxGCQHnRA1XaGDjzM6Qoc/Sx7GHV9y
Irtt1BiYRj4KplS/gkF83lDxi0hBekqVaQkKuyVRwwAkRCV/WwJQMC0Q1Xct6iUp
dBeVusgJjmcSX7J0X17aOlIIhY0b0mTlVauTm7ff643dA9Hnrn79TtBhZYm9mwKN
InsQcvE8WvcW9wa+yrC82bza2cBiQc/JVIn+1PmfpWJVJDImpjaYQYV6yNS5SKBO
qWO6ApfeBHgbMNrf8mJoj5TWJzeCOO/2AKI7tlAEI34UY/b6qA7jjqu2Y7YZVAO9
707vxvwX6gh1YL1/wqpKziXels4zN+PkzU2P6rRaaaGz466XSCDClg/cLZKN/CM4
qPNqBVFljIk8ZkDYii5BRpuZjssB6wcz42Ql6AKpMQ5vGMaOv8DyUWCyoaFpQ5vs
xusRM+mZUuJ9KUyV/zNrsPbjPpx63B3hZ/GIno0rDRVAeJ+XdLrayhgAJbIpfJrl
D5rRg05o4u0qM+fHY9YSz6pA1kx0V7fS6N7V8A9JJowwrnFWt/ZzW3Spdb4PejN7
8JwVziGKw7KoP+8+wQl4r2CuyDKLvZdnWWkMalJYhwL+eCtZ/8chvqheNTjvYZaW
x9A5AlXrbT1S6QELxEITuLH9AZc5fbx/9anptmtNi2xa87R00mhK7eXBQwfIySP0
7qBkIB5NynnlBYfJ2P9p2jdKF3dLME8vm2KSUNEtFH1JNLE2Ds+gASmACxw3+T1o
PstDKYecRhPLH2BhVL+UWM92AmgMO7sD94AoMHb3c9k1lEGOT2g6SmwS/oxJS4ws
iUOag7oBMDzpmZ1XvKYsbwhXHKNF0ClUPj9Y6YvASvxA7U0Va1YLiOKrzRDX5XAc
SQ9Nl/217AfigL2ypaJI5p9KsTPsqgpO6LC6tYMFNYh7903BItKNNCmbEY7VttkH
uLPVm1X0X+0mptXfbewwwG/HrDa95Rchsxr+V6dD5cT6XXDNwXSFi6nIC/WjwofW
opycwSJBrpMVPnSJgM1cqNIM9Dy1E7IGPYcXGcM3d3kVGDlkD1UBv8GXX8HzkoPm
UYvJQw27XNzD+CGcNsFj3DPpQEJY284Ls2A32vBpmkeizGgKd5LOCi3fOeLBuWwV
c0oQjE7zjLPLIz2q5+P69dHFF7PsngeVJAOX2mSkohwUkQHG6hVIeX8HkASUdHJc
dHb20kzI+nBFLUxfGi2tLGkx/sMAv8+dWNAnxyGdof/TcrM65wnyQJiD7HHZTkTg
l870ARFkNTHS8nXqRjd1EOQDQgEoEqAUgy58ulw7pRtp26nA25o4sKB0DTgc64UW
iP8GxsYF8C4LTR8HnC7O5p1Ij53lmaKy+Bky/686eMrGn/TxzGn0T7ouzLme44vA
CGTEiPtXF9S6RjSgeEkCWws9CtbOrkGyLmBvx7QfYLdDNasjJmPsRwYeKoIx7LGY
NC7NSqV0mxF+op8TXBNTbUMU+9nnsUKkDh2QrrJ8zglhbgFDwbBri41g0cXBg44b
MfK32Xf19JBZkzW95iLuXSaVqk+LbMDgW+rVLyEk3jtGpjFCZwTqtT+eu7lhqH2S
KtmSe6oSh4XIoTkmbtWMfFHc/k/XhGyOgQPYPMCJBh3QGsHPt2LWdYs18uMb8Pv1
t1W0MkAX6g3nSQKrUa1WKkdvTRA52OOV22m4/Z+451cRLeP4GR7lfsn22w3gYJ+h
av9kz+tpDbflfhKydDvWX4vSExAF1deT762zAwYYWqV6RjbE/z4/0iWwOXx+JMQt
6BIBBF1KWlriAvqkDFup7NaTlYPIgWbmToND84pMYZ9vg57pqmRkNGIMQctKDQdI
DUJNnDbtWILzGRhDL5Xnjh3lpccfrC3vBwthS9MbluTT+ch1NrFnABcUpSGM/ytc
erlXSqoWs4eQItmTj6uBN1c6DJ1VtbwYYWiKP0n8YKfuIYWb9iCDuXMevpeVKiBL
zc7IvF43chVqNXXjttsGzXQChHRq64eiSsE7dDwLTXG1tBZzhLBJ+H12EVtdzIAY
BDHXk+fJCQS4dGV7e5/Wm6dhjNspsSte+SbLv0EWPEBssbPeARxMso7RayXHnhzW
TvGLRlQtxrPQyRwFbDVh4cYz1gGd4z5MLOpN6L6Lh1i90L65S+EFuw/6DROyItbm
Za3Lt7YIRTncaA1CKWhNEseHoflDXWcVmb+S7QPlpy+rfToct5BgzLsSmcFhJF3x
lzenKtDPtiCcG3KP6bwZ7x/q/PslE6QnfBJnFK0sy/3xIzqHcjz5OCZYAP7cRvp4
fHYs3XyCO3iMiTWFUWt0E5doMJwjQTUl/d+jz07Z1lZcKHGpo4rV0Z6vBGUMLTJp
mdBiA+biFdOjolgSR6GxDq0bVvwy/qDSDqddqwISclYKN0lw39JSsg49Fgm6uGT3
uUPX4G4b44mHfCatfn3w+43obVgpuFBS8EpzWuBBcDtKnMZ0agI9eFXzu2ohrGCO
JkeV72/zCvyCzcPNKKoEZcGeVCL/afF26/vJmqxXP/YtWq0Ru3oUf2XSlYMvbMar
MTkBilZBIWuMUri/yrs/aeXaBcP9+k8BoDtlRLprLqvXDEHzY/gtb/nHI7Aqh7/D
X6/o4gbQmg1dXJGdvqg8hz9UgHlsBf4fc8iY4qFIbmqTtg/TH0LNxUu4pnjBzhug
g/ncI9Nbql39vdqPO23/H/SxbwojqbyP/NmSe1TRc/RiAv4dWakwHm68I/uarIqc
/FbbF+T0DxSVVNqDjE0/5KQV0FxD7i8muTA02um+FL38PxjLc3no8FSvQ0BKbjnh
9+4Nxz82KFVSdukCPjWGaYcv6ffXviEgfVSPRr6rDPi3AXBJ4M78sTjehcUb1/PG
vYyRRfCvxlD1dfDUijCnv8Pc0GE8V27Xibx3CeJ9I9ybNhy7xdsKYeYXspW+prq2
PCeCPC7nXkJF+InYs9qiAFUtUKEhp0bjDxv9g302ztZ+FhqkeSicI9vy6j5knZM3
bQeOMVRW1elGdXIfGzXcivOx2cBdJ0P7l0aX14xjIp7wxDWFRJSdzIn1Y+qN/qWr
ExqbGh0zEeQ6m3TCF/YPjbutpnZPurZIhCM/QzgY+ESgSOydQIfagtCrH7J6mx2B
HjaUPtdSTFgu7H3UwqbS5EMXuHu1VQWXXCY3VAVSZcp/7iYTbDbXZJfif+f13gbf
Il4RTG/SwxhWkuCNOynQAoP7EtMrfD12bZrHOobcmeExhKV9gxsaFk59FlxrLRSM
mDRBs4BeitWaWiyA9XToAsqZDE2ZQxcBtwS9rJ/ad0j+KBrk48YNTMhatJ2FVvKs
U+S0/3guSnWHg67iadSYoqfHEvF/nIgQqNyca/O6pEYADjNRXT+d3PHTGVCkdu7a
o5lMMnpDH6ROYATbghZi12k4vM+VO36eCMZXVVi/8dti7U2SPueL95xJKOeCd1Me
MMDP5FdgrCCrO4JWd7adUXbMueE0tWAO5/11qNxBQau5P4MwtJwUE34ljSv+4pCo
Q/eQTLZTvxnmEFNxnnI2VRXYOlIFLvT2btqH3+VdD/eZIcC41osR39kfHs01F9sJ
JgVjFpc0/D5lwnFXdl4+cqu7iEzOBp2FBrfBqBNXyYexR3BMuQTM2Yn6siEGZhn6
x/lVJm0ruBrKeUyW/kYRS1WB3JX5PAhb8jZPPL5WGP3O6fi5c9iVrzkzFCysQcd5
hmkhnAf7gkgog6HJjWX6CBkD9ccEnfd5ciWjirzPv1mGVxvvXE9paJ8FucmvpX4s
A5RwCynzLLNRNeKatMw4smbxdl+lKEZVPa0CL+PZIEy2f2lKY9dc/K9bdCQ0JGvf
2CdgRpxCfYMSOZZgaCVkWqyqeac2Vj9tbp7lATykjsOOLcsHW29Pz3chuli//pFl
f+hQSytJknXM7PEYsQN9MAISMz63a0qYMW7emZydVpNrXk98dqrZHlPj7N1L3bek
/PMn5QUQnFGWO3sfB0dR08P1+VMmNbmPSLPti1jZ+kdYHw1gjkppZxTDlaOM8sjT
8zSnBFTXzUQm/ogSUcj1q0zqM0uUnd4hkKOLTiEoATG1HkvUcDJnukCbfqLFrEj7
rfnE3zldZnITQ2X7liYGZWaR5SvfnOkqJg9+kZsH5SMvMBu7ova2Eg4WkblFuFkn
HFA3mB6vYooEzftaFoJu1mT6Rr0pEqrsPbi9XZkwaZVbfOgaYRn5XhR4y+nyw6NG
w152JJvdLcWnMo07csegPuiT+4BvPcNlwNDb1RInEuFIy1I06hP6yqNMM50GQjsn
wKBiZ1D37KMDXm1cqVrYxiXhpEbZRSeB8qzty+6nAHWJcRc9HtzmHQYK3mtOyfDE
irkQ8m62NiA2BdDVefhY2KHck9JNsNf6G2hw2KoMFmXs4iw/uEqBED2WNxvmW0jL
xyTHYwAiLravKf2s5W9SGZxIfqmmLkVLC6GX/fuGHsm5OZsE7u3+piNTnXVEQpGp
r/KX96AqmHh7FJayj3gTYMeyTEBI38edwEy7a5vVrg+Dhq0+HQm0Z0X7ntjQH57l
Vbt9XHtBGafbJE48N4yWExYhGchyNvzF3xK3MI4Mk2zqczifJFMmc9xXgmjagoCr
cC3y4Xonca6q0wERoXGGMmPe7sLbdtwH3VnpReixeQwXVcvAAW0VxyymAjOTmuDg
V8KVeBK08yIj5WEbsXG/1OLHmFuYCiP6D2dOpFXs6mmYctA0Qnj1P1rrFrTw1EpP
MC3dv46WnBnqlP7x/VexYm4O/DysasS0R6amTIr+fOL+MTCK2cRIGurrq/8y2dIz
lTrLWsd1QUPGiax0PkTq4/2bdueVZRKAdf09j0O8uJmzJ92/j2reBpTP4+Xnpd9W
Dg6NJg16DVIHQIXG/DkaDnpTKOXdMxCz+UL5i2UNIEl/E+4v7skEeCwlfV1Rbeet
a6vt43VglR3BVNA/WC+9K9I5XxUYC9BKAr3iSDqCH2foUY7wI04dqyNGM+zJm9im
4DAuSDYt4buyiLLIr+7fycahE2yIRAo9IZSMZEJDsnRQPmr8pLV6Duqobf7ZgsyL
V8SS5zN1zVO+lr5Ab/Cr1vyyWBRnGRANLQXt5mlNk6Qp6xRNMbpvt1/sECsc02X8
AxmMeodZ9rc/73z1opC19YX4X558JFMbqlD1ewu13iBh12pqJ8c2eLlZ8dnYLkqX
KP3fzSHkIAh1VZebdq2LjKMwsXPPHCo+37Ui7NoIcsMLpCdQHXGrqJ51Rhwg79MG
JDAolmzChPxWGClc7KNQCkD2I16B1OirJcaPkMuRrpXanKiq77E3iuXoEDFbqIol
TuNxWGUsyIcGKdOvWCBOVdp8epxqP7O5+YkDZTiyed8hQ5e31CfzEB7WXD+AJ/5Y
kXTJ1ZSRNASbUKm1mIWAWQuTCmQzDvqTHQZ3tHj0mS6ds7sxMWnCrTm7kt8buE4Q
Rd4ZZGXSiW6eoZgC9E64QE1hQzHW49JUio3P3YBwbTn9ECqe1OHEVa08B12XPYII
XfjT+ei5I6x0igZRiopi16sxkLl1mBjt09HpkRizlfl5TvyEE3zr1DMCh6F4z4M4
Ur5dnNTNViOL49ZIHQ1NtckwFC9aHfQ+s4i2y973VDP00DpR/gXqSPI2e5PaJg46
DmQCVri67oTIuX2fJ0+gLLpiMcu2egoGkJqBF04SB/G0v26Qd5bH+Rt5FPs4eGoz
tjMXzdFkfz3OwXojoXvVNC5CpS1lx7jajBOM0kzDxPAou18LCjlpDuRyKtse5868
VHEqEu/6XKXsgStGDCGnIpluO0TBH0qLltz7ohRUSV+8HbKrjf7ZvEePmkTQDFaP
zUbivqOY7+iJB8gLEuUkViUMJIPLqWCYVTCF7EFMk4908Z+wqCbrSvaFa/IYrdN4
Jk79OPaVj7UtrzmaCxT7rN1FB0sW3TZj2wkJYK+80ulEMgIaB7T8CQy935xFackx
G0AyDKeH21L5znku5slaURTuSA5MC9dX9IktORWKJHkvnlFvufg1zgQueqH4Byg7
evPngFyvp3YfSQOjHi3yxxib7r1TGqrQF+TrUBSKbZ1BLV2Wh4wNyXJjxWeRaYBq
JyRXDKI5RrDv8TZd7B38+NqkSM9bSPGnXwI+Rdmr23leLGuf+to55kYEc5iO4Qqw
NQ4CxGQUU4ig3hfn935n3IrihgpHlWUceeCssT4PlKbNb8/LTd4l+smLBDHm8PWW
+QuI0P1U2v26wTuqNEEY5xQPBjbc0QCj/m0axWYkH7kxSSEjuWBkmCksemmBH9u5
9SZe3x3OdpIcs3RTyCkspJlUr4mdFCixcfvavFa1Mo+W/Z9lDJdz/p3RVvDZv7Tf
RXnncs74DmfzvEBsihFgKwgpbMRrSLuc6wkSgVPMTd0wBS8GsMSQQTI5pxLjOUcn
j2Tp1HQzZQDqPN7ETlNeExTSSovBy4+Sz2GVB8Phf1g2f7WYeyFwORzbOflLxvqk
//pjAXNHBcBgCXF2eDCIgh8iRgCbSxdf3Ovg4R70Bf+OLqwRMgUoRVtFvgRz70od
Izku7aWVdLHp/HpdKFVMLzSo08cxVyFESL1F/YUZTeq+/i/dxJ1TaNFQR7L234MP
JCxjxhyC2WkNzqNHG215EG9byL0xzbi95tb9N3KwBeG2lZNt55skIU7dWC4OyeBs
Y6jCXtBjZFehf31K+vfZeAgocsSb/FIMENWcGFBEPOBICVVnP7kkHp9LJiViJNwC
emjclzlLA4mQkU+EQu5tfQsjIvHFfGU+4T+gadPdv+11Wr+PO/RisW2Oz/YATJSZ
3NweEAUvyJIbDuybtQeKbUkrJDkMDAiqTJqyDSjQdalXtYB+I0tmv+UV8V6IhcUG
y1NClo7o0iQfbSaJxl3PuJry22aPC+V3guCTSyBa1firGq81tcXLsf38ja8DxICV
/tczGv/PsMCr+onlEEZZ1drXJE3y/bFo8qYL5JycpEYbjDpJQ9I16JsN0KeNJwoy
imChe6vK+4ouKIbk4JYpsLnoSMyf4FJWuD1ktDf2U+2nsu/sjm5EFwvXUQSDLpCP
r0UAhc5WCpr7qjrTaELHVtBFLNBLa1NkWSd/1nOXJB1wQXnV3tW5/uyRG11TTok7
nthp6IrAhuN8GbmHBNROlpFCi9AAauCFH8prvPDqJZP+qjEuuQdP/SCRgEQqUOe9
4nhqE5FxY+hwK180PRaPzlDYqztYUwCExsO0ch2EaXzZwDxsv6GtAUtR0wUe0CMu
XCmx1ggDIovHlWn6Yt/HzRVUBIj9+3fKtHG8QkZj0I+aFNRTWPCYNxg9M1MkPwh8
cF5G1Lj7+kQWOXAtEUiYNS7qToFFu6bw4f8GWyjL0SFkOmXcDIx9Pg6GfnHNmUPc
ZoRK8uQAQh3v1p6GVc47KRX6FkxdF1otx43JLuAydcuCuUgY9yxm5jJAGxrrTQkA
6oooSeRZr5ViLCvr5ihbVX0buXaSXyO6DoqdTA5wAMfCJUKU2tKSV2y72wfSDpGd
dpbt+YTOEDaEFbRWb0g4pjO/TVydQUgwKi2ggRwz7HDi5JgApaXSHn/9sDcr+/UK
bBdGhhlESZ1CrlT9AYw1HWE5kb9L+KvYfm1i4cwVa/1dCUc/w8kgCDQKD6XPg6hw
679h8l1/aoiXrY/9N6L3kfVHeACYE339zV20npR5HkIymdt1BfTHScYJopnskDHU
BYdHfv5VIIytV7bg2VExq/0eGmX3/Mk8btSbR0QfmxydM2+GY8EQGaMBp+quTH2T
lMX/6fLYKEmkoJe7HNTJyjBrePrvszcacB13ZRwsjwFrgT4HC7hkmIz+lO0uV2wK
lAMm+s2QVn3ZWb/Kp/RLowEcd3HCW+nwVNqNIiawwLHHu9HhEwU24l/rxtp4fpbk
vhnz4Bx0SLCjWP7E3NL7eyKqRbyXF1G/YMSrJkbR8SxbbFTZSt3qTiyMDdrQJPzF
xkOMlnjrJojf/oqarQHdDvBf/IIKLTas1TBPUumCH7SBGle8KF3hf8BJxDJ6Wg0B
K5EsSGDt+3Chl1QkU/5+BvwTd37XJniRJJ9XJ19ncp7TYjpCZDzhIE5uCX3V7rZi
UXE9MUj4+3EF7yB+X9Q3ApgNLVk/QXzDRtbvlQUF6wy9NSO/V8ZEkjZOBGxNKssr
fN146kEwhIFZkdQxi36pPcs5dKkL8AI0KEEKfP72r5mLahYrRWWmCj5gu/aK625g
TyXgZQjfcscPFbh/7uKlm9Dg8DnxLwmelmqOs8JLo1jZoHhkTfB4xb5S1BngHiQH
KYR0two4MxcSPBPKLcnSNXLp7lKixnFGDxOy77c6JatHrXbGcLKWTW/e9SCs+/WM
7SPenlzA8yUSmpz2ztlRlx9Kl20zOmvF0/OLnqOVJASV0uzxLAIxdOMWS8FYtbKT
duv1phXJwzWNWuWVQ+26odLlxaosQqwcd10CZPEf05pNI5dgLlCnayLYBLmeuQWM
rLE8MHKcJ45cjqLVmZG24Vtclm8FIoAXxZ+xkFtaBqZfriGc/Em5jnk6TGj28xfl
RdIpyOHC+jwhRHNLbJiLraIWEI9IGrX3ac8ezmmIdhxBeiYHKWMkYCh4s2lRRanO
UptFlhsh0fYVi8gm8fuAPUoEsL/nRUNkpAAIqwvvdqG32L3F90/dzU5djwK3tu9i
CMdytYCm2N34RaJhnPViIX7T2lHaLXDLone1NGKZbEqDK/mkKePRDkIrrVyr4QTS
e9RnxUQUdpU3vWGxY3ktR4jVN8zHXPpe2UWkuOL7LaLj4N/+GpC0wz4QSaU4SMPB
tnTLJyMI6VY7ZdtOVFqDzoHKOua0QeclQ4I4Zm2cC46GpaAOX9oCmTrFuIzMCjai
lYN9TLE322dj6nL5dPJZSt8/jRtvhvG/MLeCZ/dSLUYGQ2k7ZtvIOZWA2ZyAEutg
7LUpkVglXC6tVd2VaQJ+ZwGQ/t0F1QTmgbGhRyZfStLhWqk7p7RNfbzP/PpHG6si
+gA6cAAv3mQcqDrMPWVrlbvXy9MhzqXfXKJUAxDElvuHdKCSH2QMmhcroAVH55c7
q7A5kN16C9SyU/9Ujt9QisoI8zbaBYSSim6fB3L+t9IzJvjMVkR8bAFyJ1n6cwFr
6BV8LA3wcPZi0eUjiqLqmoMIOG+q/dqSKjZ4yUi7SqZ7tpiIDBDkBMByVP9/Rssk
TNmfmo847S9msYMKUN4/LWtQzBwWqSE7q6uK3DtV/39PZBTEj49QCpk0lP3x2R61
AfBPDNQAa4kh3fL9wrZRKlemcG1Eff4mShskejmRsaawL4vlRsjw91fyKMrAKC2D
mn9gf+YvWdgsxboZDbFStThFCjnlngPKA85e6I8otX6s1OyRqjbK6dwHXYHqdQvJ
0pgKxAh7gPRMgZc6v20HFHCRP6TBE2o5pnLtmo/h+UsTUOOg1CB7aR6OEsCnDHj8
kuCDP2wMm/olI5T/ABV2b3lb+LiIWoA+s+yl+MjfwQju18D5ZoZ+D8RkObHXOmA/
nEFjInFA4cqW+LWJiGl6EuXdHlYe3H4uX3UR3SiqRSgcOqFTcFFccQpqQ9NNTuKD
b0DvldFyD2ty/OEBzoOrgv+xzRpT1dHRBK8UrR9yRPGTyVGt6QEMbsjqaBhRmBdE
g3fG9IvLG4Zs/EwNgNhmzkXbNJx3FX9RqeiXly4SKCfSRsWHedVD4M56cSLwwe5y
mIwW7yz4P+73YIgsQ43VklGuwk+fl3ZL32ZJTtHJ+zgVOjeSDpXru/ARpTk3iRcA
g8N2ITCXfbVBScbG8uadV4tDs/kmJ2dnbnNvwuJ+0M5xYP2ObZFbQ8fKfxi0O+0W
FBPrXAOGw7PUD7Bjpdt2GlC8DTE4ObypKqpKhJdZZgDSS6pKLzjKaZODyltudd4O
8ZDH6fwabpsYlBKlbARbUaBv9+iNOwnK97B+KG4yZG56CA2k/njwLsmeFAxTYJ5E
L1H+vpybOMve4/GTYfQ+cAWFfFj3tjXqOYHsIiABnBy08ClWIwoPOA5w2qTgCg42
qcFUIMGELU9Qv5nXknyx9DPYreLyRD35Pna8NOKcUE4epA82nYVe1kuFnF46bLIK
s4ctABOFJUIKMbiZqWDUEMuXJSpCdq5E4Y1LGH1Kb6HAWsjLMBrauIhb83AlrzBY
n55UDlFIjIZRdliDXDJ+qtEhCH/kQHK+aUgmeJgN+CBsivm1EgSdfWcR1Hm1Dqy6
3aiiYnQ24654ty9Z3Zb0EJqqNlOWWIUFkvuB7fCSlyjdPGNpKjU2OKeWcWoNAzlP
9U0G44oLy05Y3Yy4mq4AkYPVzuUgErWJ7GpFHsKidLFW+xX1/NzDaIhQJ2LpaJXb
cAV/6Dh1Pm6ehlVJKTSUTC8xyArPt/8prn6mLQ+bDVz370+zVXwizJOuRd0r5JIp
WjsG6RBmQ3tF9NHL/beZYPvbsypQ++TvdPi5CICubIU0nU1HIprj9olxfekeA9GL
9zUT/j6Sky7Ke8brd3ItWnV02ChZ43bXjCLQQofY9llCQqsoWTzssyMR42NUxmJH
6uMrHuhJ4n1I34qiJ+ytdxImdFDY1PlCLiO3pUUvDuR+zYQzLJxByZL7NiCi5hmZ
Sb2Z4czuMkDp9fx7Z2927L/+dQkhVXds7rWRROul6hrr/QticPBXSSag8H0WbrT3
dDSzPM1pcDwFu+sk1ACSx6hEW/qqgKEvdsTIaR+rVvnyOaHvePFNfBCzfVGrs8Nj
I/5XY/vekexAH20rX/Qvjh/pvAzUU8MIM2qbR2EQLEnxk3gJUZ1Sjsl8TCCK2aWp
RDpVn6QWV8HLX1g5BVVYCHLAKOFUzfBHCJVV9qp3HJkms7rG1CdE1srW6Em0XSNm
+3UY7J3PPeHb71vqjeSCAkQxf+BoZajUVTKngslu1/Jk+XWUarXcjMd5cLlMDPvB
sP+0ke8645ykmhA0OyotmS0PLEq+V/OaDxHVv//MeP5yk8sG2AJ/iwhqxqidR224
h6OztSp4dCtMtXUOg5FTljLZzU5JH3RZhXerj0l5K0Cz2UPt+C60niE/uNGTV89S
4bukGStID1q48APPC9nW8jBWgTxeOjtZ/zMQWeOdZXiLLL5WuKr8H2yTIZiwb5lc
qCSoayXdOZQql5LNQSuZMWBRUNdJ9CKW2dPzOKpxXnZTN8Yzs/OqUvfKjYShgiPq
fZPFd8JNFhz++BgnUuZ+kI/DoLab901gGOjGCnHFG087oPX9KTNlVjupbkcq7Rb1
+RoLQw9aB5MrNnDsYWDsS72/OSECxHpznBqiCKvBygST4aLICAD6u3kow8Dky3Cx
EEv9BvomLpmsRcMv5VuoLM1AQEj/h25ka4wU0txViP+H17RJlFEFRqjbSYmpwWcx
znRCq/P5nhsJWKQeTc/ZhPzAP659q0Cf5jIT7Ne4GSJXyP7IPXwHFWqdq+C3Thw7
lrpvWbxAoBe4p2wij3iO/IV+4P0IOy30oKq6/R3fvzCRNGN+HMyzgk/S82QHIExB
GM5S5U4UOC5YbkXpQ8C99AphrnJjNrwzNyVkaYkb2NIRnic3LgWG7qB3ys36+aGP
Nmss9NMUqUo5QqOn0fNHBpbhNdQLlNaF/W1ryrjWYiq0JpcL95PnUMAE6owhaZl4
Q9I5Bb4htmZk6wGlfFBbjvOFKd+TMYDLp/U0Wn0fy185HU/BYHI6omr8RMiNVyCI
ZplHolK4e8AfPNBbflkvd/LCefrAbk3MWrwJN12zao7YSX/srXGyYY+kT233sk2p
CWmv31WSUN/wcH1ddmXow8exfuVrRnccB2kobNG7/Sg3qdonyqowo7s9Dr3uCjJT
eNCNEceN/bNkRLBko+7JtzpPZht2SDMG6Wr16EloSyXUWPaq5rRcfsYRRlXB8h45
dSLnmY2eGKVk/7UxeAnO1L79X3ESpvtE2FuibTKReqNeR8fkvOWj2j0jlisIyHMm
JIr2P/FxVjKkerUCPF58PEg1xdx3py1BlM0vWOEw+WsDSODERR3MN4ncG5WRH8YR
gxLRffdSMQDiksrbAYJaysvA447pz6FOPfEoGZuc4jNgNP/GyIDsXUULCMGpfpXK
ixWGyNdogHCqlmVfGU7IsG+KpMhC/CIV7jrdBjimiTID3V2Xv5Lb+9Pz8zdubuU1
LwJfxqtkmU9ltwoIAzok9N/8JYPQMp0z8g35EjcPNhkSoi7SrFdEGk0RJZjMXL37
QZfcMwVYVxcs7GdSSsBlody+GtJU7kUuaGPj2oKSzWygNS/2UIxij+pioGCIznBd
xcjhOWWueaNLg6zsdDTiVmNhCw0yUQL/KB3cXTUWczX2siBGiEmbrY8C20DehOSn
0++2xMiaN6sBz7uxfLFZLcFqU9NDfsbJTXmCUjXp0X4N2hKqzCj/K5dFlzkmrTit
G7jtwng70zsGQeUycWP4SSrDiiD9DevF57k/aTkCqkwmkGGF9mRw/i3tIDNcaYU+
KmKCYj3xc0KKpMU979l2UpUCSvkVSmnXJXrMxSVCeQT0+MGZL+do7vm5bNNU2vs/
mNcK1yWrnB38UKHfcrk41Eo0kBpUfeb3fgjFQjDLjHPW9B13Ppbpycl7dNCXszc/
zY5l1YiaWQLduwewNhktDgtHBDx3S/Jwtwn0v3Jfkn61rumFDw3HkBEkQHWmqqOn
nw2ztXIa294Z+VIXY+Ga0ZJVPoFgjIQrhXbVPHQKSZfE55yadb7uWyoooP6kLGYU
zh6tzvWsW9+B0nOTHaEo3XVvWZikMW6wbcC8hz74OtWnuo+tyWy7Qc8IJq7efyRE
M2U8mbgJxdwxZ6aT5XzqOLMLjlm0c6K3jmGNLOOHbzEEYCokrKWXWzm4L3pj3OYF
PfXx/78qUeZAqDfuiLlquuQUnX32Nasg2R0wXGke7KMCabiWxKxkmRiYd+YZjF9r
q6Rt44w82Yg20cVicYG8Ok3pBNDenlLh4SwdU0siaA1B8IekWK79cUtd7oUgpLss
GCvG04Uo1PtG7dEOPVGXU7I0xLmXHYoJ9DP2INmVIKTGBWozIptcw0HgNwGXLCUy
ev0I0TCfXZC5kjHDQfiGZFzmWOhQdscjfVl7o4FkL8SMVMn5KiMjyRkbbNQ7CYUz
guVRnCuJp566x8QVcAdwZez7uzV7RScGG2rtFyCAv2yZeqxus0nFFCqmfLZpdAPL
7EDdZiDugnBm7SyMr5hvlaiK2j+hiyNinxNoxQ9/ysdH394rKpqQv6F5Y/RpD3T6
8BK4NsSRBr9vzm+5EcSj/AhR7q0Lm1ugtCv6CCNz0YjBkFnndgF+nQIojShEYYDs
BXIgZsK8sh3lm21/fWTbDhE8cBPG20TZTslvPO4xZVzKHGg66KIroOnuRMxml1+a
dVuTQi6mwoCLetaKfLZY/64gVmjWmLnhY0yKWRl4Vnew1afOa5eq8bJcl04NcVH9
O2rtr/Lq5LGfIbemCyKsQIOiB53kndnG3ViJ01ULiLTXL6BNAL1EBXSj2CgRIoU3
CX39K2iM8CcojBwwnZfleBayXAffDB58d5AzQvZooq+y76UpPLsUHk5C/hW8Yp8N
cDP4SL6DU8SzqvkT2UXNSiZt2A75z+xoAffp/oRXID8M9XHfq4o3RpKrOocmrv50
MPPxfrUxXY0y8cgCzUS1+v2P3GOF4ATqiqUd4+fyfBfrorG0fKDpkF39CeMspM7r
5JOjcWeJkRofTdoPzTRAx+f3UbpDSg8PrK/ejCm9hG1uXLrnUxmoATVRnXIxC6rR
5A4oOZvZxzG0Dh+WCNB8P+k33/sQAYJKEjkN9v0zLSWaHWwjUDxWxWf6YH92ISJu
lebpOah6djEEhxa7fnJY39eNR3Xns3X9JA8HNPu1m+ftz6Ch9sJJgAp2tLvlmPUe
Cvx6gMcvM3830RVMcdDsItjnkjby52ECHwiV2/SIAgSB4JFGXakW/6jvp4nY/Cdo
wIZQsPZtnD2SLWyfhePQKGpqxKvx6YwjxikD6wcmY7WPSFh20BAALxofbHEHj+o6
lVTiJKNxD89eGOHsA9G47b+p5+jYKKZ0Nn5rMr21ZmMTdjxhM9JEhGCqeSEVGD8m
HKs9gsS6x56npeviSTPaG1g4e6/hbYwxEoa9Wi+qg5JFMbQYlbtf1lTIuCICc7Hi
6yQbpGOEC1O3EdgyIdo/hS1bd+4TuxLLdwGFYD4hZtOO1F/Q5xs0rX7aL6W6dvG4
bBRLmN0Sd16iqvZggHO1Jt+pAMIyTV9TXMNcTXyWp5h1mhkb9j6jj8pTnoXuAhDt
YodWk9J5nKbWV+41ursbUZ1nP+tVzRdZLorPCZw6SAzG6Fy6vTimsoewierNU7Yj
tMN7nct1WfuQ1YOcW3ND6i8LhDcFZb86Tyc6mxWRSh9mPUQBTnacFXD7ZzUUdo7C
z0h3FwFsBCTbovf4wpH/6mOfodZQjwZAdIvDnZ6vWgBFHkB9+HFSXfjjypCpPdXL
TvFXX1GIcQHwna2Ns8nuyse5GJ4kSiaPT0sqRorIAv5d2OaVpezCBvn/+sVQ9OOB
tHIH0N3fq/zABQxCCgfnV8nH3VZpG9GV6ky1OrhxBTVC5Pvgtz7EDd3v8dmZHX7y
wamWyS+3w6clT7bj/xZj6urldgkFgtY1jokT+GFOchFB3OcA9Wo3Xn07jJXirQfU
BSwFA2ujj3LGSMYCW5gC/U/aam5ATA934errHcTDTwfqwnxQxcBreVZLn22Xrgde
npmO0uBdZ1oc5y0hoYilIkPOAFJacGqkZDETmATGFKVSxUpvx313aWEKl6J+9K8a
2D0o1eU+IGEaqdVIxAIX2mdwZu+37qItmVwo5sXKoyIC9woLnqvfvesmwn7oJDMV
MdUivG/IQQ646cP+RreX6bUXlxpIAWEdZqp4RtmDk3Kib9lkEZChWLyJJVHrt7+J
qTO2R4bNpW2OZm2uS7BltQoAMP5Hy8FOeTAm0vxWwnMrLPrFRCalt+SKLd3Gs85V
RT1gk4FsJaShVwvzeXBALoydFzVTH16ZTKTUQKPQwoCE63utk1vsHPVw0IPcbWBC
CtWf8TuO9k2d7S1A6Pt5x2Dh8i5eO64qiBhI48xYUmJw1hLPQgqdPtcw+YJTHfad
WMep22GXLwZdYV701cgTyKvKSDdQ+K/blsC4fix7IgI6Udo7L81UEJVqSv9RnUVn
CZkMFmwr6pXqKvYAcS+uxJdOwYxFJcLwCUGxDR9tTEqn2I6z1Ck1L15vpZ3E4N+8
E5tEzdclKDWn8TvAuunONG2OkM16RJByCAxf5/I3jXsCp0IjRb4ofoiooHX6Tcrt
phVXOr2MGgeoIZf5l+6GLh4hWJ0AJqy/PxFy3FW9fy1YbncKKdkGpL+frz1K4hbO
gbZ0+PTeh917P0SCxOKcDzqYfTjkeCleA0yrjNQzJh2W5KrEfFGrmi1SZUyKkUp9
gVCJ/0RUZj/Lc2Fnx0Kt3JSh4YL6IdvnB3gtf6ooh6ASIaGT1+VT3oyqV04ZCbSO
W467JIn4OT0xsUKldZ5cQJa25wIei98NByYnm/js+H8iA/1WPawoiuA3Z1vZlHGw
p7PPbKr9f6erjr7VkIhQosmuIrttDjMzkFiBCFHhx5iAPNHCp/+XazF+A3cIGXoN
qYEuprsaWUMK4qy3/D3WdhEXUiarIZNKQv3rXPmyC+ZTp1gryDcuiU/tHgxBocZq
nqXEbdb0F6ODFDFUZItTx4h4+OLpTP4yyRSBVZAk16hzLMD2IjgpUgNzgTO3MQ8H
9SkHiVKnaMA8eG7qUCnkHOLOqZ3COIckEGphRA542y02phgtcu/f6xXUX+xs78oK
Z/BR0b0/YO+nsllECawPsZ33+feuZOHXYnQT0QHPyK6CBae/z056qVdnZ04PVIQA
97hqJYOOULFUxusTrfBhBpApC5RgMNcNVmOKRV/m7IErXDPWF90rCKnZhvOVZ/rR
2WC4JvFgBR2VD5RzezHYuTeNhBchD53iKu4G9WR3gFagEV2bAEcXVSLbEzmGrkuZ
7Ef0JAWMa1FJLYbhMuV369xg/iLfAJWHEfXi8S8SJNNw+PRB5SQnXZgtn9elXfJJ
VwR9iv4XvjOrWSmaYIhvn7DEToIm/QUwHc+c5LbC2xGgJn2f4hY9Njkz1+sn7Szx
RhINHeJ4JFQTSKaaJ6eew3xlz1m6BsnrOhWN5pJ0t1MNAC9ToRW0Ix2N3DGqXRl8
4wdiUsJFm0Fp6Jpj7Z9TgGhm7h3r0BZjQGZcr+DRvvFGZ36KYrpjZDb8pa8+7zlV
3hw2d2Uey41FRVsqTEbUUhJrw7mzeuE/bP9+/wd6HhfjISq+K52ZRFYmnUJrDcVR
ZkIwKJ+3tv9MEdaeFG89milUmFlA6jMV3WqpGdr2UXVwlQHjSr+afSDyv/EB45Ss
pTzyuTP5TYE6O3ySqH9zKo1YI3TgUt87PU7NHQ+NZ7Uv4IxWdHSBkDxFfE+/jiHu
YLqIoDYcuEc2JJPzab0jJTFIux4+qG/ATWcRMMrY1dhgmcI6FsDzu79NtkqWdImS
hHcqSqzzPggvEzU2/m4MKgUDukfJYElE62yzCDUQmE8WteNZYm6dCPz0Ew5hmzt+
PfXpB8RD4eW/XToFzvfkMunchL3JqqLhLvh3nyWFN0zwQvM1tXoWpPTUUjuGpsst
XurDb7YlCZ98hVcKh1dVRxLdrsU/nDlAcFeaDZVRF4xKopi2/9dImTslDs7qtQyh
E1G4fcwChMYJTfQPHj+BPu0gPhfT2ulzTPq/ZMM9b5a07bzFKxF7s2tWa0PB/Cs6
VMIAd8Z7b0pyD+CfkRoWkZSCyTK9GQzxh0QCalOAne4OdQEAqr4L2NNK4nGWIKQA
n5YJGbifCqC2cfUoxif1SVR6ic+SLA9wzop99MozYQY9D3qPLXlSPQGXGdScvtfl
o50GGVmm8irEdvEzBOzy4tmvzvSoHkkuVfwUxeEC1mU0Dl5CFmM1FG0jDzyWjMI+
Nc1xd1Mg2f06F/DqoW2DrGnmtSz+WiGrkXdRa5fF15979+/UG5MKWSdQShmcXXo/
ayVWiQkLq/cPm8qX06Lj8AVMkEfjespGHIsd2xVQ22CKUGWQITOZLNoH1X1M0cEw
Lh7XyTFnP+q6LdUb5H7aH/epW+jml4yE6wBNlUlZ2SQoLbwGK4FLgPvM19gktFc7
tnNXj99HWcgAmF9pdU1V8iVKHontQWwbhIDFx2bxNUOOtcJBB5ikHf/GtwHgvGp3
4za92sl2D3vzEfEny1TUEg+ak6WVahSUd1SdXM/dtRE/Rc7WEEEDT2t/nsaOGV7t
cGOc7BJTfarwSk7V/7eCOb9HOx82FmpANfJwCHNuMNJNWbp+TXx+JtKyWEH/xt/M
1/18b4DHO5lK99KEzs04qhJrXKF4bG1UjLxNy0WFZIr4k5OG93nc6qOkDqo65rIv
7tqnvA533Y0ifn4Wx+5YZvpvo2V81X6jAV1r9uHhNlRYBmlQkXLlcnWGojvXjOXa
RtP8ziAuJ/vDAIno+8tdqUmhaBa56CP2yVPwZ/LqjqxsySWDjgoaj7RzwhPSiejH
PXYJduqCWra8DtfXZeZHNaLPJ94pqyPvOEKZiIwk1JyIAWxGr4OBSZredGIBokZa
+BrBKz0ZXzQM15i9pDVMVSKmi35omehO0MwG+vaW70rBOv/4EvYwMZDrUl5Ll/ew
aydDUctJQXewbC2c4R5EcwiRwCf2dUs9Dwv6mUEuxrkknqaMd62zVJNJ0XRPaS5H
yNY56JFkn67WMdwdllnA3XoqpOkUwnkfLjZE6q28QcCwJPcrLpLO9tE26ZJOrpow
k0zeDIb61P5VeQiOmdyTYEUNIIeKO+rrIuIbYImonuZqFr4eSKROw+I585rHmeZT
kmZg6/kCtl02MCINXp3Q7UQgadQ3WgrGcHUpKkHAg6dpGFXKsIKvm8PuAENvUlTZ
Mx5R30CouAA8STYYoEG1S2tRuBuir4F08OzNt3cdTGp0+3Fi9F7pQzpPP6MqTJBM
Bxt+1MtMTGdXzbzZA2z9Vkq3wzEaSSIXP5fsimWrTxGNbOoKB+NdgxYTth60zniP
dhPZLa5ceQAE+xrrJahBNM1SBImUkp2ZoRzOBk78Gp3pMamZXy4CbtvEXfOLfjMX
95o+U7nV3WRWPp8XKIBSwcAeKOihDtyRDXNH9nAKh3cP1ES8SRmztV9wmoKbvnzc
z4K3sBEDQNHF01ILoyfCf/ZUTRMpNK5nIpCGQFKwMNJTJZxDAXaM3bpX387h9si0
Ou9UYVKSYKSDXX+VS1s/i4XuaPBfLV+WAfvxy7flmxEhxlJE/Kb6bNLHtYP+j1lT
83zhGG4bbP8V8zU5KJ6YInmw1rga7fJpOLsgDNr7RQFG3p0q2NkgSG9AbSf9KLY2
zIJAGwxwagniIb3F8tj871gcM/zQst+WelnOtJDSbEYfjp6mEE+qx5xdpwyIKxAM
cQD1pdcbiDL3oWf+oV520Xk0PAugNbBoRh2jqIm7rpH5bN5TD2ZZyxPopyQkeU2b
KkMLIUC2IdtmjN9KEJds0fjRwtZclexoZlODUdQakkdUhLl/xDHYcbH/ocE7QAHc
kgYTd59fze3IfveM1kAnFphnZSO1l0gG2LNm/C1fWU7PpCoCo9ph5HEWOd+z/TMn
k/gmcoTwny/524H4kkCmweSWXuBax4kVU/QqNyiPkeQzjD6v2Yf1bk1Yk7ULwsPB
4aHrq1wji+iClFvt8w14INB9vDTX6WvbteyrYJjN8Xoi01fYjfores79m6z1c2OI
y03R1OMSR8PNNO6YG03eAeo2EsMZnjQ6BAjV1G7HoeWc/YpBUMN9Ls/gcTIlNaY6
+DKuZUl0SRdl8/MCMtIuHrd3ft5Yhg0O2ymBoHez/unGsYbgsCeIFs1HvSNx3bwr
2+DbxMumhi/FrqRMmUH8LHsJJDj8KBTMBV+gEqeeWdaqnuCiAH9fffLn1+8zb5Gx
YNlZ++Nb4cTD87Mbnhmff9vh3YhwgmlabwyQazNCfC7vfJDJ3zpGlh4Aq4SDzwdu
zXEMV0pIz2E8mBPDIIaimxigainvggoR0Hr+UFQY6Xu2Rx7pPGLDm6MQefhp0egA
HVKcVt6DDKWUCorqHrvA2JzkBgAXqyn5LAed/A1v3JCKrdF4LdwJQhxKYgKeqH+6
ddInYS+qJEnQUhvsCFx6rZBABYMhBRrcnOhjGMjYitnWVtEzg7CL17PLUq8+buaA
SD/4xEvtLgWvJXNzDqjxLZUNqbuY/XVQHU93310i0PunZYhb2cTm41sTW5vmRcdS
y+3yAm3UEu7Th9D9TkNNlQz5IS5toY3ge68Ett7W+woBP2g0BiknFQfjJUTsaV6y
tu7Mi8CmQDDDRdjB9q0FyOFQ0Xhpca77qdR5H/UezX4VuJEZM0P0DOl+XPg/SmwD
VDFbBFL44sl20ZgqAhOMgeYyiOr+bsyXa9GFIsJoYEUFbWkdtG9g0dSVJzrmLs9S
VKJMhFQULVMfn4DaRADNHQymSdsrn9Q6+Ig25k2TTPwe4IWlM1FnumJ0O50J4lZp
heWc7MenTztsMajnRO1Uodqgk0sa2DH9VAWGfrY5F6P1rFzVYWmoRvmZn+wJBZDq
eh6MWLvIddhbYDgNFe4H8VZP14zpwcGl++ntsny08Ti/0MiiQrYy5w4Id30JJKBH
0XsdWmr1d67IGxYSsnCF7DxIkTw3GoXxQcGeQOS02KjMuvFUMtgpm/pfH7z3JWCK
kBkPfaYquqo8+c6YbaiGyFuSWAqcChVaLwMXs8ZfKXbMWLI6IO1yCFDXz21pXvBY
Z7ygF40/KP1SOYg1XjZ+eH8DMzrkfrtZvnY2xQOiqbcMs0MThgTQ9Kox27eIiHRR
dW5jZyrLSrozSaIjkSnCcTFvuZWmJbbJPLgpdtCdW7YNBonZCENaQX8S9nA13fgT
H7R18QqnK8nwysfCLAmafcAs+zyu3XSMlRD9MRntynqK007oGW8fT6r/isH4XiJS
iC49u6UEULKlGsTSn8rzVa2Hpn7p4XaOmsb+dqYlKVEkD6LgHtv51jBtekqbV91U
CjnaAHxJ0WltVxGWd4BNNO7EWGkuVliAfzqmCtAfUtXNJSAyaL/8bgQCWeFE5smd
2GqWT/8z8+602E0JmvNJbqGPconO2wsGjMMFyq/5C2HdTqciGd7oJnqqykSslmi4
f5rnT3nbCfzSVTQFwDZRpnajFlrJ1mPmWOsgoy7YcO8+HG+o8PFwoa+Oomsaokd2
NGHOY+3NKKLm5glMdxYBTWpv+kvFUqKlZUyllSSXQDZinUUMkYUTeyw0Howg95QY
9YxKr+Pr4sPvcOcmhd3hlImI6XFZAoUZizEu4/F8d8WPRUnHnOPhMNRPXlS85s5y
cGfm0r347vs+7sf5A1FldGW4q1ZjO/w/LZTp6Lxid9gwZEP50tvkxY+W63J/F0je
GIdmaNC/EuyVG/YjKCVnzv4CKRI49QPEwwar+LWCvbp2Li6MdN8g0aMn2cX6gNCP
qHom9FGS4GCQgg1kGe9k3Ewc9xohD1s2jVRB8kR8UHbbRmGIY4GlaEwzec92EOdt
mFSSphmdGzAZhsdiqH/BWA63P677MSV4ScYqHAOhD7C6+im4/NlMg9uPVkbCugmP
exzTSBfMaIWMFJpWFT0OlD9GjaUSCvzdvT/89q8pVfu7voDQeEfsgW7TeQxSDUva
zkKWvmt5ys80neVHOquTgEKKE0/nUOcY3+l33P05Iz6MFOrBt428sgMEMHwfLgwF
dVZmYIQVofLljgjVdbXYii3Sv0fGPdR9RVT2gjeXVwBjF5QJ35vI70nvijSrHDId
J627sLZbeHlcpk4K0g5nFqDzHOPpQq52JYwIeo9lZOuVbLjDok0eJ+xhhmsuqOTQ
8vKc0EUuNJgyozHyVd6BPdb3AGbjYFYSGX/Cx39UeZjpepyrXACraa57NSHtSp6M
OuAmxJ4O4EGHNJqHctznz6KGxC5WcEQ8h8OTgzIPqYgbQhi1nyS1AN9jhrzul/4O
a/g95rbcECX/4GIjzHsfokyVlkihEMkKvb3ttKsOCLKzfmwfgKZByidLhdF3S6gE
NBQ/aBFq1jBgis/Q5SiAO4UiRue/7SXT81Iv9Y1CVH2BJlZp0U0btcgLgLuQTUw2
ZUyURpvMzM/O7OXAJULqyLAquqsznq6nU8lWGNCUbdIKrxiiO7cyB1uLScisjeKA
Pw+09OsmCgiQlpXfTVR/+/NCWrlis5+cg2UAQ7nnHLK4G7qcqIDo7tBJBIRv0aO7
nfOrTMq7eUvnZItzx+RabCLN7OxGug5Z/N32nFgUD8SEpEJWOfbgFg88AN/I9q/Q
4fkMeXSCUwymialiUkZXGmstQEJBGB4oiJeP/sK2JK5fHyJjbykzPumQ3heNBZaO
c9Ap39DhxeWF5iGL7BXANjIy0asmDSfyoSWjsdZMQrG4sWMHCxp/haO2eSQ+fAfn
6hpotUmUDvZWZEeKOVFoKT+xeexWeM7Ra2NKfSDrLLX8HbGEuz4bMYsNdglF/21e
+7vIirvkceJOL6LQ3Dsgjd1LC6N7KB6uIZ5MZHiaFO9ZLFBLhZKLajdCg+u8tii4
9Y1kx2KliHr9cMOq9DrPPLkozwzgQNow7+rKoOt5xTiqA4VZIDRga+Protjq/aA0
MIqkY2l5jPnLfAwfkibiqrTI2UFkqegzciIjvWAIiBbzl7eqRzcHBt6PawEXkPDk
wzutpLuZxGz62NdKMw1j8hd8xOqP6pgYKFxBXOaATErBK1vHQrqMEVTUg/41haTF
XlUTFprs23WScsxNYwoZlnZTVW+CNVktSDzdxy/FYF3mNrv37x8xt7hxpnuczYZ8
rdctIrnpAoJ4FEoGd+2SnqqCWOG72OESCKmwHRu9HzFEXMONQKMYdw2y4b9S5IQK
HD1J3vyidMTYursARNDn2XVhB6uo67AM5Y8mUKs0PHxPYntWTl16Mpqdz/ujbBuO
1Icy4juK+EDCtij9OwV9zGK0oV13w9KVRkZbL/FElHi/qxu04Qfc1rVKEGK2EMLH
XDPyRmUB/S+/2D+b0SIQh/kuuHLQjTph8ZBvoD3vLYO3/z702a7T5BsPSyA5fZoG
exJNC7y50Oc4dW6gv+r+iZ3rbJA+FwsldWAVYX6+MDCn+W9Rh6owmmHHwlcRq1dX
b+Vq4n3c2M8aBlQZfiRspfdtZQqQRRfj88dX10D/V2jm7+xE3nZPu4AbXUTBpiDm
xXd690PPUi4thMk05Mcndhjg7YVbvsPzwSX4JUfCBvrOD1cHr9gVVIuxj1i1uDYw
LGA/BrN7PtOrFZNFYAJMIhieiNbovvbGFadf/YgNjqsLzd/teDlpBZt4dJrmnCkL
cFssb2QLTn4asd1muGMMdmUrw3jy1w9kniwNu+auBXFmoXcUzWHAtc0UQ1BaJ+5U
IAlsdvXAW84LwXqh0BqiGjMhYg8LcaNXkuvqhZcaVTWv5cmQQOgkdl5mogsxrCOW
LGt+YBATooIeNHoskCfjilXAYBMD4Sk9wORXog5UP5AeCzlntc0g4NDfaDwN/wfD
rAcqd4l+bHnDk72FOUbpi5vXaNAvcI5n1k4aEwcXGHjH+dTFGq/E0K+yjmZKbvVS
O7Qu2fvseEi+TWVGVsSVP/wvUlvngQ0K2CbfKGS27Lru8Wtv6De43m/bkQWWm9KD
vipZwN/pCEwCH8sN21uY2PqbmbXG4VwdfF2ykyOvLMPWU194dB8B8IRleHVOcyEb
Xu6hWsWlBVqyyIaVGi9zRCLl3cNen/hL9BPVplzs4LxIbPNRZ8aZneh9BBKyImvj
+XEfglVsmH0wSOmGAULUsNtFfRVI5lh/OMn+S+FvBhSQvL/nT01ovI+rkks7LNjv
HrexjigaK81wmFnI5CaLMQV8gU7nGM/UGx+okut47ajsfwGZUSXNiokeDrZdqJnm
QPArFuGlF07WXFEr1h7TMTEbMIbsnspbDZLyulYb0wG75mPXqI/K7EZmFy9edxRm
FPya1KEkhGOYueYITWniLg2K3tHN9hB8vUF5J+XH4nKGdigHwi54VmXZYEABYcZ2
iObEg3pEsgBXACE7W7PooLVnyfab0cVEpsd0WhXvHrOtEtpQaOL8ecQO/jtOvhoU
7dNDws5SIggP5lDDpFl3WeYY+0yzHMFtosv3+N4u4Cw0h7N0yCrVoDGVUbxc6Ijf
eYFORzFcUFBC7xp6DrXjU2pDXvWovNPABXHMjO2ykcWQxh8xol8oNqvp9AsHQVT1
wmkFXiHJ2c/CczK6kHS1Z+ZEyrX7Du/Hp205PLSIUr5GDB80NlQnLfBwUssusA2d
yvVvpw5HPvMX2JzjGMVvfZ3MMult00jmEbv6x6S0Wnj5092h/VdWqmFb7zkBmLwA
p44c7/dXwhvXCIQ5KljUCYTSDwQ5gRyVnSfKVEgR0XLQCJfEfoqLVLN6/7zolJEQ
unuDBNa4upCqzaW68NNU30lwqlnStuJeZ/Dffj4tY0KAtL0Wq3JMUWruxWsckCoW
ns+ZAB4ezPUYAsq7VOF08yH2hSam3rN/1fNfsERKg0OoG8KJUsdffRo1PfzCcfQU
g0v9fJLKm9MWDkuY2bbZVrDpEWKQvqs+DklcpG0OYRr47ezwcgJ+nBTDvnwfc0IR
uoCjhcqVcphQwmDZUJ4Ne1JvQVVn9yKf2CY3ArsIFIwRjGJqtpphYp8yuRAo0nBM
KZP6v9fhlb+PxhP3qvjkfQYpVZKoqLbO+avDTSHpbZVNuwpgvr8jpIws4qZlwBor
oNXuvByNVlKGtl55vJP1wfKk7e4elgMgnp/mn1k1j/czXiEymQdmqXeSvqsDjDIo
c8ZKlO5/YV/l+47TgqBosO0eoYcp3gzJP9Oz2zkpWuX53GCbhU2RMsV1IYzMwJrz
BM6eKpesuobSKKOOQ5cNckearNnwbXsr+LU1R2XwjMKUzGxm+NlYbG0ZlHmddekR
aoDwOXWvnrPaKFgQspI0GbizolotNHwHWVQKbWD8H7uNTbdP+wfSSrLkBoDYn3Vm
B2dnOXf9ieByTu8TgKlZyspLhofiDAYmyBtPFHB1nESOs/mnMjdBdf6WthkcfZkL
Y8cGK2COnCPxS8MUq1pRK/6+8n0vuPXndhIgaI0Qw1TgRSppSiYepZFHt0gkQy7g
7RwPdi8Yuba1rL3rpu5A1MPWpYMqBTRYZovZICD35Imav/gJHvbU2HPy7i4TvWrC
uy3b/HZVpar2suW1s9gBSQCmfEBAHsJqCb+GM4S8zuHX0IahMdOGxwxVwOPRewgX
IpoLdPsPjyVYgZrzS6FyJZv6ed3M+WsZbXgQVr3EwpBhSTNzl1HlsjqN3kqUzdMv
6IGrCkrKJ8PejSRBt+jiDV0p5UjJ3Tl5qanmaToPhwdvHz5yvk/lZkTa/xgLAl/l
b01HGJBouJKqRVCQ45SymRmnAzbFUsThU7OpPvM94aMLpT24JmM3/gdnZ7ZPT/5W
WZPJJfyXM4yGZ6BwnoV6GVecoeqU08tCshExjJ8Hy0nA4Adkfqrn5R/ucGTd3vQb
DlLwQv8l4fYmd393d55NBtzqXQNPiEo9z6j8OUXxNVVoRmy0mnjkhzrLK/HLwzFO
CuB+wDLd75SN9hgw+KJQ+L33oGLdMc9pcFUcE30RUpvNIZbbjzL8OfNUkS2vzwFY
bBHvcOYdBWsx8cLlXc6FP/rhYeV2cMBSEXSdiUA+nirA0fknlyXiNRJzv86Oknr7
5s2pfDJg4PxLU4qP15Gi4ZKG380GooTgNF7kIO05LPUxhDnFSo8AyZCWfl9mqBJY
s6jhKiDlIC7+624cVdmh6m3ebVQzG4nneAXtzZdoBD3+YM0LJ5ZVcfUF2hPkUiRn
OoI7sDakD2Y7D2Do+qs1I25i1lgKZzQxDwt2XBlfISFNPKf3xZQD93doGFiI4bX+
3ch2ygHCVbFepoZ/4IJfUeWqC+Zp0FEwjXOaKENl7QA/oRUIS9tX6EM0fAGCPBsP
f+SpLwiyK63FRlZ4zcY4nXewezgVDYUB4eWXtZ4EFW3KXghPO196gJqdsvtVmWnz
Us4aZZ3DRgzdj+WcbcyV/xOPfeMyA77M8lI2oKkpU1ySXNdXQ63PLnogkE5KO/hM
77whY2UCWyT5xp8nXWPfFF2CqN8cgZEOqRr22o8EBEwrwaeDESfD1ZixmLgOQ2Rw
4hJgtlfinhfN6bDhoMXjHGuux6cvm1xbLVwsL5cYKq+8UkoB7v2W3+ySbtflfw2I
ZfMdgfDoekvE3EXU7P674/V25343CHexfy80usUnBRJFKjRf/jR1cb3Ddquv4oY9
aH7rk+L9+HORlSjDgzgljbb7UKjqP9H7XEk8rH4pQz075vJDT3SLs0YsYWYRfttB
pNBmoEIIqks+wMCC/DKbu25MY2mT9z9Hoh7Z621/aT9Gde0EzF0SSRfmU9mLPHVp
W+fCJeLSIr9Gbq5rfIiQskgq+LJx6X18xcJJTdiPWRsY4U+FSmD6jeN94xRSWMzB
msmyUdSJSV9P1pcvbw69wofYvGfXnpqxYDfGrosofkWWwlDxA6dzuhKGdpxcmohi
lbtmqm98mtclZumTLznAjCTjKseLvKTqp8OrOCUhL/uG68+roDH+uc+LbF+bnirI
nVHyREOvZD0qKp/N4jMC1kXB84U/LL856DhDfXvqNv+Umb9yrP/mSsLlmwNA7cNG
+0pKnmtLyeYlDkWAXJd6P68FrSoAnYfClNtLXtUEFVu4Wbl+dWHFp6qqLmPQVXQF
ZZWYwUGrV/guqG9t1KZfd1SCmSsSt1Bv6mjcXoSpqkXeBsBuyzOrzpyqXTY9Cjvw
ouruJLuu3zf/PSh7wUYDNJZDGGLv9kmdz4oDcKk09wa5ywh+79hgtYFUtZ0m4Jw7
dYR3H2rg1Mwx7nJ17KnYpFLyrGQLHsjH9TGqNpLFEwSmMcSmAvTSUHGQQwzWWMTy
ukcXEEcSAvpYWM+b+UAusOUgFrsH0ZzYPt123eDV3cXiQ8MB0IQz5+oqKnA66fms
4okj/8SBQfcQRQaardajrcxzJy9iM/4mMozPPZbdeOfoIzyZvxfhBm9UwObPplm0
rBlIH/EOeNvLLz9LZ1Kf+DifWVghpjn5AyMtdzQguz0zQfuZb18SnRGerzNzGWRh
yHGRvzjuVWmi+8UoPc0KPCRran7yuJRWa8tRQn1ayPsI1ZTg2pFqQKOCQV8Bu/AW
XhOx6PZJEg8bF63j68rsurpon8ek44nyppuJzayLXSt6fYbBonInj3xqC2lwLvOt
ugjO/V7gAjZxgtDJqeuUyv4wShfggTYBacCYzEWBQoIPhKgBFkfI29vdDcdV42h3
kPhW9FVW3kd5OpUJyVmv3//iwkggjPzZIlmEQGkZbcCL2PhzvZ91NJe/PVx/J6rH
P/KSlT60NUcLSYBfn2zyowxRnEeW9atNixk59rXjzAnrCmD/qa/AF3E57FOiiT8Z
G2fDLtY0oxbpvZm+UuXkEy27rTueS6o0KpfgaVMMOGGKf8dEF7bhNvmdYcwCF17o
fE0faqIcHCxz2rrFjADrq4uOq+yKNJUO7hNyuRYvzPNQtCiWBC/UE8HrE1UjN8Fy
AM7t54xKBejHF6Ox7RCXX7ZmcHWrAt8UqP0oHz0R4VpjvnTYPKw99/rtMegN00y0
ZDpETu6z0KEzicwB29TWL5EEbaEQFDcehy59U3Ygx1UAb3ivx3kNJNuzz2cq66lO
Sq67Ozuog4gMm2rmOaO34sCWFvKKQoYUgvHFL+bbzhOsPaaf6dF3zQKkUNljMUS9
Gg8FmBQ8JTcqeuxE/v/xm5OKFXySOq9+TfzdUZVJ8JI0rnXU+QHk+UhwKbV4bld0
/tKprS1v9+OSaub1BuMKhhF2rVIv3xC8tofKm5GEEkZfmdWPtT320Ii1xJG2vlNC
d9SNsdJBBdV71yxZnW+x7utS1AddfwMDBCexpWjDtzFK2bjNTJ7UKHRTomUDSevV
i4CgulbpZiEizzJahYrXAIk8DMpWSdUvSNbj3j6naFFPmHrYwDI7x4K2hswS1ROr
onSp/BrgfxkA7rmG6hJ64xJ9EcSeba4E20WqIs+u1ksuVqQkwpae9QPY2L4kUpuK
AqQuB6mM0eHv5zs3sljd0AMMmAqfJHBNyrogPVWUt5VI3OarqcKIdI3sKfloh+CG
8yHQAoM7A9bbi5UwhJn+90j17lo0Kc6KtSRu9zMK8zvihQt8KuATSI0kLky+9F1g
gNmrZk/cJW+noMF8qPKiMSdHSORx0eTEr2NJA6jEzvVCkq7w9tHr8U8p/XdxSbaH
aZhWxohACIamibRxtYkS23vz5L2FDw33x1r4sB5ALRSu+OjNcC3jZK9isIie+YTo
tFO03jOK2BajQHgXVjJtdhJLmIp2jQIZR0g4Migc2wMuFfrkQbKcDDxr5Hh2jQep
GtdVZTs243RItEUeBZd//MBWedXGINM2jcQ+IAti+GLra4MzB5J5HCz6QvTPDMkP
4tJBGWpVmxA3SSbP8uQg9dsfZ+Mxx5FljpUnJ+dL/ng+ZhucI8aIot3SkIuk/s15
bg+cETaV0U+RiAhNxp0+9B+etk6A/IMr+s1fLQJKGw3Cy2hkK3zGOFRzKA5rp7sJ
/qwe2QI7h4AWvcqCKMWf0TpqwFC1iRbbQsdcB/BqXPAsxX1sfBDuKJgGYuHbWjTu
Fni2dO92oGmOWtvvflRGrlyI1wMiFxv2KRocz8qvta+yfhpnLt8/JAYa4DYwwDtA
/PkYhRYMxhMqA5h0023PB9+n5QBLY7S3P5oYnCc99hgrUNUiBQHULiaS/UJkEn7a
v306ZE+e1T9yAySLfxkj6/+xybssmeZTDWP6gJkzuqptIEAJEuoYp7OEZ6finrRL
a8LSswwLX1nYZqF9cF75HMrJ+5DYK/tfd0AF1NOMIl4lUxbhP56lPLUnx3kcHGPv
MQnyXPnIIH20GJ1vyMrXi6n6b/mZLHh8QbxIEnk3ppwm8n2s4Z++hlKNaQ+461At
dZPuAiDrC1Qom8AJZmU5eH+LxwgU1m2j3MMSxR2NrvydyAMpRFXVQhPwCBYmKRXY
V3/0ZiCrVZXWv3ni7+n8k6z2VGTAnxgj6oRbCypn22ILXKpZch3VODrQFalu982k
PIERql72zzIkzzyMv3ky/Lo0IInaygtdD+lmPadIvUXYoMnDU5FrCUD+T3+Wb5D7
fph56dBpfeUlOQ6QTXVsZMhvXJBPk+tFgc1UGjKNj7v4cIuzIiy216IJXqfBa7zY
WanRnadjxWMFqq3SpwmCE1jUxtHmSiIzQB6YsVo9FfpmHROEOOSeXxtDINhW8W6j
SQC1jXRqqdsugRp8Kevqpm9xs4Q75eZRPcT+i9VJ5rTpcb89gObbJvd8U0O3jmVo
+4+FT5p4lfKFl1c1nIY2ky3lr0or9/z5aFi8tQnwTxHdMhIr1L87vMQ191wjy6wt
HpazsizclSBUjI79AsYUiO8PmbjZAsZo3TmdcwAA2cJ0o893ARV0JBs5DSrlZiou
8h4pjtfLNoq8FNzPzUaaUZ7qV6nuiuQs3UHXGQIJas6OUi6FfVd/mgK9veQ4Eu6Z
gXNpOUFXH/9U/uVz5n0rcwwNQ64obirIR/xWCu3PmXKFOWhP1ovLIKJ5v9H5BoY/
lVduwxTUM08aPEpROzTCsxUfTIyTbYRSv4kAzLprYbAyjSwtkMyRpHGOxhM1g2eW
7uIrauHY2ZesNIE3v9BmW2CoLyaygvknQpFou/7k/hF6kcLIfUWARJun5LL5oRoy
OPyToqzdYl8OBNaellfh/dnpbQ0JHh7TCmIpq4UDfquiO07i6PvbpqAOCdeFn8DE
63lEBhbzc60370uFYtkHbzT3V3zlNJ4afUC+RNroGnpP0UVytdtbFtQ3KVLmMEV6
LStPFKvVQQgdvHFtCe9pGpcj5Km7l9HY6ahSH8p10S7VZFOMpE79WvZOswMxMRw7
c/KWbEO7rAAAVr7oiNU2nYg7ejup9Zec9thxt+ILrXOGi3QFd5O0mwfHi3CbtilP
h5nrelIXus/3ukyyfUrcdwsppAFOeMVOyagdUuu8cRz/JNDzmgmJuR1Vt6MvaS5b
8kexZN2yhbq9677VJ1SHHRIpIYzmFwlfIOwP/IEV8SorTTRGA292H0TYXFg30/3Q
EsHiaNDjbcVuKQB+NtDtH5GuJz/YX3iYuoN0Rh1gzFK1sUARJGQo7CZFJddPscL0
XAnkvlTnztdN2Sw98Vvjzd2z8o7fjeCqVd5ch8IqEhe6bDdS3hBHNIa5q4cF16uW
lMK44gh0w2tM+JJK9n+2Cet/cwLcqKaPMcLgqqx/Fd7v/owAnz5+UQTVRtrCNOG2
Ub2kC/Wvz1o96y7MWRE5umP4tI5cVlsj4/wl6eBDZfv8tSBeSQDAY5nyPpFNg9B7
Yz64q+XKDs4jRdYRck1RxnsyS1raauEtyPKyxjXCPIkzcTBmCuFHzYNzftihhVq4
hS32+bF28a8WY6LytdBGqgFe/ynIorR3KQZad8WA1pd3ktx84uHFoV7nyVfNkwZ6
uegu5ImKFb1g7rsI6Qw7Wte7pIos07tvwhFQgZnWa6s2biQlVjR+Er6gdX0+I9iH
cA81ypE6R7DQ2SEnb7KmNul4yovDc9RcYXPC7TwB/W80vxKmieN0q4wWMHuDmNOd
3tD6qINR0CdxdUnTXGKp9BMlh+A2Vs3tdEirOFLREdhqSZbA/4W2SK0YtSzbLiXA
ZaKtPagAsQP+LdhUxvoBwaYZbtgfMcvsIhmaraKZOfxXzyMHRJyUQb4IK7nKqG9h
dSAj/37tVKi8i+xbQ7XGepVs1L6pQkni0zoIZgTJhZmZFX1EmvQRI6bflSEVnTu8
dtGGABdJemR0JyhA0OW3J2Nxv7tYFh5AcOb5GRJSMOoN7uCK/6w3AJY5gzXf1Fwp
VdzBvBZZtq37PrNgXI6SJGDL540QcUdLNsAPKEL/B7PZHXzk1B7Xk8xMUPBS59xb
mL6A3kU3zpQVx0XTzVv3yCuUqDP4fALMIfHIP5kDV+3TPPf+h3pM9OMM9Lekclf1
9F2LkjVkDx6uuHnj1XGO0LFqXUUvetkkkBvLfWfSxQW+APq+bYBt5C2MyRACwhaE
U3lPQzPUm+bVUXXYe16r5GyCW6Ohj7n6Onx2Pyawkc4qcrBTp2uQ4pTd/fBrYS9a
AR+7QDBz+6GETfN/ztQJ3+fELCvQaGUzdbdtRo5wK1CdbV/bBX8dapUsLMPM6U5S
LKOZP4QtULmGPHWoAacH96/TRzG3L+XFpn9aeEFmTDOI+dMmxvWrRvAB5rgEAUwB
7D5wQixcSxuoRXu0pUq9SjRM1Bru8SFAgbe47GNpQI3iR4iU3Wi259IU2VM6zfmi
ahcJ/QbM5s2kr4E+u3YCfvn1WRD78/GnzkE9kYtoadMpgAu08pGydsheeqUhrTL/
TzA5OzftXQ3JnSUck8yKJ0rnL0liqGR3aNTEES4Qc0TAeNayOC3MpkWIbXqwQgeP
jaTjfqh6zdfYRPD2fjYOjKggP05GsU/fSjvD0vGp3AdnXLL08tbs7NkB7LrULR/7
gcBFYby6oCHPNOMdgIkZmPwl6DsdUBSRWCeBybZRR0zwvcT86OLgu/8F8sfhpbOb
V5JmiXkYqrHGiu3dm8CU2rMGVKMxkdnN6CGtEaQJm/byrwuk0A5ODS7ouDtptofg
LBO42Rd5YdOOQnccLgExFRqL+7XybPnnzqJYY+vmKzAn0I+lDUM7dITvKDoRXxu+
NMhwtx3hB7+g9aoXxR0bW3p/3qyyBiIQt2SNn81ileVAFmVFU0Q5FKAoCpCgWhEM
+PItrR0I5FSG9S/xwtQ+Zhxg91b6/H8Vo7+/JEAPiK3/cuIrJaLbXTlf/BRJZYcH
h+reE+rZCdpS7Vle/T01o3VEoNlKH05jHlUnLQ0qHHr+o7WEy3uGJVREPlD9WT6w
20i0CBHCXkaifnDXbYhFcsIrmy0kb42Vjx9b5+cuw5JgAXHN+qJ0p/RkrFzt6nbX
+sZgNOWbv97fF1+fYj0A2CAtzkORw9dET4D3QujwIClUSi/UKRoNXQwUXOe7tq0n
90796RBtH0yymZPNzLCBTa4ZPuNApWfTdeivtx7fgAvNYAKZ4hJjuvddAInZvWi9
GsVKfgUEaYQrLrqraDfvwKB7JswRT7b3OMCO1gakJVs2Esy8KMW5rEMaEs5il2zF
Z/jdgazuTe9SUDiojQEHO8efSXZ9lhVevRtIcB2N0G1V6ate2ORLTpX20N/b9d2P
SIGMKC+EKNS2UcPjv4R7NkOQ42V19iO5JDMHltbEDMkuQ/Wb+JE3ic3LghXj723L
DKYKlTUk8Lg7UCMJyCiwyYGyyB+8f/HcKu3gbl0s/QcF6i4mtmMJLCfSdPwkxgb9
DW1ZUbSjwbtNA/mFkdNBjgrNCHutggK+GfWnfTo3/jwtQ2YJGKk3IHQ8ih8XiAwQ
H3EITFfmpJwHewXYdbNPpHnyVIdBOuG2fsoCcgTCpbvV0s+1JXkExhFbAC0xa3MN
5VAfcaRTzd7Wdj7pjxYyh18PXYsAXyR1xgOsuxeDCGwlYx8IX47VCb3q4Dwe0R0Q
0hYsKl902u8uWDRdoQ8j49JJFfzqyCBPzUJiRwQTbk7/yRViFtYhalGL5BKup+M+
XZJkvxdlrW6VP0mHdDcr4iuWyAX6tQ0Zc2QA6og6HyBoMufL2Vlfj+L2z1ZxOKwX
EjovrjsGpg8OUKBpaqVJrMVPw4ipIPnD3k7l4Tq/2Zizt+DhDeBCb2WSug7GY9Cs
1BxJuFuQ5aUQBp2Iwk/yT494CPQjsnxcnnzlS0M80/jbQaP6oa5o9BE4VjKWx0Uh
hTo1ehrpFdJlDX9qmnI37bNxnB7SYFm31ajJhVO6ak54VvlcfU1wR21LCGBUZGcV
x2I3gWsKaWRLPwDCyynque49UxvGgWrtuQjQ0ufhr0s8aTpDkgSK2mzRVNaSM1Am
CSZRmD+3+pTPSkp2Id3j6aLKJKwfqATwm64FxuHGvof2yud67SUYdm9YBOdpfvpy
x/tVL7ck/oAGPsPzxSHlRJNlUBXvw/8L4phR3h8Qf0HNfDsme8s4ajokduYxPK3G
DUKkahF5Y5YSAbjWRzzcisgiWqwo+ttsnvPAkeQXZftRkuuN3by07BGDJ30hQ7NP
6joEwUjl5DfAIP4BWnd83AYuFcInpt5zukNFR5N4nHT2tawV7ikbVZjaj13z/n0Y
8XCrK4yMTx2I2IXlvl6vNViHlX+wEvct4cz5OwOlpBOkQBVeH/jk5gqOSoNQqNIs
Wl/Mr3r8xU0olwoILAVOYliUrrZDhdqIEf2awaDXSjtuWCbBhUlkg/tDSmX6PBbC
n+cgFFQM+CCt/0Lxu1hPjxEnoQLaOrQy+59IVgZW4Ki5E3ePEpt2KxMCplE3OqBu
55PrjhrwWDEW9kQgEV0LYJiUXURS7FdP35p7SCfk9BySWrDWmwwPjOrK5QFC8kcd
jnQkpft1aaXLGfdglgctioFN7AIX/C3Pj//w5EUQvWanJXC8Lzt+7N5YaoRhUMtP
1GtrDCaYGxYbTJ/SSQt0uSpP3cKG35oq2qsGlu4uRZaiKyhPAtSU36AY0245376R
bJ2ojzDPfp6hxagIdpJrOlte4jhhpzfLuMnH76ssx8Q7N6OlV3WONQH5szndDyJg
0v7IlhTecu8re5WB8N4sKobfW5raoeVJg1KPa/rtCk9BymT1C+2x/aT5vlhFoSM/
E2arxqg9HxVP3kowsu9p4YWF8505Vwx+vH1j0uST0WvrIFRHjYYbTtG5ZdOhxDyr
S4wote18Jj1OiU8wAs5mjegfF++FU7yqDidO6zl4auMemkqK/DW8EEFyRJkT8JUV
ilZ+t+97Z73J93uE6DsIvOeU1UXNh3AVDJiQsIr2jGiQIdKckgSgpDgN0/WabHkn
qZCUskBzyxqS96faAxQuJTtaNfJFTddzhqF2YTo4VwG89b950X6cUkBwGNIj9Fj6
vi+gtcqG8JfJOSpXbroJz7TMZtOyLVRpcgjbdOMciAvykxuTNrxlJ6I3EVUSwfuZ
5vEV0Lov0lfR0gGk8iACVjLsZ6psPmMzKRrzCSc2X8yNQkgWcAbfWsmXQAFIjX4d
ShPBlkQfoDu9aPVK5cpN3PJ1z6p2bwXVpzgoLXHktawWNGw6139CG+/jOSnpTuJi
zEURtnBdraV5uNH7Uukfu9jp4Eu/DbWgMB6rJmWk7NHyzzwATCKXkYtJntGorXYX
WwDOZYup9lJ5Xuf8ZaZ+ZqDwmcTj91+Hku3XBtUsZUesorQ04UWpb2jq1JRl8Xld
tFlxpOdejgsjyhyhzH1s19reMv8mU5E5F9Wv6WtEpfNKPLPUrr6xB+svuKMRnjsF
6vavk2e44WRjGAWotpIYQ0OqJcZ+6n0EoYVYGQbTFSZ7WJM4Mk0k6WatpwrYOIQ9
cLUGWTa0VoCvCFcXCLikMiETABl0XBLmQVNXRwGKdP6INzMxFOpzVN934NSa6+rr
o3mj9bPpDGBfbXdznjM03d9huJq+f7vJoDcI/l2fEzPl7Iz1msca1uqULVEwbPo8
XhkJdnF2KrntxCMzjlnDiMEHIXfSpBskXz02odz8mEIErsATqP1/35ihB6UXWYSX
FISaFXl3XYCzPgrla991pDs8/1p+cm6oh4p3QwhhToajUAiZkrJHh2V+iI3LSWML
ksojQbdXS2xsR556qJUqjawh7jH7JryX7qissOfCyUte0R5WGQkxS/HeGBllvUnC
qx2TocNJeA4t8MT5oUYpfn2azyvfLatAMlIRFQL/VqTIdvavlvOPyjbameJTcym2
wCUCNIwZLTvpYH2Gvr8i5d50ta77YHVChSBiGbDTEJsCW3FA6FI3qC1le9I66f3s
aDbL6DyeaAJ2O0RPoJQZfEETY0z0VKOMgWxA/knIWGMJW/qzs8UDOVZbY9yngXvW
lFaHLln9kauy6PMOjwAeFJyqGd7asixFH42o3CdcJR/UENKw7QjJZ5hiB6f6uFmh
yhWnXkQFMdz5vb71OzEGRNrCzYchEFrgpPoQWdjBAHZcywIxwYsRcWcbn6UttTOs
bdk8Rt7nvQHty1OHkaJfHe8a1QFGFxruncVKDu4zSptT3Jl07q47Qp8I+2GIhIQI
SOVDcIwd9QdnOfLh+EC/jXreePFxfjiHPAquyEgGuZkZ3+f62RWU9n8rLEqqeuxd
lSxqgICf5L2o7YtpDNPdhKMdzCFGu1b/SF3X+pGil3o9e6VLSVJVv5Z0KN6OzUlA
n2ubUsesG8KLoZx0XI6J28sYUf2jA7Q0GCPBX64jVMy3sbP/uKTuDNCl6ZXRZBBr
7TNujcbbWQiGnQLahh6KeFrFBLGiEq3Ko1PGP3fqgQefEazioxxLTIiCQiTxyxcc
RMPeiAsQBW4KHsTCU7hI5DaALoRtiDtUNQ3aL+6bgRsXzKpoutsiTnVIxShWyuFt
n2wI/ui/mcgHa891ek0iPDSABxnFlPB0Y3xQpw0RviqwgisyRj4w1gGA6p/VRrAp
tKCtds2Am4stLdpfBcjKsA+yodAiuHxlvisC5bSqu3T/ijCLm7fkUJZYZ3/nolnm
OMoUj632+UzaiySIQbgzZ6jLyNWbTB8463zmdJSYzjR7XFGTvLAz3t+8cKJ/aI+p
zH69g+oxE4XrUm+bdY4ITsSyIQc9qvzTSH8mjIPxK+yLiKic7PrkIih3pH8WmX/p
RxSqSiiuP6y98eizNEPrWgIVtSOq3vVS8M14vN6+NxAzes6YArcI1e8XghWB3jY1
mCXq6dqgdZNSC2lOtgzUiIBlso+laKZgvyOcX37XHgHYW4O2IUgiY6rJQl6CIqSK
3L+x7KPiORDilzsa250m1PMi/v7pQGCIBMrJ+tizNwGc5s7wG8R28LwAlOZZNtYK
z1AtmzHTyfkfoharJ4NhqONY5NfbEgHA5yNX7/QE0yzR4IfDlZ4VVFShvJiFhSd4
KRGpGA3AijKeTYEzsh7RQeIjWc0+uqmJn+mwHM3dc2cMLjjZq3dND22yqIpELPEQ
g3wDLVZf1hgZQCD+R0GkjY0z4aKsQ2oyncyvgC4jZgtZY1f724IrK6yQbhazjTOi
YS+n/ulehIfFupylsf3ek9Je7f8YtwAQQvTqe2oUNQftbrXFYMZGP0717Ax/Aal8
JgcntyHAe946oHL4Xo4rc9LcS/5y4OohB6DV78QX/kqJpUkDBy/r/ERPxm9+lm+A
0rdP/bLJVIPmAtbKz9GNwYTcO+LJ0cSEEjT7hunHKAtLy8nIGTkX9MvdBprxjICg
wBQQRWKz8KeKSUsrvQsjUXCt1GtUe5dS+iBls84AGU1ydRpPUDNexIpKHOwD2w5/
qBmHMAG5Rej79LtNNt9IjpgIXmsDDHKvUb32JwU/pp9/d9b8Wx1LvSRfMLCovLvu
SpJl9WlVJERGDyzo96MmE4L2upOawKiogEuFgBPlj/xiJEZJ9yaTelClli3wX1mb
oXhNIxZjsdtM78ULsqhQKG5E9IiM2LLMAxYSe2r1hX/PNatwDvSFaMK1CY99QcMU
5RCTCr9LlrFnlsYN9d2irOzpybyvxRovU8agLTbREVi1s9QBq0SYTKdyNwI8uzD+
P5UscZ1kSp2NInjJCbt76+WCd3jgBf8gePgWpDR2Vq9j4RgrGFtywL/Fi+Gyn0iQ
ou0UTbCwZ/iV2FLeFqRI36LtFdr5Lez6FFeh+NEoDZRtgmH8etDUhWD79JUB+xn8
avOJ9HzlywHyHs8gTKYn8BKmPW4PQqW7G9bwYPABuO4bw2d0JdL0y4QX1TgKHqaU
/CHwV5/9Po2y2UiOsGCHb084V9+NIS5/ejmsgIGjws7+nExrmmgmEelLX8sgfq0K
IQfGBiz6lW4ddupubKZv2mZc1TU2xdnNLX+J/bOTxiIA7e5WD1UnRJVYikQQ91TG
yXprqQ50WvsNYH2oLv3y/175owmYbO15ISNMUqYQokx3hmhFX40Xgrf07+QcMe8N
+n4cE7qI/r8vBQF44nlGeKMIN4cCuyRJhF0HPLUccGr8sF/oLusyHQRh1MAMH8AP
SnSI9hAaT/UC6yxNHqQz3GK3aovmrkKAxLFVxt9Id8f23aOw1Dj1JOfT/IB0YtiV
Lidz8W1YKEmywZly94JU48rOQNlj0E9CJi071ZgvZ+kujX4WajJ2yukZDV9DHFFM
VjxXFxldt8+oBXYFJKA5JH5S7J6rIap8lRXhWmP6T4KE0FaKRfY4Ei6pbjbb61MK
3nTNyfsibF/tJtuqJUQN4OTQACRrL/mMydLuGhzOPyaZN2Xn21Qt11qTJGHUtrX1
bpl138amjPY1t5ozCNjmf0zWtVrEP544uNYKNDCh1e1cNXNcKC8RF955vVl1C0AD
QYLw3cCHMRnCLFkzBL7YEhnSx+b1A80eayr9wIfZrE3s/NVROgCJDLKDlpRg8kjV
yp6ZnrxAmmFYDhDv/Hzosr/L0HNw2AqbfsPz7KYYgyNWssXdGrGo6wp/hB7TzhjM
dELfgsYuVDVcBZLQ7T7eQw4fkm0Jf8eVnLqnppw2Jb7T1phyVTxL668a7eV88zEc
l5gTGxGizCMviH4KuSUbpuAw2thP0T17bED+8Arx+p4MAluhfEno6m2bafOPBLh7
U4THStgJb5U/zS9U6QAnUPbq+v4pNyfHbCjc/Alz9A3H1dOREPT+K0/CF6jqbhDG
AwiDYm9Txbb6GQFXBxokSyaoC0p/Pqc2otwl3g+eUeFWMTpfssq50HbSRYcrdOIX
miyVY30lmCnLBr803fXUUlYOlO86aXYMba5HPWj+7gCdHbeIbaQ7tHmU/82Y+svE
y9/leuC+t6Ado/c9VZrUkN2L4+30k8pGwW5a7RJW7/2EAo4LHfUx878KKfAjocMw
CieRPUJ8eGR3krRSFpNYIzcCjg5qFR4fru2gvXN2Wqt/uxE/R7U1/bBmRMZeJkX3
8VqTcprl4YgfkldlqFlD5vR0OaBxP5jiWuU8SR8Pqpj8JNiUGZmRAaw1B6WcRyW6
Ah/dyAhYIrcbII4inIwyOf8BN9Dk9/fG6K5A7In168YThKDh/P51CKH6a1RwdlKk
IOMBRnJZRTXMRij7DdxVgCAaaIUk/4t02UM5G59Iaq1C+3OPojW41HxilZLM0rdp
BSnY9z1ZGichDE4WJbZuA+t4aIqEQoBU96cnJsznfBuYu6oS2ZAeTedyIA1t/WVQ
Xqls8rvxuYtms8P3WS1PTdbsyQn3W8lUHb/oFuPrZhST6icfHs2GWhiy3+2f1cU1
IywXgwq1QFnxppQ9OJq0H+AZEJW89AKANI8TJUeO+NbOQozSWYmiilAHUiESW9tr
T5G0gScLLawhAoLjAAJPvdyMKpxVyJazNfq7xv6W4DsZjuLgbIsWztuczBcl2xWc
db4z7hoJbY7Nc6aJpwJDsGXOmerfblVGHyq7eC1dDd7jrVCA1Yg2MNRGKsIy/68/
BpXXsmCPh5JeL+eJ72TndyTcFTE1qqGSNX9on3C+k06hmfqd2scBmh8EODu0pApH
yMr9vZnAoz1gQTYdU9I8LF78MW/h3x/rt9ve9bZM7Fruef5H5TfQ7ea72YtYB9qt
QyG39jrsFRcpv45jssoOY+BtFfIpUy37EDzLoRniRx8XS+uT9r5OK2O3FihphE8s
hAwSTVVeGiHn1e6Ix4YEDWSAG358gakJiafWPayVMyr3vDlah3VDfF2wqHLnswZY
FSkO6Lfdt7GIvB0s+UAzqClFr9U+TCO0kQOqFd+2wAeZ4VQC1KWx6jpf3bdnyB1a
T33iTb6twxtxCuKJ9iVq1jwj9ZoEjY34K850cLHNRMN6JILQanM6JrpEJRrmSBXc
oGgLqLfop3d67iWQYT1yNTEPG8pw6LiWPZj04siF99MgAySPPBJfC9JVv1C3UOvc
lxkaC0em/5LARZ/cUEBp0rWOd1oIHJH59/kba46Ha6EHOdtwrcgO8tpcRJB9OJid
xnZwekBRxT1EMgtID9bxC3egHQMdPxmXsY3UV0/OacYIckCIz8DmbjzfZYkTQyHS
XrUt4Tc9PTzH25QipvPg3/xIKNZRhDIcZlD+7tMiaExDG69N6cSnZeMnGQft5lND
alFpjkzTaCZcWxOE7Q+5jBMOMYw/JEIWvNFAIyzJIOIFV2HBw/dOIcMaYWBi7GVD
ke06JWvxl6ssljoFR0QNuNUKrPXwV2J679E03xvLyN41t+9s8aD+reu0o/91Xn4a
qecgcOwnhpeGCBJtjAOBBZPybOJnGUBuskeuoCl8Ttm+j+OImT57ran3Fs7coqtv
cfqxZRTuE0ZjdV/MKmOjSzbSZvdoOX9Pv0S9NPq0irCQkfVeWSeFLnCc7BWHgVJU
gfxlBod5RUAe9tvFCKPF5MuTBuOZTJ8/L4BvuVLCHLaQt5BSYiMoyQKGQBOU8+3l
oRPOghKGxDaxxf4l5o4eMrEZFTr/P7Z/l29p3ASRsWAYG37PpnyOutd1IEIoy5DA
YfqjIspmZUZw3UW8eKqyyZhEnL7zNsqyU4Ulyqj2t2g40/t0voXVJQBGUv06K4Rd
wHpc/oQdG1ivCbowOMPyHqwn+sDsv8nXfrKzeCBMbQQhv8vTS0AGPPvs+2gZpont
IrHFTCUa+AHbBua+6qKCEUGpw+JECGfSBEe1uDC9c3s5VQRM7CwwHVr1Y9jURq9X
tKIm6KgkrEhvFimOIArBnMVj3HiC/ymS6JUpLndk/0zzF6sMikMPtjoaQdy031BY
7BR4FcBNOoQSr7mkcJ61qAJ75GeFE0Mx1EDgMm5WbTCsM3jjT1r1FDMn8hSdgADk
pmuFc2XGfn+COtvAYVqRlMhKGE9cMP8ndjPfQ3pZbRiMbdtosc+Xfr1nldaf/H+p
FQ43yi2hBN8F4LSU8qaMLGBqoVu4t6wpxdZJQ97BDRTM3xafYXxtCp7sNeA0J+tX
pIlsw9aJjcXMPfv3LeEBCl8wqzaugvIZYtw9x9uGQ8yfXo7xJPZdML/KuDP0sAHd
ApgfxY+Om6hJ+nuLTouBwo7zgrzS95xEo7w4QGqACQ+x3kJ5wjiS09tdeuEJAWDr
0uHLqUtCW+55ZVEpy9QGn/6jCzQA4rQVgHWQfPKsxMx8+BgBGJbtrqp6jL//2d6M
IRlWXpYV/tWQydFn/kZvQc5Uf8DViCOkep45q9tCbe9uQeIqmg9iZZcdYj4ep/G8
beswA+8WkYhr6nVczSpNURiUXsRIVRIJcOp2oqvQ+kcvhHtF6KrExCClZVMkErSB
5+IX3QSNX2v40ZOc/up0ZcNOG56dwRlcqPCCoFkDTaa+j6OFGag5grXOvNjFlLh8
oKwQsoSiJFXmk5DKGsKOwhXr2ilxqWghuGHLTjNgSI9l7Lx/XNmKxa5+t+uAkm1p
HFq6JxPgrjR7dLML7iIvSmcQjyEks/6fvPtiAmsczOwDQur/9n2mIa3aII0u6/Ys
dliHMd9WxtH2tOpIPxhAfWoKi4gJs+bt1GZOa8LFarxxlHz1D8hAWCjh3Rx4gj70
BSsSWXWESDRJpqSJtKuyt4tlPkBEZXU/+myiAzw64h4yr/pNNW2mA8V3MNsjbC0H
d4xEklp7rBlRAjBxcZ2CZZFpKHdxZzh9BPSk+pk1qZOPEDux1KlDKQzi0vE6SFDz
L9fdI2G0eHr2XXowNX5MLHI6ahT5mAwrHvmTb3TKKzWClnS39u6H8UMEd80NJUZt
c1svM0UlcS9P8UlmiMFg0MDcNx423HXgiP5G5mxZ/vQ6+gEBZ86OsET8Au0DX95P
VMNU8pC0jSTgZBkB+Qb96n5A0RiNIUnCy7w63SgLP8PUz+nnyn9Rb0GqN96+lt0n
5yEl2Y8C+l60E6fkJ73MAyJTZGVWimWMwpKx079oz9Mld+0u/j1XHE75vWk/MYnX
MxziCIOF5xmkG762ACE31SUfp5s58m/vcFEEdhR8JCC6ZJGcaE9ubNw0OJmTX/yh
mNqvZ5SbcPcxh56RBkQhxj2uS3Y2E73izvqB0pCpUlO4qtWbLyWNpWlDyxtf0+UD
/hYA8leYDh3LJci1WZ8OQ7KXkRRYnMMGf/b6iY5YR4EURekyJdaEBElZcczBccyH
S+pihIx2nfsk2IrYhtDpmqpuP3clBm5g0Yr5LCVcd8HGITEmgIsxaOv7mtvsDUpY
fSy9u+9sE/suZPj2nrqKNt++mAmVqkId55nQ/AuRppJmO4orrh2E+I5nff+qsPEO
OreLZYsrS3+RpXzzDZa0vjablsGIOGvOKpAih6Mf2S9NN13TXP49w2ytHD9VzeR7
Qmw0N9uix/x9tyvZNoRtv4ZVxyIObCuK9y1MaSDo2j5KJFw9MXe6oA3U2o0crZ6B
72hlLFUpcqe8YUfIoVphTJgb7XUW1aQOfQKnbU72WiWeMOjTw9nL9UvPoW5Xr5WW
8rbKz5a4c3uNoTFG/NNQfqLyquwk7J1lxs2mFLZspaUAgDX+TFVHM0ivimEpWZYA
ufGpr79Ca/z4+sOrJYnR2DSL0pj/H5Re/o2kGiPI1AGfqjxt3KTantNbBEGLublp
nuYkv6EmMu4kD/NF6ry0UhvoMG/bOb91V5kVNp2J/Nfgq8cD4DGz4xQ72VQJc7ev
G5kvR8pAxX5UnLZDKA6zKObFKMSPx9zWLoEjECf1E9oQzrpKskSO5I7x+tG1FZ3c
gksVnyP5ADTG0fNDAraA9pqQ0zCJ+G18FV8GmWOyoZF8p5WPDQvMC/H9ji/g6d2G
SlwPkH+Yp/lThmUUMf3y72iaOC2I8wnnJT3Ick2JuSyg5haItR/r8v68vmO55ZDX
mE720uXy5wlxfNUAIkmZzLj/FmDNEoTGubExJxfOvebKF9bYaOfZ/z5RbLme59xt
CmKVZmxSWGJg7dcWsIJTCYB3z9gO5SKM1GGOCVyrBT4sWAh7CoEOyhnTQdOdzwWw
ROagvGzmTEGyJBz8wjWf2v1ZMGf4IvlIJyme2fliFN82FvKMPzjSmi5HPGgKqzWW
1n3g68TOhvph8LxMDopka1AiIdTNb765D1ytmHh71EnOWgDnetHAYJGzYeASj+F6
dQv+s3anOROaSA7djMbidVXrZgsrLCQZQpHCUpVt6XVGAjYKisAcDWq6SlocKoQD
ecAfVkL8FUh+9yKrSwB+nEMB0gTVcH6PXtgt1en/NDWNNfFTZygkvT3oaArG31TN
VvTgGyL03z7gOLWpWVqPtRCglSo75bUErbKhUZ/9AsbvZnazwCOmLphFa+tG7SWe
fSlg3u7vq2ZPlKLA2syWQOZr++Zvfi8HTQvVqKlcNWqSJCRaXoWpNFmRZ/Ot6Vy4
YybrYLD9PboSloarJAoEKadueJbQBPzSK4tlPEB2qdZqtg3Ox7zH/GdjHuRJ1WUs
ysOwbHU6U05RfkhWTsxCJ8BayWuZ/v2Q3cb3zjys2nYeYeXz9fEQuxFYQq3/nLBj
vyGzUrFmNDC7XhXxunqEMpBYKzs4gBEEBG+9gCELs2fsbBRxXDryE/AaSfZYTDOl
D61iN+8bu6i+nCa7BRnVP2wvRoNoFKFdeCwTMqMX1bOH0RrELfOa3FxeYvaMwsjy
rvBouIR8SMK+dsatyrN5n9WyicutX4zSCC1kk/spv7GDc7d8CGvzTGbVFcI8F0Hj
5W886eSf4EQ3+mmovX4E5wPtZvqBsgbrSAf2J8IJWw6SSgFbT3bOCVH4ZHt7/b86
hQKAGhOip3mg9Zy2oCeioFWG1NY5O5L5Co6eIwT+WCEwGvRUpXZBfEoKRskivjbQ
rwqfxfe53l5jXLznMzEEGkwxRg4WPooZZlz2J5zOINjOhU0ZU7r35f5y9nXGq91k
hBmvUzI5loFquD3W9qYWYmFu7HzLeTGeoj9IzexJtRZZVTlEBg6wXIbmKE5Nfk5B
iGG7kZuwi1xwSKKbw03ND4cFk13Gp2pTM9x2AqgQMfh3FOMCCFnFUHkgi/SI5yQy
i4VgYfjWQO9b94V6tWSIl9sMMPTz+0eIgmcTSTOf2pKzP6YA6l6Os0TPwRtIWT10
fzPaLmyWswOf0irfdMCm1apDE90dTaS7F2NAp6QIZ/EABdjnYTpvoLt5/KWUFGYn
BSYTROAKoBmsWoJBDOwBleoMgGxc7S5u5yJI4q7li20JMkpDTHHaUxFoWCHd2L71
l+k+Ro7vThPutQGg+52s6wt5/4NYyBrpQPOW3OLnnwqfm+Kxj0ewt/fpq8V7HqiJ
KzsO1XkwAiJrSM6zgp+ssemWkNaEZ5uTRfnOvE9WWjcDezYwQlqlAVDsB+3TYAOP
+qtlKmzerQOm7YyAqht8ZmUsshtocD2+iXxc1ZZIhq2ditFyLMRcZgoM1W9M6pyV
QIYL45QFba8EiOPt8Pyxv8sGNZDNOcp+GVSbb1t3ca/THuBiNH96ddj24ZaOhJ3b
j+WogoY8Xn+MRJv0wdcrVXMwgd1F/MIeHcqkPOZy4vHyX418SqWMKEddLu8czCQo
1pAQI7tcf3iPifkV/fWKeG8Ycincw5zAY2K+Jo+bO8F3RjutGUeDS19J0X3A2aNa
f0b16b9gdSS1B1J/Y4106STErB70opcCz2uNdummxT2F/CieLXTSMCOzl/HE7u3x
L1iLhDOESWfNb80Cd+d8cnFytiwuFh8GYByvOJ96jpdhqoFPFCiZdBURaT7rJect
U+OcZ6rO3bsevDXChg7lr14vgaYIP33faEerM1QzsUptAfQQx73BUjs1LXyMKMaY
IOGgeOrMr5ZifzKQZzAwnVIt/aLhF8X8H8FthjX9fVvNev9vSlb/bL8A22AYW4UG
cW4cwwhvagFORoZImG3aQ3M8B+cWrWflKxVYq4CcumTN1jKDEdhl71DyV31KeVC+
ISNYg2JqZb+u98FOIqdQhltvVMWj8ZR4f6zkv3gfCemWDniLX7Eig+xFMntPivN+
W1HJ4akBE9EfC7j4Fhzithz8fNiMjEXmEF27HZdHeHLPpJ+y8qy4PjJ8iTUo99cW
+0MJTA8BoK29q+sgQpwtzoje9JgRyoWeyeXTQ6+wTFljCdur2YaM1WP9oZnE++nX
3aJSHkPhMvSc7Fzn2pypV7Mh77rAlYti/lYmc1I2/wbn0gLNcF6c0bH+PrOPcQ9Y
EKVluXhCL0q9pLv3iyntJS9TVrzHjeqZwmdo+Nnmn7S6NqMHdHwGae2HpeRMw9/h
r+SyqLZSkj5MsxZeMdrbmg2JoUCsuD/S/uCWjYLUNFd/Hc9yPS0ZvuORFuUbY7fQ
cLIKByiwpt6XOe4NeTnvCLd0BYsGzs4tqPGAJb5HqBfiubGv11BsgZ8JCyjTE/Wm
sZh9U1Q5g7NA9Wh6bnAh0Ap3P0Y5dojkTXTFHYtek9sAWhABCwrGJeldeBna4J0N
9QpSGq1F05NPe8aeMaEDUW8iyPo2PLKzMCxRJman+f9ujDHGwM+RGw7ALA8bKBOt
Reqie6jBNod1BFYh3j37NV8Kgvz5vEVxiB7a1FvDl1aZ/NWlDrJ+h6taF6Bmq1ep
SSTyGrAJQDPWGk2U4i8Q0KTjiR43XNkgwcsgjnIyHt6hn6rtUe1atx/gLl2+JILc
dn1NZtc1abcrMb/bcfe1JJRBYCFi/ptz5j6q7YCjxn+XD6pWa3CgwwNYqxn8mroj
id/Q1pCPwGFmoVUhKdBK+24jjg0DsE5ZMs35pibX+SiyMPTIO6v/b5j+OGfybLNR
DoP6HOWmw/KHz9+QShmU7llc0JlYEyNaopmi0Sn4bhakxuYLMRUqajKHnFRMDfZ0
7gO5xN2acKnjR4OcMELa1gOQL/D6A61kvPlOtll2V+M5DVNa3q8/Cm4Vn+rMJ2zg
n4LN6BweLST0BNOKMDCFQt21OzJh2HG7QeIUBjCcWZmJkU6DXZVEiNMZAjbIRSCl
PzsUt4m/ULLI+C0yXHKfdP0da/JYfE8skW/tsQvA3ehxx7wfi6EQQQcNahj7XsD5
37ppQhFBIe1Uo+S3HkevJxA0LTzaiVjxc6hXkJ0lM8HugXesQHawU6BOe2Ab/Eg8
c6ir26eeCENHa3hJa08Lr/WrKGtp/rNnYd1a6YnV9BwjOr5gNtgGZb4IgkMIoixV
zNBAySy38z4qRJ3ioy4k5f5nMF1Sl25NHBk1DiVoReY18jRqcLxhXPp87wR6fTjN
6ftyA8A7ep7IMpk2yzVcu5odQONChA9Ply0LBys8mrDoFKWruqsN6dYbkpzavuqM
u8HIwbNgfsAFeybhH3Ccep5OpvDnXfsc3L3OlS87cJuuww1qF7NAMR5IvINJJLFm
il+N5t4zRcicktyipJTWnGggHndAXSlsq/oe4tuqk3+VaaKJLxzRaCwcyT2gE3fr
j027Jn7zLumtwj+d+zFNJLGROMletAQSVA3ELWjTcwUfaAdqB87TaJvtUVdT4PJs
ypELMe59JjbjxsVzG/rzwLrQh0FWHJZqrm4ogmRbaPC+gJ/Hkp5K5uAUKVXJlakk
D9k4vf9wcOswo1Aa1vM3Wg9gIi+7EFyruhQf9m9JAYz349ZG2nlmLlWprc2ECf2o
bqOPqwur7fHiytucv02a92e5fe8cuwaa+067zO4SskbKbMBp1VguO2hVGnHStHma
/LUtRrSuGVL6SojsP6v91mLH1dKJr/KhGZpeKSNV3RBPkf7T1foPRA8ao45WoMWc
RvgcTuFAwupBQBmnHqsrvTF3kfQkOPVWADH/hcDSAFdUQmPRifr390WgxSib7WNg
qD1Rfleqr0v32LAWKY2ODYcjHVU6aB4pOSqgT0hO8OjDgmi9WDmtZKVAFDXo9Xv0
SAT46FBDbcbCBwjSjS/Kmzal0Th6tC/bWruLLmUtg/blt80coY+lDfCzE565DvSn
bit48IL5kMUBVeRUTp4SEI0u+HMM6EDvrBaz04tezC0G8f8B8ibJWRN+MV4DZXtx
gikbQhCM2RVoU+oNAQhlFVlfXvtFY88zbVf9z0FQB5kYvGdc4dYypM4N9Okn6q7d
GQ+AINvMHkJrWiknwqcFZLF5+u2iLmraz1l0o3J27ysdwdlpoKAWPJQSUS29SX6k
wT6QRFUbE7awp+GJaigex/c/Ry96EhY/00o+MNgpNo91iRUXStTBdLb9n8aE1GZG
2dBCfKlKUonSc24+hnGjPnbPFy+D5LmutshUksKYIKHJ/nu/DZerZjed2J+nRlpc
6CQBLlMsn8OBqSlbklkQz1xBxZ6VZtFnv5wNCM+o5TO+VGSQZoiTIzmNnUg6K3JE
WB6HzQhdNjwtVWVdaxt9JHkWZ7g+lUPC5qOS0j1yvQ+GtkEvABHyGaPa3kyEfYYd
UlD3+6SWZxdtOKOKSD3mZwoHL7ctzfcgRL0sG512P4fPSnHcby6++Lx9FntihOuf
JgXN6RLRvwl7ifDqCYP7Cvmmre/+TpsTqSpbr9jOi4DvKMN6B+PTimS8Xkj/KNOO
U8uVwPE0Glv4k7fz+Afmq4f56i37MF5tG6El3+QOaSnBu9GRTDNdL9j4NgphOT5j
tu434tsR8twyiEmMos+CKjH6INZ9slb+RcJB6DHylpvEcso6q3W4zojn4s07kJui
jsFZEqaOqFCThbK8n508kv8PeQ+tNp2ULJ+2RJ1GqF/9E+UntV9dFfkJ81Zx1b+y
ytrioI+VjzPUIfgKkeyNcz9im+kCHtoWlu8I8JaVgbs8e9OIFKxxYTlu0ifNodYw
6LDmVpc+0sz68YBB66AsEUC0HKRCK+4mFHFiJq3sLbv+Y1wiS0OL3lwY7XfQZBfR
RDTtFawEHgHr5SLb1mhE9cLpYQZqeGyyULeEVd1gkyWZXIJ0ovfgWOaiUDuVjHsB
bbdDq2cheYodVn+aw6G3MZNIE+HGpsfsqvaXW8a++f5vyPGTnUNArWOzNy4WYRk8
EUjIt61MXiP94RvfjHsmNFRMQatbzRDq2LvEQHFLH9JRgL9hwXdGHx+AMQthKiQ+
+oEz3arhEiWZyq7tn9oPibxlB9sOpP+dy56hM3qOrmSe/iCg/sf7ZgDiDzPy4sIW
39B66XmQluHW2Nq3b/Lk4avHKxAimtEsnRFdr1GQwU+q2A8dsBr0eugYop5grg2q
W0gfMrzyWT9ueaMnOb+SWSneUuTDO8ID3tQPo97nPm2Fb3n/7pTd5rjFGhOQkc12
00iyFPbok2EgoZdlTHW6sTqRMdsM2y99Zz8WtrNsvkLg5clU3VQ48kgUqFS6I1d9
2WcBLIpiFF2GbzahaiKLG0xKOEkr0LApMx9NS+CqlFHfU1dLoVT6ehb4qWu3mm+i
ZDRpvgVBD60HCtwWvvWT0qeZH3s7nGsjoKaaOyWcuqfrEbdOkifR8ECvshiSfIsi
xNaRPwDrKpsA/zY/+UirolYPetax4Cjrw0y7iZDk/iGkzzUG/WzDcPoO2Cq/6QcS
JcNIlb3VmWuRV2biNa/K20w+9/lim4QM7BL+Y0tqtnsYack2dvwyoZRirsnjEXY6
W/0JnKRR2VndB0gC3R8cm5FMIdxLhTDyBc62W6OcNVcsY9ct1aUT57jng3OEMR/A
s8nGFNJka3xD6qdpTa4s07nVjrXFB/GrSVmOaiEFZEXbyJJU7C+lyQgmeanegxNO
eyiAjc9c4cQDStUUPiaHULB1o2OBUMhjf603sZNh+hr8ikQYJCWdR8USI4oyz822
IwS149cpEvuiypwCgXrlC03tYtZeh4J2qNQzFAq9olDuxrzSadrtdKhqXbLwcnlR
0ALX5SZWRO6ABCYlLDtKe6UVa9ah4AZCokbK9eA9bG12/3gqM6ngUn9trv5Yf1+8
60LPx7bslJJckoynxwXGWG78ysvY/tHawJau46VGfRpQcgbUVM/NYPWNoaoQcykP
MAD59wuJ1yK1vJEk6hMmUuZBinsxJynwy+EqRPMFeAGh1L2dfxrbfHd5AHcMG70a
+HvpAmPgpg30ICyLyYX8Wnn5+zdQxN86c0lHkv6pCG0xEGeeSV7TKWLBvMmeGj9d
EzJXDRILw0XNps5lkRGCh10i4GxjuIpeCUZNYyAavcYN9eXWrwmHoG5m3AFpH0rH
bLZF2X+V3TWYke3JmIZOTEutWvzgwYn858mXWew62tBEEbGyNa3Fb056spgY7XiM
iA161y6JCMIlDrjf6oq2DIOvwso+zWH/xqtDULkP1AKPETgVEfkU8upThCYhSQRs
jcHYhBRLvV8UBY+LURnHKnqAzwuDxqqO120c3LhS+om1uFQDh11PCd9M+KOUuIKc
vYFBBynOvOAtz48jmCoZtNkkyRcRCkqoFB2kl1PNUuYrZpo3tnaSsENohu4XdHVH
4ZlwSmYhIWRsvxR0Ao+nA6SqF6UAFf63B0wxPGrl15ExMOTCvPJoRmpURHw8DxwR
IzyPDAGqwiFPiN3b26RwI0B6MDzVx3Brr0TDNskycuYJmxnDO2ZOg4PMJT/LFfwZ
8mf4ajMLutb2A6S9M4JMwW8B8WrWTMwE3Wy8sYqreJXHOb59A0x5g6uVIr5cIfxX
Ghcjz0v7HmzLxSExr1eim1x2EFWaZ2rdx4qe4+0etmMvAuCjZfjX34UaHdaHN5BB
/LaJKwWkidJsJeaZAvkmTI8EdGwXGP/APSMSmXJSef+ZHqhVsBBTKTfQUibyYPHu
ToumHjm8EqvN+dQ5DRal1mMZWnFL/J/T+DhZ6tW3vvcyPLEcSZQYhiqvqA5n5deI
sJMm38OFhzJcQXkOGGo02JhxxtupRGB26/MZoygjDok0JLWuzY3rFzui8RsOCZ/X
zDFwnT1dL5sa/LfINaPQbIIulk9FRBS2ndx/qXj14ETAPPMySrS9R30wpVfT8HuI
M0nQAj/sDugj/DIi6iHigJxucCUrjiZeBBAThSk1lQjwzpkM8L04kjlH1ePuKL6Y
IhJEEx8cNmOmovR5+Ip8WFXRzIWn6SHap7tkPbiimmbY9tXw8ht2eQUlJdszuxSQ
JO0nIG3gXhV7tLMNk1ukqNLDVtb1+cTluh4EyJj/sbtCCSaDRvrw1+VCxxy3jlfD
C0CpFTWV9F9IDAt6RphR9nNhUQIpysSL0hkr9mRskXLUl4Kt8BCDSdEClC2iduYo
V0yMIm+yvNhwmOeaBYrfbbal0Mgu+SW2OWlza2gFMHRZltvbwvbIQJFS/D4XPqwu
Tk8TccvS2KQzSzlpt1O9N3w+BODB4WVSHqOKnJVlPBenOOrZ/SxGJmmexHGYasOu
fEl9agqUl7AvQQy0SO5Lew55n7jxCcSOwof06ZnZhyys2JI/aBnnzoKFkdfY1cDH
5cREucMiCLgU73VM0juC+r0xV0NgTe5igwTkLT3eRQJQbsLnOKiLWDgLUiq18CH6
3sBsCKCZ5ETgBDqXVTsMqIS6RIc05eN+qXqy4ikN6fkFYeBp6FN0MSAI1eFq9tyh
+WzwDsiBDSSsFHfw6x3isQxu/m2YjBYEqygVrT3sjp8W+BQIbbQB6ljouYXRgMJL
V6ZUX5yGZJYAhsaDbaqIiLpfs4BMzglSIByWvmDpxLRXofR88NLnMH9nEkhontps
UNFhkgjtehM4mFs2waQGN7Fgjf15RQDzReQI79Ey8qtt/KFKConBhrgu4T3zUgH4
it4AhxO335qBXpW9FITrMoHi1TK/XSzoJZ2VqbvKrA3PVHQBAXvTcHNTJciou5Tt
Pc6yq2DXkG2coRd0yJqhe92cfhTiWaJiWPEFWyOT6SDIjVQ6PtTFXtPUcGVmFcod
6UuevpME3tM/XMFmOJ26toDnvWN101mtC/mvC6NJ9rJmREDwhqRsQCu9dK+KczI0
jUMBiujP5lq1dl57Mkx/73wOj01e/W6CRqXZ7uJSvFcPgjM55wP9h+535i3Uphdk
cYiq7y4CLshw8pjxiURwiL2Zu3d1KBilBJozYad4fEGCfIg9psXgz63W2541qfzU
kX9xJiSpjs9MD76dqT2WPJaSRLN/sUD0b68iOVo9rSs6s/QUyaVwQ23RWamDorBo
XjmhwiAMoI8CoLi1MNFkr1+j6FmLuoHduFkMl4pmMPJXDSVZxw8Fj2Pgh5OJ3zAd
JaM/HCQMd6VxoKZsYiT3iRyYxTMmc6QXyipGa4wZ6gM4HpFKY8NfPAfqLI0rJ1MA
nSPbqwNi/g09HQSwJILECLAnPj5AqVHVggdQCzeOocqg9Ak8RyYvHebbNohMyGWn
0wScRT0ZXeaUX/rMeuLgoL5Xqo1vyBmB129/SWHceoj6Gi54HhvMgQKkaaazxixK
BpzbyN/pZSGU7BBf6kL2iIGlmA6AJtuwhcHEm87y26lF5VIAazwluaIIM0TD46yh
MzQJb0gnNkmX+61xn569iMKJvdVi61v9LUHFNZuh/tUDeoiet4WBFTG4OcPWzaKn
oirHroqVhR/YZDXjw5FyFYTsHTW/aYRyjLlOKDlrClEA26txSz4RPD5yTQh4EgsA
IqyyFkajdvrC+nyPgJD2RCG2QIyAsr7a1BRyIQW/ZspJQfsTFjWlzvZ7LsLtLJbw
IQoReNgyTMAVNBbwesFf8gx9iRrLvuIK5TF84/sNaC7IX9CWhhtfICtiPLGapoZ0
qcQvyDFUsmw0JjflCBR93nUwgBGukBqehLZhvD+wCxw89aIHTfaMY1AFn2TCLWDH
FY/28WRNeKFGY08tukIv4LQsSm1lWKagq8OwOP2CWKj5laIlXRJlkyz9139xFAf0
xZplgM+os8ZAHkm9wD4DqMmjRWRr2kD4ueZX72cQ+r1W435x2/r+8AJrCyUEke2a
0H1xbJo0KY7duKn/wuYcxmS9IX3pdkCt1YbMX+BnVqOPh65qPZ/SVQsygkm4za1t
kxVz2oRgz/H8aO9c/PKfoz7cDhVA/X8DsS8oag/mZZZ3fuzOQ/oX7hVfZxNrW+cw
ZyhVt0cTT3v+rGo+fq28DK7ojGeNMltbOefQ++sI71TWiIIcnuO/adBDLEHf6jD4
ZHzcS+5kM8SpIMVHfnPBOis1wGNj4N77RzFJizlkBkHd1WlCwUld0VlqUlRgChJT
POangqIUBffwZTCymKJwlSiqKeorgXCL1HGtMOkfXslXOY6WF7pC9K/ne49ql+z7
ZYKCLdP5s76nTbrcftvmndxc4OE71ro/RZOAsXjrMUsHDuoCTUmD/z0tpXk4N2QU
W5vtjgSUVaqJyXTXv8zGtX6UOMJxVi7GEZmoIuZ7hCFUvo3qh5mlM+7EEdk1kipz
JLTk2UlnVC1apqCSebwzIe2DIPhi8VA1MkcwQuUuR7dBlIMulA2F6noOjti3NsJ9
LCI3aSEjj0R3gLSBE7VMPjx8PPURW574ue1fIJIGPQ4+cbWCZPP4REwYQXbXpHRO
xCwoM6B4k5FaQ4XUsGinuOEFiD2vWQHSoq1bAfCHippz8cxY7K8qO2XMLC5dZkIo
t+brNx7ZdyvPfKHCDg/32BppCsSgBMokGXyRBYpm2cN0sx2O3Xfq0+JjyNg9y7G7
vp705Gl+4Va6MDxDM9onwgqy5v8S+pmgtumayoc8ImwG117hSbgN4a78flzHoJ9L
xR+IxVc8t1FaH4fqTESW/mBAffCgnhbFjC2epDyjL3Yniuo0HG7NjJL/vhkZ4keo
d9EXZyX/zKvwRow4CazPvNl40o3PaMyKEUy5D6lvIKAgYwclXxVC4dixneH0RXML
gzHfEOXKLqiFsMKaKD+5YaqtNp9tS8r1Htxiwnxq07gL+koe7r5HcqeZNu3fxvDb
py8cKINmobii2Qg+ENyiqRAJeLnMhF4dYWe7EWevvSOz9Z9ohD3oRSG2irVaSLLV
KQTWYtd/XeKYKEFGx8xoFo5IwrKic6Unmu8JLX+PsGDsXaKQfuAllZ10tU8HIir9
jyRvOmHvARE3qcf9QDooO54LNR3zz9Etjmml25AEE5aIuOPlOAQaI2d5asM/9C6/
gp2PUWd+a9xxL3Ka0oxtiehQkdNvLhQ3b/NfzEBH/sjoTz+cc0H4Y3YDtSEG1o/6
5Ymg4h3h9jfnkxK7TpOHoTL/dCL4NC91KeaNPEEYo+jyHMFKMZjXa60giK2iqOy3
DmmxAdO8GDUnXwor7y7tjhdSLJKf8TKTFbofp8KYR7FOOz3RofkMCRH2x1+ZyT+V
JkXrTKyuVpnDb00xnvRa6PiMDKCs5XBaxSk41VzQMGB0U6okbRwSDf7DDzjoKGuF
UhlCogJuOXoLPByDa6ynk0o18VpQA2k1gvhdOleKGh3TTNnaD5218c1Rj7r6wWsU
zz0AcYOfKvqb9eVg1umUAuVGWYEWxEdm0Sm0AWflYTmhdvakRd5xq6OjaXQvFZE6
K3A/3PzBmrI48r5nOK+D53t50t/EIRoIROPB7HvBrLs0AB6FsRz873DXehjCefiJ
6dPvjUYiejjdedK34hLJH5LzgxBFcZy91z761OuKUkRCf5EA5P3h9m4+7VYzVGWp
W8hkKA8yFMdvwocF+3Bj3nFcFEfZhZ3LZeGqgmYPtRaRogR3NeQd5ytabRhU99L1
uP2KETg/oolfvLj9wGcGXNZIK5Dvdyf1EV/b7vcsHECg44/cerJ2Cil2S0vtk90r
vdoy2EdMsQ7BBJUrTDUsbDX7hTnFUXLDipJnfnRgsH5sbFPv59i79X0oUWtG55mn
Sf5JGd4neoDyPox1d90mRnn7h3ORrn+lfYtK8xkCIjnW1H489vPXMNuBwtEeDLGo
vJlmFUF8mOzY3tDnJ/GyP+6MOwxzPBdeLfM9UCc6YtwsOHsjOreACB3a9xM1GzkM
BMXpyNIo3Yo6lpmnJaDXlA80+jMADGTH5IHyCQ1Tfem243vyB5RDOiNnnQvqg44v
v/lSUKFjL1adPl66WfUNaj2cWAFOwtJAQKH+76ayXupJq8mZuLnLJ0VMe8YRQmWH
dUedIdZpzhoe3UmTHOTMbscDLE2zaV0g4fxYMwAE22/cmsE4K3ly1L3mWtZ+4K8+
Qz28/EqyhRWi9AybuLGFRDkdz/Ked0HU1AFtAUycEBrF4P7uAXfRt+QdIAEAymz4
E3csIVNULgTYr7Y+L2BrIS2gYhTY0ldigIqzAF2lrundEjlxBeotLm6oiX52zbV8
GCwgMIJHP7acDGBcQKUC1bGSZiSajrBb9N+5eZ2lh8LLAWQWNhoHHwyyhG2cFPuo
PZhibn4FWFn5qnFlJcFajjKsv6MjVfXpQVhCdwlG1qf5evR2X6X8uz4KbszR7We/
+NXy5oRb9pOPF5aokiSWn8YUoG5RFc8lPVKTnezFn1yJ4k6dTgv4wZLvbu2SanML
bZYqMNLKOu0LKUS5d4kR7UApx1Wxi5fFxQIw0S/anZ4x+kJrupcS4Z1XL/7X+YMo
UL2lQgy7F5TMARGpbacD7W+9yXtZ3gY+LHwHNt6MBkUWi2dcuwuNgaq5T04JXDBe
sggLWUtpaEH5OtBDhuxc8HUbnoRDSEOA+escRGbYWGQgjeJVBzyCJ1kcQplja/u8
+A4Lcfg40BBn8hmDC3heKnQs0utGW3ViHYMtPXE2Y10h8odfFrqNMbbmxB0tNH2Z
ybf0CimIx388EjYVKbUvfWY+1nYXDjwh5kAuEyjJbm/vzQ/mkqYY1lzyPSGzfdyi
TiamPDu3QYxo7BkKkjxLV4erhxTrOdcYxGemXGdIrxbyAsbVrgOvYE4QbsbkG5Xc
vh49HtP6Y7DJjCl/7u2cl+AqYC5OJJ32bl6tSE8rNuj5BxAmqinMgPnh23x7bnZB
BztKFHZjgvCxO+mbV4JBTvRSjYW6VqoWd1Xd2w/0vy50vS58Ea6/dZ7AxoKwa6vY
3aO118+G22s9fSspFU2VF4bXi1SbT+Sfnl/szm/WOEgHtYV31PylkmIPEE2LQQrP
14XmCk08G4IXdDWrnb+4xfn6xUdgU9OhEIhQhX8CWKT6IhT0bmGBqlzgcQZXwbUQ
73mCTcZ3uqz4rvA8j0Ck1LNEH2hGkDELhpUN/h4E/fYUQIKBhSHgUgZnUHrwbSl/
d3JnEJT9sf6CaSBUkwe8tSta+LpP6hROlnoBcVYWl+4lHJ3C+AfE5T0g2PQLCoT/
g67psD6t4D4hzSaKFrTrwp22P6rg4IZxGV4LtcIboF85Uk6dHGOO4KWWNHNMCE9p
3cxr2a3uYtNjxsRLX1ORHznOooc0qhNZq3i9co+0fk0Rr6cwj6EVdVH2DKHypsPP
auU5cEAKlqjStXd6jzzPPv0yujDgkvf+9nCHT5zdxsft2aBTnRAVg2FTJNPJ9DOr
MmsRztI4s8AxYjQAlYEKwcdeGEjicrF/usddSvda4gWAX5rYnpBpsDUI5um6fycr
T1gtDx5XY44RcRdYIHDlZlTUfxERSAPUHS2A9U1cMkrGAr+YSMRhVX+gWa8uVLbc
jX8A3xqtmEV+wsVqwGg+BPbK7tLdQdQ6I2aR65SKEJ61IFWU5bqv7FFR/SC0tHAY
is5xO8bCt0b25aMGT6slSv3wBjg0fONxxlbqBQaHlxP0U269cbxLebU4y2i/o3oW
MdxlcdOwy4RzZdhueevpjfu5yZVah2HRFpzKXjn+g8M8hfpgE8h439P2gz1InBM4
GRKlK6e55aBfNtgOSUajSzcUSaxI1tmLfbWuRpQJM3kfj4/GMrb0lYdZFnh0toXZ
uzgzjTmIZfKV2qBTB4pIQMIStEAfak1QzNdYqi8OWZOWiYwq03uPDFhk7wozCSkf
zHnmrdmo1bCVlrVu0rW0G2WDzaiHbEPbByfmVuHhX8wbiWc3lzWRKcz4ZCmGyjtL
dQDB/yXdpAUpQczF6GjhFrnK5pHk7BIvhl7BCDG0kqwo5Y4F6NYHIIkKH4LQdWzG
LCen2011KlVDfyHBe7p2BDlWO2dYQ7ZlQSAsT20W2nX5iEDKbw1ROO3UWnpb7rmf
ExHJvauC5CdysdHDzEWnZx5nL9rFECSIGOyA0SQBxFQU/p0DMPzALv5bkbCLuBYP
gsT3NiF9XRvJGT3U0kTH3CJRkY5UtPCtX5kNyyctMjtCUzfMBxIOXobHUmI80xK+
T7ZyWjeTErwLKM+etBA7xzAlAb0HhPSZ+WwLn0d+atkcwWw52UzCS7ozh7pV0Pwx
m6v5xOBzcfS3ZBvLKrC31orzdMGLABxw6n+8LpnHSu377wVgksGzi7AHXneQ4UAS
KNYwPJVcIbHhOs8RGcnb6jMwnZi1b5WJoMv2TXCqUwMnEB7HLkeUdRWJkwN/fV8g
IVwWSKKlWRYtpoTtjST2tErCYYaN+u7OHSt9WdcJ4bxws7QB11/uNU/JIl/4k4Bk
WUR/0w2uchtwY+MdoWgFNwguy4x3zKqNEpD96en7u3amdXDR0raaDR+n0F5srSFf
IRctSmm7fKTuYPiSjemfEtBwdWNKFrMOc0F9gDCEByZ2gRvVYNqSU5KHEWLmAMhH
z7cSctLmhT7eHMIdEUyExxW9xnWxVKk6/WtyJvebrAv7pa61xc9413NcsOMOYDah
QO18zVtw2/rBvJvXGBN9knWu8JLBIYxsbr7/KRs4XXQMSm7z7o7cZxVTxZy25zu1
jmSwZ4wxnzs41wmQBOXr8WUEuGfyUw4xl2jxTbG/o89bXrzpkaad7acpOykfPihe
Y/n5X4Q6EBWzUecSBHidwAoR+g7FK8gmXyfMGEsK8L0oVV7jmLK9JtkI9fn6qUka
4NPXmro8ZHDu40v2igrF8riWXQdbZejObOrdXOQrzcxXL0R09c83hQFrhOWcsndu
qAfVwNZUPN22zKGxOwLiEMWlV4C5zLunNlY0OORVUxC5JHo8nXw0J05g8IBke3RM
vnCfBwe6JC1cN2RtUCcrV18z0EFOdCjvKvfqQW7r3euAociosPNHWLhtYBLZOcxw
mfZEkv6VprvM6N7TGUAdyr/A2qyDuNvMEXjMwVNiczBGAzwJvSLsyzJBx82vTzf1
A3bMHUPvZ1S0G3A5AKcQBHH0NG/MZ0w8YTZ4fdkI+endFvcQGKn9OeSH9QSo7wFG
h8B1i/VuUc9KnxkBDkjSO7PgRFuvh8/LXbOTKgVzUaKbpBO+6kxVANhXfX2MFVjB
jDeCP4iBNXBHFyr8bG76r8o44DzIoPjBo7KxtvBKHA7bQIS9ano9qc/I1VJ03qsG
Q/MKly29qc9NBAE4pp+iuQgO8ckC7A9bb6ply3+OZ6j8xtkzAQJvC7rBQ3OJIwJx
759pFTh3ofUmkdU6xnHA1TyPcCHcW1vsjg/GC2qakHmoqlnNG7F6GKsIYrTBJb4L
zzzEKT7Yv93oncCLMXbvIroLuaF1+f19VyrfepjrLqWB+Z41oea2RiH4NS8t4akG
Mhe7DUxMz4byFrPv+ZrxFMuGYUala4f4cSGkde6lyOFoDrRvKBLlppe3/NpM4tMd
jDaB3B4viWwNbb+sHKhLQHJi3Z7q+1HomeiN4MXhx90X8JvIpqJTO9tHBEhn6LCz
BCizNBuQs97HTymFyovh2M57qbYlN+W+uzYTtfuwsByw4dzVnPvDBxuA4QwjpEW+
3y+aTLV5jj1zrGLMA1jJF0RSKhDy2YYmV9WUFxLZHLkRHhae2ISfFh4CLdUQjawe
slArW3vrJTpAE7cRAh2ysmGNDswt4IIzHZfLfw4ZEbd6w4hWlPrqOJbptyhHckIf
5OWBvjU2eln1bQG1QGSzXMZnUJSlgrlNpuzJnaiffYWrj45E4nSg9L5McWY+zYuK
ZDwdnNxk5SX35Ho35R+rijmdzEu0HL1Tq3d8e7y7L0eEaGfElmUoOTnxUdMhADzA
ob6ILRfCO2X2LyPtkzYIp/vR1EIUUSOknttdGHUWivaFy5aiMT6+1h7MJWI9f2xK
rmqjzfnup0OjBmBrLkCYQ/LplO1CR73wIuEHbEghppQ886Q8S1y6Z+KvosVGDwG5
W2Jpu91NvS4+drwyucXjveGqYsuMnucEcsWaSP2LhDBxO9l/9opSOxvXQ56JFfJZ
x75uGhMm3LKA4FX0isMjGqgA7aa0RporV0YAj2f25y1zhFppWYq8CfjKQB8PwiP0
H2TT5ujRA6DSbdEtXT/53K4Ub7XfeWmbVUYb4O0oXz6AGB73RydkRsd+cbVUxOg5
fiYKvziXQHSDI2IiZhLboRnk+IMI+EDfQOHC0rpxwd4BmMkp6cEIWNTBU3MOGcUV
E6oQnueI9Qj0yr+91NqBY2FzI8i7ov2ee4gNS36gJ0wh7cw0crs6p3VAyZMBkmdj
UjmkHyxHQn+6Sc7LPZbnAA48NQwBP7imKBZkEHRBNBpUwZ3W+vwnGyimrli6ofqG
JcP5bPCVUr5ubTJHLEcd7nhh1uGwew0/N9quD9Fvj/RwN9V2F5fu+VkWfc1oBmdK
F8YRKxLYUETePMgJOaVjmnqnO55Ptpw5pkqO7osDHYpoj+Gyx1U/DSWZagTD0G5X
NTIJcqpgWz1zgTP8KuCcCMRH0OVG32TZouuy3RPhJ2Q7YexwSnc4eFOEJkemGFkA
9rNKnFft34maQO7vnVpuPKDC5lf4STj8PCNtN34BJN0Molk/RWrdxey7RVdacDrz
3eaVd2Zg5Pn5Qf9WMH6hBJVvB5sgI1ST/ZyH5VQWcA/bBtuEjnJNxMz/he0ngV29
0upyTsBjdeW/P8G4ipX4fNy5Uel7ZV+80Gv6v/yHJjCacPlgYTbZ9XgrCt5Zk5Qq
/58IrIrBxMazegN3WT7FyuJVnog5ZfhGLae3PcZZRbAKGCaaHE7WG9yoUdsYNPLh
EyuJhwIV/SnN7rxQDVowcUxEnbhkPtovCH/y84fLF+SCDvp7mHw7EeNCZFuDDkts
TLLKSXCHO4VE0AiwhswS3ukWbBfWIzVWhRyW63Ok8sQbguqcjKAw9nMBIJXTJmoS
w1+66BR/EOxLfMluH6zDrmzO/iBbKkHxdjqSm1a4rmHWQfFOPb3PsTNh8vaZkVDd
+D56sEQqJ301U24Q9K3gy6lC0U7yYS/g533bnGnMyWlHyxofHsp/ImS7Bi6BFwp2
LDOcTqskm3AH9cvcE9QOUNYI13DpW6JCKyrdG10Tt7rVYNINpVQKwdYUUmqq3mkF
1knOAtP14dtQeqdwhGGKpiEQ1G+a/cECSQzTKh2Vt9xWgolv56BU6u7KVbIP4wAb
lsJAyptQv2pr7f5vQ9bRBrPCmHoI5mklH+ESVtpI5h9j2OHizfRQdD8HhmPNdQRt
r+vJ1UrGWLyWiINoiMC9ssY+1UXmBMaHeNYsZRsi/BEYDBSLQ+jTa/wpzkYZ3cAf
aGKtpNs/MRMktazKE87njXSHGMMirrDJRQM2FlcPMopcpbR21ef9FJm1KvvDRS0D
zpeOYGpSN3YckksoVNmsyxKCsI5MFIcvSRFL/bFhW2R7M/o4nQCJyyElI+SuHaFP
o9DjHt4KKaQgwpynkWN3diCLL4xMJ39xPHTxZNZmFdwNLV+iMQPfpSrh2I6h/wlb
aepT73ynMm2IPQK+3lQX2+7Uzc9m97G+MNuZ5sner+/7MX4lisqZnIMrUpR32YuI
LdfYTlEuoHKDjhU7EMQcNNBBvjff/YBT9I8HOZheUQiRaHQ0rjaajP/wlzcGh1Ig
d4wit68UsS97rJ9RaXFNSsleFTbrc/BeVWPQYCOV8tlsGCYE+2pZZTOuyLhqxE09
/MqeXsIUdGJ3iIJlHjxfs7rKKIlF7S90hSoalXqG1qwRrxrwHektMtVXxxyD/d8E
KL8oikuRBYxoJxFQqaTKqMJAGMQ5yrVH8zuRp8vWC7PMi0UNxr9fG2mrUeAT4oWr
2syyuvSgmbjMUNptZv0kb43xEfOVf6p6kBGPMMQm2XN4G8ULmogHR1640+pwbwoA
RGTxQDRoDNoYDcusOwibahxQgrzjcjdF0j7BpvZL26sqt16eGHiZ/fiyW1lOWtFS
mWxL82KPVEursng27ogxcXEQ7WD0zU6MpWlOx4/4H7sCW0k8bgGbpzBpvjkPx+OJ
BAV02P6eOCJ7cZ40nUsWFcTumuhSuuFkZXTKg5AxWr6a6ZSweEdIAgk+wtV+oYxy
9RI4+Ki1Jsqp6r/OCHUB9Fmy5fytdEDw7eXgi7mW3+FCKOGI1vJMTYyOQXMZqb1a
mkAPCA3UK97cXI8kGxnNBezTTW0NrOWeLCLpD5NNHqAIcQX4FAhItTNsQ8ygt82V
C1SU6nhnva0KFcy8VnEkRdBdu6XsQu4ioXBaG7wzTYlRBn6wqd341VIir5SDgbpT
k/k3VnXpr/NMKmMsW2J625LjZGo5lqjJUqHqUNMy/PEeZEJpbCI7aXOXvJOE84W2
wzLzxWetxQfTOuWn/2Na0UYeVZThb8dmZvPt4BYjgFyBK3YONNuMXsXkUKmIq3E+
YHgDrV1Z1e/malt4JTH1rjp7fdkwFyZiPT0PQ0rW7SiFoFCCwdhDvMHr/7RRB4UN
dz1ITmRbfgzqM9eDuTah5c2SRUQgUT+E5/Nr/dEMbhsCyMRf+SENYoojVbgTha7+
K295fZlHHBQFDZ+mUC/8CnDa8QWHb7SNbf0cktnPkPxkTjX4FIW9InUT1c6ciFD0
+iNArwV3n1UIfVQsosw9mw2wtzNoPJY8joIBk6eHVHzRbyeFdz272JSoYYorUARy
cPkE1znsM/x/aqj5+GIve8t10hu7VZ2CWL+VmBTGM93mpnc9Fihqb69k88rrSpVx
Jn6sXCjE35fvEL8RZLWGriG3epj+GOmieCxkwVgIyyp80ksHIQR38fKdbBYsNVLH
6gEVvXOzU5SVPeXrzZ5YrdSqffACBTOTQGcQTypSawVu9Kcsc6bFLKcy3lex3k4C
Qr1fZN/c3OuFEbJtZDey1CJPxKVAmSJFrA9u65FRhFySz7dPop9uR2hhbJTP+LVD
fjAUr93Hr3bh9NZldUPRskz2jrgBmwbmyhwGg/fhKUD/A1KfFy3yuGU5PrN3IMdy
A4Y4J01dqeUEI0/jey7CJx1309CpDU1oQqJB0nVyqePjB5it7gezBIcyqV17Iiey
fLuu0JX4We453KYW8gbDpnLBLhMgsA8G8hNPhOBQZSbOPfb6+KANfrY1HxQ9Wfq7
3bJwfvDdpRUjfJxy2Zhe/9DBHrl3gCHwWOV5NyVq78U1PfszK+nvNi+/E4j8311A
T7jRSW+haJG5/ZgwMx7blyuFUK/njCiwoiCY2PHP2C+Wf+FgQtKsENwK2BklaeCJ
ibgMtvrAhjjw6lgtT28Wt9lGt4BsLbwCKUcQNp25+W3d/DH3dvQE0BN+PR5rYLp4
RLg2rmXnMiHbyOWJRowgR86R5LYbaIUB1AWOw3yGeA7qgA18z1w0UKCQ7ajj2tap
vIMEIUTgEp+rBPNAI25EaWzHDSLRQMAwwAVOt1yFjFQTzQmFY83DgD7JZTzi92RO
0JjGfMYJtwaQuZlogccV43ZZ88VWeiwS3gl89LmC1UdpdVUXNDxI9mCpLRkfaGet
uW1FWsxo9pp9doiZG6eF5Hq6slI3wsTDZGz9Pu2JBY66PltU4315/nMg1YfNaW3h
94B/GbOSRsP3cyu+oMxvqJOU6qPZMc7qNQYsxxyZD/DK2yvXN43SQnxD9zeSlnEi
1rdXaHezOm3nW5GKxVYJuv3+FcgcEw8HibdqzJ/pVgXnGkgz1WIviR4MmAobTO+6
3otPJPuXo9vA3zxMZvAfdEjp4krYFPdFkxZZdtSnfcFJXM9qJnpMZQZgD58DoEHQ
QaNdgqw23QSIFsUK70lbX0w1c+oqzWiPEsHfEsI6OzRMgpLWw5kvRxIovnV7CvZL
+mLbHTXdkqtrSBkjXm75gyZMNgMF8gGx2XfOcJls8c6EYG+qK1p/JkI7/bZzPOS5
OjlJxgrNBsxeXzPlUE0EAowFJJAlPrsx+kTI7uvsYgWsiG6s00QS42CUhYP0c/oZ
DTuDtgrxIDkrqh3GdWrqAowFu5JQ042I6bTwbQHCX/i1pz0qivNZ3vwx24Wovgir
6m4vbX6zwEPStMmZQRHP5qQBPxJz8yF/J8BpnFATTB2rRHbqKxBEG0MLBQRRDmRn
qJOnnAk85aTbTW4wAbmacAlTbjOl70IM88Bcep+jByZXkFuQ70spxFef5NwagWCb
kSDkzRcFcopUEePcKmKxz99ao5rS/EpkNPspvynXWAQEnxQkjcrHrEFqLZiXpDY6
7Itxja/L8hnY9Kybt0NSnCYay/6xqC4vIDTaGgiT9h4AREBIcRwb6/m0pMtYD68O
lxv+BBqE2oiXkpvzBu/l4B/mMeg5ec2UkGKa0/PEprB3JXQuyot8PQ77ZYRR85uf
PhinJ9uZdE2cPGLm8h8DL3kP6yM2gkMNKp5egbKELJb6ZEf4ORU76b0pVQiz46rY
FWsIrTimuOjPp6BgmIUttwgAo4RbSVK45YpYpc3N41+KNmb86MKBXXwnpMxByIPw
4DR4B+J2o8t/jiuWWayN/gw25jnIqlpif77Do2TelP3/2HMiwIxzXxtoZAA8KW+A
hXUHbXNzH5e1BGo9XtXrD8rIpfKhGEq/hVhyLQvcLWTEC4VXVD2veHeswV0GWcHo
XKoFD2XsFZPZLfAhY2+bbHnREsQV0K0MRsBOpnbUaofYCx2VHayrwQsKWaWjcNp3
QrFZEp+w6Mt2U6QIhXJt15eQQaC3otW2/Mdn4sgdsNoGrgBTPSbfkBAN45M/vJF9
cbh6uSuqCgU+k56p4zD2NfaDz9nS13ZQWYJ3pMHdZ4O7//UlfSGcpPuT1mLHNSh5
Co529Jk80TZWuBhv0oIYwSukEkHCq+hJlBNsEofUdfk6QTTa0AP4WRWVJX5Qg2TX
bLaKIGMOyxRP10eVJUmGCDvGMaH8ZUIMZZExxUaQJlYHPPee7nRaA4rFjvhuHO+l
QXsLAYm2eW7WK4K2TExs9RiAKJRN/fl90XAeCZUJHP5eTICVkgl7Zf83CQGV9M/o
SiR1nkFpbiiHFVrkjdISCuPt9RoWaZ3r89UOtOE326pr4ComARUe7g+169pdhqge
f17cuQtnqQheItlLkVZxqsNzY+z430AxJF1C1WTffjZnR6hsKoYUuRgNBQktp8Pn
tPCKyQgXkY3SwbwVXhOr/t/GS9oPhA3w0EIDgdQj4OFOoml1vODtwtycfZgKUmHg
9Igh7FnjoanKKAWMTLp05TNsBAy9m/867z6W7do+5PE4MCBlS+0ZHzg6JR+BOmh3
E80blgTUT6uBNkaCRbvRtDCOFtI0Az8U9DY8+4kwIDztr3Ci9fuXeT5/lATYhRs9
sXYjkE9+8L+FpoqjUYGdoMiwjws2jTkAxDHtixkHvicJLttsQOqreZv0u/P9B/GT
GDv0DkJegB2Bzm9+B930gAdVVelnitXYOdxQWUrKss3FoujUgpb7Bdm4HENDgFeW
ejI2x2O1NZBbepy4+8I7V2YQBAsClUO0343MI6WSnceAr4cGUwi7v/3jfeKQm/SD
BHz5p2FFE13FLROSEdoSrLkWHonasJw2UpBTtAMGCPmBnu+cIsiO8k91+ucpU2g8
b/2fIVx8VGGjkob+yKEeVXaiNfqLk2FxwD7NBY7t9zy4Gylvge+E7wY4dlqB71Bd
bu1d66KoJcKJMjgLRJbEED9VPwsreN5e8zvq1dEspy0qV73tozd8/IH0WiC/2KPb
rC7TC+RDxW1kXlrf508nWTImJtnNLQsccratpN1o/mz5ylQ0rs4mu7WIv6LXcdR9
rf9XpaLKcRFhxlpkWi9xCRkWf8cL4/AW17708M87pJaeFX41Ta4SiIXXll2yr1eQ
MgfQKOkNOk5Qp1IGJ36jUDM4lOoidXYLiIKBV1qHPQPZ6J0dfdkspZHgmXWuFr7f
FEPU2Kz1thuOd0zfat8TWybniWy5iE+l0536rS3jynedb2F5qvfX7/HVq14XLA5Z
K7ycI6u3ZFVrKelbcokgu8/BFfJC7dsEtNRIEfoqjF8MrGFUOb1A4tTEOM0ylNcB
xj5qu3UA81shuZvUY5njAl5IfhlU2BXwFb1oYXfAN+/WmfOp0qvnSM+WEpfukCB3
r/wedngTwdRZECrjKMOumjYuuHeaUEYJGACsE6KjlPKHAtl9Vc0OJMcQxLAPmuuh
KMQlcIUTsOCCcg9zOg/vnWfe6q6HbOknPKGQx6r+Y1M9YsXsQ0rmdMKzzqGFLhCe
kZMVEhu0k6FVrTZxl+AfhHZvYOKho0zk6gbkZz11Gssjly4F5tTjh7rfAtaD06wT
Pas/oQiSeTFDpx4q63P951PcpwBfo49Qt0CgrJJiORo/GChBL2wbIqUxG42c2z0I
9Dfw/S8JLQT1dD3WtcUI12ar6/7MUPls+9MDuo9cO0RlZMNTogIP2BXf8cmKPle1
HI4mephaoybZNJIrh4m2e/hoyLa45gBXV8DwI29Nil0v/Pitao8udyEgI4TLjkLs
fWDk9VggTzN1fGwLYW79bCcFEdEQO1oCPXQQvzzCLV6LL8NKZU3BeNJTSSPhQPmA
wp+biWidxEP0yFncm4Wm0zTVrj2EGrkmpW3ytzyQtxZSiCRiQSo8QxSGR0AB6LIY
eeAiCBzcyDVKqxdrSmfucMwoRgTzlhKUw2rjx45LLzTtJmWzJFSrbO4N3AeZaSiT
5OGcbQSGZ/hU+uIpflmkdVSgqjd2+IFZVJueCvja8bYGFmK7HoORhK+u7b/kH0sE
suZAFtqGxm4nJyPyNGgwUCLyuo+Ia2gbL6EmsPe2r9maPbP/LYugxu5p8Xpvcv6L
ehMPfzwi2jrU4wHMp3R5ZzXVb60aoubsh/5mOEcy1NsWhUmOXQDZ2lo0pdqtYpku
MOj2LCDUflBeHMPsLZsaCNkt++3pM8DB9AvKk5JLDa+6vJhKYqzY8lZdOhAQAcBF
PMYeoE8rm2eM9ecJajZU6jpMBbZC8JefUPOSBKBP3TX06COx66ROgvu33PF4BmkF
iHQBhV8bUjXbJJGfFSTxDSmxztmG0X89oxJJnZwBQSg43htBMuqmJNVR2XgUOCsD
ZHxanMD3j5M00g7iReQxvNfLnuFsVSkmROqhuxpHcV1Xr6m5KgfbeYZTCRoUIYUi
r8l5MR9T1tABzYX8VitNu/r0zbZ73PFiUl68B3id33IRq05+qtgfFvcbx0fnUFjy
rdDc3Unsgkqv8oXLg/wYduF8q3zZJNzvGckI5fw0HfLilnmb8wAnf585cUJUevjM
JClbTqXUhiuyRbn4btJH2p7IVlh2cIgSN8NNbQHnihpoEzyfKM61/OI1988a/Oc/
0f2i4C212TNUBiHVTsQcMpnNPToRgkp+fuSMdp+5ORxalMknkyqYHY2cdwxw9oWQ
2sniQbN2HjwSj2txDhxLtICcqLDo55T2Qn02rmrWJ1wKVi0Wl5Wviwtp0D3h6oRn
LBzcFlGyM8tGSchbAaboUzsUMajUNS2PXJHU0ioIQ2gyCDV1nde1rQ/34V5YbYH5
7/+jeEsbaia5go8gtA0JQoUtWpT4W0TajOHK68+0hFc5AiAIV8uOeg9dP3mQz1qR
/o40/OYU2GilmQ7NtZRXI/WChLFWGuUWstK4ou9+0IK6L9nuMbiRjb/hT9eNI5XZ
qA8cpTFw3FUyK/TkDgXP3xVkvN0hQBHGC6oFWi9t1AEDVphNRbL4gIpManj/ceTn
NY/v2GWmhEgqLsd84ApXWfp9j8ghmZGBzSnuTrJnrQz/VNaI9Z1TiNO+UcAjgQtF
KMhYtwAzPpNKbvG6wuMdyKhPGQ5PBB3FC9cH2vCl+J7PEQu1rvZH0lAs33p0TKap
Iu8LogC6nhFfoReqrOoDkJIiO95sTHAEgTRKmJpHg2BFeU+pTXfEPw+w1Pd6m8ff
WQ/e2L3OS6LGNkGl60Bqhx67B4QCUNYPIVM3f1u/0KnOk4xFQeRKwS8BkG+rRnSz
DzztEdzNy2gXEg4DJWorlKW6/QP2s2kH/v8CiUoP+8o/Ps8BNtwTUCHn5SglhQpw
gBvNVOZn5hai8l96P+lEwJQ3OgcbUlUdHGghrzuUy5RAzaCNFVYdvKlfXnRW+0ov
Aa5wZhSLjI+pat3qMIO3RtXCwJvpGnMaFp6KoZHaMmwRWgs7zv/AW2v+iDmSOcuC
pkjrq1TppMFqiwMxBoZL1gwlHQGf4a2REznTyBwfCmd4SoWVVKwCfpAWVVnk+ltn
37Zhcy8Adp3Ts06KbLYc3sB6Czw3Xt/QqPigBj8YJZv3IT8xluotYtlk6pN2NKwU
0wjFiN46T2OwE0pNq99GSFthHSrVr1+CeuzhIPj+RJk/mORv75x3498nc1aGi9bO
RWdMykO1oLBBdy0sHtZqZwh613AWzwNS3klC527HxtoioL6qqhSttHwIcbuJV2fC
We4G44XudaBObzGAU2YI+bz9sefAFOpPiQgLVcX/shg4CxmXxAJEkyWA6AI91VTO
bA1Ru697RGWMVjXf6S30a+0pOM/OeDM6w4RxnTmERgfG2Gh8rNu6naQlKkVZhaTE
WAAPXCwdOd/VkRhI0E2slTPpBdXzRehZl0/yxicv3OKRFeY4Hx2GWji/ZvG4YJQt
B3dTDjrMNN2E/A4L587LE5Yy7r4K++/RhTodhVPSwzCNTniyEvXxEdJV23ZgxOz4
V7/OZQ5OZpbGnmc1eAk9V6kTgVebUyaX3QxfpEWGSAx7DHwav1WnvBMLj0Gxd4V0
SsZ4ZAYjo3z7g/NmDg1tMFUHbMFB/7G9fuW/a6vRUlsvGxYw7+Hu1Vq/hshbpIr+
afyBJooCJzkeT5uld4rTwgPtnCghgM324sQC1AztIGHAnzrIk2yJ320Lep3V+Eyt
xxRbtSHrSS5afPq1v1jxYQcJAZOmhzOLMXwBDNHg9fQ/5w9YONBJR4fsTRLZ7/Ty
5LUGTe2X7m4RJIitXplLVNHSINmgXCRDQZxzCyPREaPvJW8vvnbAj98u7LrP3EKd
9BWyhmD+/67vZbcAK7xS+oZ4g/NkGe1vOUeXrYRSKXgpInTAySXuM3uD+i70Lo0K
6QP5T93CZY9G6Ppsq9r7SARpZyRwKduCSs36FFci8WZ+yVTEywdS2TU+PYKZ2W5s
axp4yZRMFD6NogCL1hXdoCEw8tFCpXxI11ETeCRURhaGiF+LAb4USC41/13Ln7mk
iOP1eCPahYBv/lyXQgHA2RKrSecVAN8P/YEsBNN8e905jfeu8TiR4GQpmhRUiJOC
F11oO6Ju72VA6sfOPcHmm9tLAtYEI5Keu1hxhI0gTG2HRWQ84hZ6x0HhbHdyM9/Z
jr6ZaGE1ZO3pSXUcHPogihrgddbddRBm+CQtVlonZF0cXRZwp3WNVIyks27W+sao
Dm8pwqyGJ25whakC8cp4+l+IyGvGG4cT1tIvVYCMGqTUDnU3KrCOVxOhGoG6E460
fp9iAORu0BjfsfqGQNuOZvxbJygZjV9orM8FNUIyGKRNNZTPw8blU1vhcYL1RriR
j4zhdhq17+kMBHR6+dHeltUGn1Cmn8WZds20S6AoU/NDNgdKC5CAbhqmPjcshP1e
Mt9P5fUqAYKSAnjT/QwTPUV+eCiI1dyKKbsaB1tZ8DaWvFD9SCKKm7cYquR77gnK
/ZpRpMxQv0bhM/Rbowvovb8T9Ntv9Z4oWU0jh90UkCatlK8rG3XauJKz0y7zX2H6
5k/M7KnVd8RLVgCsVey6OOwfQX+C9laAK79oMn1wQGFgXr5P5iYsKAnfom6JbhUj
6ZQjoh236MrIp3x2luO+JiRZgF9NYCQ5ggJP5sUgxI+gt8sPOYQoHinhmOHuiVGC
GkPingZgfj/7BoEiQYOXIEo/Qxx6Qe4feB6G7RxOh4LG/ods4LeSOt4xdae1O0zu
PI1YFHLBWnVwIjqaQcwM4zirQ2S7U+hMrUCluF2K6zbz8rFF9Yk0FEVWTkXM8oV3
8ZgU8rP3Uon3VIHMPKrBvfYJ/fO1ssRpUSmTcNoFOpOsbp0kPYHb8CmGinDequIf
SlrpBRt7NtimuTVaJJhYz6UBpiS0pRfXG1D4IOHKkjWXYRqS2G6WGK+y6Sj6He27
RDqxYRJehHpXB+wOiWxNZe9bJNAs1fVjVkgRqfzgwM8matzVWDY4EswT8KcHGZpc
4pmJGaGMGfWyhINN5NAYffI1izYEzbU/9bgRg2FQLZWubqEGquy2MhcAh4bbkTdB
SOEG9MUV1Aor0Jwlhn2E0BtuK7sP3dki7mS94L4UCfqTAUnuS0+V/ViszcbLxckR
TuUXgpncwJgZa4vhMJ6lAb5LgzvIGqPGLVRjhaWbRipkLHbjlRl6k/JVRWB7yNvR
mqvdYp4nvpcilRi1P1tecsRcE3baOMMb+QIGRkaLtL6r2O/weYgFC2W+wqvlpPL3
8AdhOzkpV5gpAe7OMcHmNxy2Z40avahVeJ3WhzJ0hRpEDJekZ45/uJvEvC0mpaMh
tn4t7d3IPrW2EyiHAQF83J2KDHpOfo0hP/9oLIydmIo88HYqyPXh8gx2A5XXyvzI
IeBuKTU6Kmj9iLZ1hyHtdsLbtEFhK6VIC0fFIBv/fCWAcOX7uU8suPRzxlkw8QF/
gHuDjRWtPGYUFNq796xBolDgxA8v9sxhM3Wfrpq7QxXiXOrXK+IaOCw19C7BtVo7
/wR83mOQpn7S1yIeF8AZ1owkKwv7mFA05TfkwlbAIbBVkbPeZrQgubm2r70hnGRA
W0HhMN2jxKzfOhK0dMPX9AX4376PnjKOyA9f7fsx6ZDBs/ObQSZ14r4FmlOIlIiL
xC0PBX0RNgztuM2r1D5pN77Y0hmAY7AYQJZcOnqFn6Rb+5hpe46Sru3vxg5Vm0jb
PK2J43m1KKika6J4miyDeOmJ4RmXdGxCCUBdvYWy//ITlIwZv5Gi8FjxX5xaFPzQ
wyBH9vFPC3xUV5h0o/dzaHgQU2h1apwXfgcYZO724epPw+DiciYrns57JbB0OPeP
1fNhkXdOafpk3fDiSX+ajwnWhNz+a3nt4UJqrukrX1cn/PfNB7W61G5jYQp78umr
aHXzl0zkv+PXOFIH1lRbLYIPKK30xaHI7aX4JZAYeZJALvgPrr1lPfPOy5vlv/ni
JuQKMLH/kew2BdOcwtIJlkhIgQJrB7xkvdl3WjmLKYJ37xNsyLOuQjFEgPxvOkSF
hbERWSFWyo0NjovbypDMIgTKrvvGgI6zC+aO2IW4U/nh9BGSwTSLcRsCq29o1lmR
A6yvyCvbRAegg5nFRyxV5vPGyjbxxqeSwg1wtEoJN3Nuoi807HqzdoXOuAgUuQc5
O00/xdjexX72d2MWIwNjG8N2S8ZMQ48qmqnr8cOObnFFB/yDsROW2r9f/3JA8oJ3
7lLoLon1G61mQAGtWlqS5cekcIGLP0H/Q9eaUbZ3ArjEXfs4F8ndHuL53G27FVww
z4vJVEZEOF/Gm2iSm5EhmBFitv+2Hvjso7GbNYVqyu4FzBq5SrAuB6Bu0OuLNA0V
GBzDebSWJNEHavbv2UIGjj0etFo7GbwOnPBBFUFAnNre9k8Q3GTzyoVfFSV6bClK
UMB1Ytc28pQ3iQu7U1vWzq6dg744Qvp3RkpNPt92tMvFdE61fVz9J03Z7a4spv3b
VxK0xWoSNNr4MehDN8CjUmO+OqJ8WMvFB8UYj4oWuMOwtFtMebPwD/N//Tv9EhHK
rWQKWQFg99ezlkQzhsMUbAnPmJRUhp9Ng8Gd60732inrRwxeZ6aflN291GVC1Q5N
2hY5IhKjxOVGN6+UIpU9Wg0ywBoVrviofUy9e/nHov0iAdxlq0NCbezbtqQcju1e
9yvYQy5Eq6/vh8sWeEXFMr+zBKStUKaGB87VWGadsLzxF4Lg4OuWex6BdPb1qRx0
0zZLTHiwI6z3ERVDogTHecwlRX+rsN1GmDoaz/oCXdd/BQK6+8Uysx+UNsy9dtta
v+FRyJY/pkBJU0fdY7zNeVng/bxIW8fZ+uEaHdykCkk6Y2E/iWI1N5mlTI3uheLp
6lMuLdClXXPNRUB/5gvhxFvhaN9vrBPEmJVAAXJT0b4NVXxm8jIiqFecedkap5on
k2QFsJuXUPqh8MSzqFjjVeWx7zVUrYtqR3e3oTIufAmLHM6PYWLjC9L2Qayd79Ck
PXPIOK4uPeg0Yr4YbNdifYJNLe66g3CnIWRUtpdhLZgBrLo425LYcUd/MfzOaoi+
qOQ6AwPTWQAb6XOWPjvoGQQRcqnyrKoI5fQnvAHKY23if6qI0QCk3pTevxUtoN7d
xz0UUKli5CuDaEskVbdjU6F0nKqhWtmxn4H69oI1AaxzoGDZqvr7KOCTXTRvd5/Y
VLYkYqmk+dRr/uVVMSeJIq+bwDRczZJctVxf5cH6NEq/x+GgYR5wdRPvV4XkUcv0
uf2X5axSEWFwPE6lz8HcHlsLtx5nJ7HspQrn9CA7Wmr5v0sHXOXnZDX+LnR4xHO9
iH9WPkDpgCGvb1SGQziu65xyEc6nePmYQ9VCRWt/Im85c1MAcZUhXYxeclGiit32
/GD8ima5rFFMW+Dx/6KvNnhAvRn5Xxcfq8QfRX8y5Eu8zCebQbZ5HDWOiWpnHwun
9Hu4ze/OEvNDvbHJdYHe5q+jF7WqR90HExPu2UHa1tpgUuCumdJeIbV/jJ0i+clt
BwIeAQc1nA8eVZLKwxuUzs1On2vI/gGjrlCmfzZQPcxwhXX8xMhZhtc1zQsgvWER
s3wL5imMSYjxwZr5nzRA+zVx3+J5vaRqXVKzhfeEmr9SzcUuqS7I9xHqgyS6XKbi
G40l1kDdQ65y6JoEeT0bj+PeiPguw1WleTIRbFi7K8GVAAUVStS7qML9XSy0prk/
3/JKhzPVI6PB/0go6LbD5O4aCguXAKIfTugHiT38GRFzVn3cIhmWepiOzGmHy9hB
4kTQk4n9nL0h9uOiP94LEbgMUoTGMaXWaT4J0YdRobRat0bGCkUXy18nKZQ/H0A3
fHTfHbaWvQ4pBQy/b8RK8tEO/lhEDlZP7MaAtD77d1bb6jbNtccMuQ6O25MMpedy
YbTSyNpjxfDmI0jn/qp2yTsofaYRlODqYCKHKg15FOxlbT9oB+drNL0vLwDJOQPm
0baLJGGbHUP3RCIxlt5M7qkwh52SvSqasyzvOkq5/EWpkyUaEcMrHpmSPlxiL1wJ
yYj9dOXdiYPWOp1rIjmv3ie2PiseX9+z1AKmzAQU9/ABbKMsdxSWLJmBgl2dwFxH
UwjwFP6IWU5wLF/2I2OtlrtJW+H7eLV2x82UlvWn2ZRFhG91pzKhgL668mR7xRwP
e/kmIDPk/+mBrieydhUJWPJrz6pEfazh+QGWjp8Vt8fmfUMheRJlKPYFiLoLY/hj
54DP+0AZdd7iAqb60KczyB9HdMXIXOJ3308R4j83PMQVP2R13R1mo3KH/GUdo0PT
3Gjm7xKpepfiN2Mmhs2F2SbBMfNqR2XW5qSVj7DEh8KbyzOc9v2OmAkvg2nfEmNW
RF3EHrk9E+qNE9c2PI57o7OqRo4koJclrGGf30lA6hvEFCTCH0zVa9yw2cHB6Dke
XxgDAiUXEraMBNd0zIN6zuerw7QaMhBAHphUi/2eHOtIPtsUv39HpEUqi/vGKMPU
AqdaQNlkM/qukmNUOW786BPuR6+GUqnzi47bHPzpCHtPYNb67bj3hl+0l7AhTpTs
m/fBD9k1x322nlEhAwmXMgHetNP9PXt9rfYgfLIqO/+8rzMVPRASLn3z/lwII1Gd
Pe5gf0zeGm1FdQFY0UiY3cNBxadafyfJmJ0LgrcWSPeouYddWCKL+mKkgisHZPy5
hB42r6cYkuwm35fG1lsY77rtMPALhtOBpC/Yzg24Zd0eQTUyrw35CZDLQ3krkEj+
tkbObwYSb4eQowCQjvqwcKMpbfGwuesDn18gyxOT9h+ikm6crAlafRh/MVU+k99m
eb5wIX1TArVCnBNuJZ30fmSO6ZekuiBNa7gro4xK8eX5UO/RPdfivimIk6jZp5E7
XA9ZJcTiCkEHyqKD64Io5nRMGljn2BuLrvPJJsh6L3KUhGbc7hWvZk9nYHC/8+mh
QmRH8QWKEhuqRrZJcm0z0SLdEkaKafjttznXkzfKE0F7pOA/9p11ZIDMxSO9Wuo4
Og9fk+cZ1PqosU742xTu/U612X4Ck7yCyGwM+I8RdRklkpmIJkWzm37BpvWjqFNB
20dSyWViTJGcB6eYxyc0E4J08FZN3IlnT4cROzNBZfxNyCRTWqFY7BSsPGvfHQVI
CL6yr/l3y3BX57Ap/bdpXglpTkmlxkjJn7rJ1LmIb3t0c0KSC1koIp2+hndxlOXp
oDsNrBAUFHcod/4e7MwLwHvFRK9PHIuYVA1LGf6AmgBybdQ7ZejeCj/Hl/B+WMgw
yuZrE1G2AfwYCSKcX3Zqr1z/jGeLeRS2LD73/QS1m8C9R/HEYW7mmAkCRFzAuBRi
P9naWUW+GCqusWiUmK1+DcE6y0Sf48wcZeOOcft/JKyX9V8j7n1RM36G9fr0Yn0j
iGWgv+Bt+W1PuLf5UYtoTyLBy7CO5/xJA+sei680QZvngoujDJe+Cn5zEqbdNqwr
ZOwvvMvstVCyh6GySKNvDBuZcOAdC2jA/A3pfs6z+c2rU97u1MrB+DVhlVBjQWcD
8/5AP4gVwdPuCdcyDafhHUqoDgbuZ4Vaf0kZqAtJUiEyFt0rPokwcTDZpz5LeaIf
D8OFSTlc3K6V8Sq7f6pcHWjMoB+WqZfuI2+ilBQeMWzR6DlRvnO9E22UghR/meca
VX63ePwBB6uwv92Phb/jpnPbs1VD7Y0yRkjTFem6Cx32eU4UZ0/0jmcFydU8SU7v
hUcF5Kdj6VDX0UTjoTkHtI9SyG90w2sLXxW4L3QK7JqpfG79fxfOrIFEUXArTUm4
HmaXqsGc/hA+ySrKVjiw/m8nQU3ufUjdCmCt2XHiLqvcaUw1lhNyny82J8D7tHfH
XBVt7rOudsEyz0EolrcLT0nnY2DKFFGjB0oSyC3b77DYcCa5TZhl2dxlM/UmkNZ4
hJMsBQE7SkG0zPlQOA8zA4nftdSqJYD3k2pVHpxoygu6GWl38yBwgCHNQ3wy2SOh
VLZuMzdcBlB6elcGYjXgHJBdZL99GxSmYuvAZWUi5Nb+OOnmPWOuzCgn++3R1z6T
kshRoKIwZfpp90HKAGVqeFlR5KrzxJtD1LNb9IL7ndTUJTybEDhaQDg2U9vtREuc
ezSMwYtes8awWyEV+O+vxQKO7ZdX4f/iKSOFhxFly1tJdscC1jfuMasjErdS1W5n
IreEHBFXGpn9H/kM7dDrVIreZ6iaQ6qrGOtEBiCfUUJWWijPurIg4VQ3NyMc9lPm
gXDu8V/hZMhLT6mpfjLudH95C/rhoihOiJ1Zw5Q21rytxpUKEJ+8l2HFqb8ACuyb
7Ppe/ULn+QQ3mTpLTth0500AICCF5V5JJ6CFOUJDYOS23rZqY4AgOOEWG8vDCpwK
cSflBG5bjEmL3XnB8WW75OUcZZ/BQCHQ4BE5NfxsLhCrJPnm2P2sQoY4dywBOtOR
i62TAOUM1i5QN4Vzti73lirquLtiMqT0SCBRtc2gjUueIp0f6N5XvAqblXRRR419
YfDI9Txe1NseJLFuJxmg3MbG9HNzClOhU48ilqUzQhM6XHR86SE5Jb7vWx9QJZi9
PvcEumonLrP6ZrWKXG6hhEW84cU40qqshktHiH1HXb0nNfs0DTJo3NbnGPOsbW2V
+cKQPnQvE9X3UIH6TPxMqhh+457hs7YNVdAOxiSLLdyRtqjvOgNXNPJybvEPvabJ
av5FqFuTQmrRvjnfm+Bc7O7IqGIyorSG7JLqZ4OQjljXSBFrmRX3HWSdVEKAoFuA
tMFyihv5ujV0EGJMriOTybZbuKMs8YQK9A918PN32crgTKRLejQmFLJ0Z305wc/M
3FLx5AJBjgTqiEkv3ATznLe2zJnWWh/pkN8ng6U0XbfwVW5jL9OpXUx4CMog2xd/
R/QAyKy+dsVzoVlSfc/DzlIgFUkfDvFVCiG+Zxr8GucNmRTt1p67QhjclHXCMonf
UJyoBib5VtTqLrDk9wkjREgI3y8uV1I3DrJXUbwq3ZAlToNVb9+34JEm74V9GUZ/
8chovacfXSQ8knigsY/6g2RwDUlEN0n7oQhQ/y5zp4r75aQ/kjO71CV193y8sxSx
Itp+IcQrM+3AyptXv559xK8Ejpt2NoGx4nCK6X0ssVbrSJQXqm4yVaB+fjB0Sf7W
/o9k6rn1DonzAaY9lrqC540zwp1ExvEcrWzagiOPX8zUwbgo56a7Kvd9CwJFYh1N
izl+EwkcZbmrFqYg3uLdGgrsliEpCGKWe692zmjs51xPI0GAcuOQYVCVReM2vSQV
ad9Ap2ukWmnd0ownbJZpofbmG6pzgG6BGk6YcNt/C7wo2Tc/a0hPrf1DssJiG4RX
gyg1/B5aPyIQYWrOJJkFCFCHP0uigtXt4tyN4giImMkYNZSePRC2CEjHudlUqyQi
KUyjdvRWgcGU/oHWZ0QAKg+ykNpsYjHanebow+CRs14W0A+Jb7JD8iDwK7kGVpuu
tWchCauocjV5qOY+l1vDRKMZ1iBGiDYIiG/ZrycBuIpYjOK8SpmxnjVHPqeMYy1d
vBpo51q/bX4/DiVmB3FQk5yJ3bMX5P18V7gcHVF+hsdViGsvdbw2Ruvir9fJTs3p
EgCGvwicyaEXIxiV5xZMrWwepAOrWKGpQTg5jxMQgYM7zG8hx8riFV8uY+VSO5az
ynEBFEp8f2EUVzkLFyS8rxfGeyB3StvuW86J2aa850PfcXWnaZxpiTRl9WrNDcsQ
0m2C7Evt8rB+bp1YudSybifIYoFBtSY91Vex+au5qw4W86CwBaFqGGMX037ftDMm
+umLDX+g4j045/9ri89Sg9v3k86FciyERCd0kV7if48eSVIjFadRmvM5Qdmllk1z
k5WmpqAz3BJfwUMd2DmYDARxwsF0wZBzAQREL+469fSnePwd1VUxeck3WJUvFsEG
N6rJxS78r8CauWpCVdRKPAZYr81vO0UO2zJMFHACA8vEnV9T27n6AFStto6JQM6Z
4AomW6jzXcpluGWPmG5digK8nGZbzrikwrmwAtXyJ2+V5oHgiPFVP1HcOGY95w19
jEU8qXvzyRtJ0SZelVyVzMZanEf0HkaxCS1AuFMBSqTJNND7cVmtEQFMhu3JEOyK
Hv7Kz9WJSsUPoYWRnCkT3TQOU86F0FhhVriV/qeDkcLxF3RVCHhfqpp+4cneRzTC
N5tWM8mDoEosklWCzBqAR63UNkzytKcgU7ARj0LeSGOdGh+LlEliSUu+yW3tPfyT
RxfH+NWz9oDyKH7ABpzJ5iU6jDJ24mbBAL/QVAXDaPKPkaQ8dakps4cqqrvcgmq9
NPujX9elNvTg3vk4XIILhhNct+W0OW0mdaaCnAKwhpBzoHqnn2vkCFiYf+n3T9vV
moCqSnBf17ZfdfBbZ7vLV5jZrjh2ogaZN7k/ZSDi3Ux+FhI7bkHmaHo9zEVuDgaT
UI6EAcVOrXLkX3+iZDIUi2rFwCs3o11DClJIYjoI0Pqoy2dPwqZhLfIOU4mL04I4
VlvkYvd/d3X+YjMCb7HikWAbAkwSRaqu1zc03gDISwu2EINHOBpNiVRO5HaRQHkD
vbRU8hf5w/w8dKO6YHd5sWuq180zyefNqM7a3GKD+G2YTRKaQKyI/gXKHrDD2tzR
bgqjQ2Vhsa/UeqaTLBHYm0epuYdvq1t7+6/412hCwEhs9WnlAxNDnCJ0G+sRnGt7
i0RcSsTE2dInkBNIB8FqbsBJemjVQXTnLMvOLCW9qROho5QDWMTKqFikh4QThKH6
otTe8jepDMrWR8B5x1Y/jjwtBVndeG035Zm2i0eGUnXWk9nTzI21rRLbkHhLqPFs
J4GXpv7WK2InDpZsnnFMOY9hISxOfvDAGUY7c8m0rO4Xqplxjoad2dmZ15TzpJFO
mgsABSFm/Cr9GHLOueGNOJmr4Z4HgLi3Tc7s7TT3Vemx5UgYSZbaTfLgLyv+GBvW
nAetIka+RYSFPO8TRqp5sN2BDmfBDQr7BXV0rzC9015KG3W0xCUee8J2AbPi0fN5
4+PGISqVKt0mFUSMfMBe5nNLDev8qYEXt2TIJcFr4ZOsFWk9hDYKgrnXzJOYFsvs
24Kpa3FvBwcOZmjtlCJOXF+l6RgrZKxD34E8+iYowUXwgwxvOljihjnG/ROO7dwc
pq6KEqPzBPSQbi1kgEqQZSjF053e0x+WPToRHM5vOtvzBhwmHC9e7RbqQPoMhSP9
cJxdUozJmPdaoIzKpqhM3Nd8AioKEfZyKmjGO0CEHarwXEFvby1lJHxZEx/S3eK/
EJY5Us3YpIbnchWhfajl7l4oMDh/c8b9iTE7QkIFEW9XFY1/UDyfzZW2ve6zi2al
HzbnVLImzo59rtaejqrCl5/Neay77J9x0lXVM2eo2cqUK87rI6tAEoSWFOVHLocV
/0qzTBqioGHcm+hn34ve4sABPvefA4zR9vO2CK0hhjB+EfQp4nJtkaIHgEtC+UnX
g7u8BvKhUH22T7g1EMLpaBioAOghKrCuGtUlpvNgrjMCkNb3ZY9qgfHo9myaUDK1
79fpQ91IWIdwTpkdfoEMgIZo4p4FQg1UePIVw2xo8PwzmtvFX4ui+4Nn1bazN8wu
K7usDOTk7y9js//QPeL2ebv0RxeEp6bhlxbND5KoRvqYvs9f62oMQFImAFn3dm8O
MAkkh/XnJ/wzwN7ynBcWzaBvgItwXIYK8EgxVnUB7pDVYoFPeykY52JbflcU/eKz
TdAk7SUr+89Kr87YS7qnXYoRmNc0ihaoj0U14I8gCsTQ6qjEuswApjsCdEdvCCi0
Yz+pvqG4OLcold4PL73vhFKk62M/oLfI4ls90u4SRnDx0CwINFp2Llj5RRPVAg8y
fsI1FN9tKrXKe/MDkHS1d1NuaiB+e185Auln7aAckN9rDQ3xOS1bpL2b6AyK9XUo
3ZLaRLPJu4GEWwqIKCkQZjuz8zdyzB32XxS7EbO/bO0ZTsLVRNJLqq2HIZJDGtLX
84026wOHjwafZN0yLT+0z/zD0RdvGhSZkX9Se501Ywre1F8lxu+f+JjHI2bHP37o
QRPuhgZd0j/m2rTetqLVC6TAyexZpp9vDzcG9DILPUNiN1UK7Kor1mAHYxhr2G+q
aVLk/VPMWfbB+xdWCj2InD8TSqbiuyH7liMMuwjCYQ86RvUDVms2+Lo3/r2reZeu
MhyTMPJzqXLZeZWGwKM8mQlgz7PHHzPKVow8lKBvCO1VieuC2KbF9fE6W4ewL6I0
S/tk2xZ6qhtU3+mke51R8W+Jus2qanz6EgJtm6gH37zv6vjdUUqwYHLbUzwCRDR7
SOnfT4t7NwEm4E7Mu1qXl5gRjBvHiAISF1davA/yGiCjZuu9tUxgbijuIkbVxL4c
wgSca0nZEXX+RaLDBkicD5RgSW1oRIiED/RjGY4pAeJNuAU/6u5larSwY705VYks
/d7Bv+BmJpIW7ncjWjZXdvDocUpgvnjkttjErEK7jeaqcCtI6+LGWQHR25F4dRmA
nVox5CKO/ZkH4hIIi+YM79mk2B6A6MLgy0Q1LK89Xv7/6czPY41VQt7tu42DaDH7
G8NMuTx00CJEltTNc7nJhr1VgzTc4WJ+BWh+lzYH1K25Q9zcvccJeq1o6GclfY2w
MO0OM1gNepT2iqg5GIAzRNM4NV2+YOe6ykJDAYXAvNeP4BhlZ8Lve/yrdmmSKI5W
L+1LgGUV+I8pnxwEiB13vmbcggHaxMZ3GXLqauWe+lElu50vY1UpDmcFc72/mfKY
EVreK6iBofU6S5IpXuhd3QEm88AZqtJmseGYfMcL0xFFJAK9760An6IjJ9l1188y
7f2swPpZMg3L5Om+POKUFFCPxC662MIoO11GYl8gexPEbNTeZ+xseC2eUFJ2hBCW
DFWyLMFEvv2zhHnubPflSMyQSu6E2DfsD2w39d5R877je7iFkKPe96hU2tDj9ina
HUyXRgaDVe1EVGpTIeBkm4LgoGCkneBJJsNY8xPfbyu9dbJBpOq2edlvkOhPnell
3k+JWimVYxJOVYMksY54iLQdhXxwwk+Ayl/SPay53hbK5+evhYr8hGG+DGFz8l/F
2QzriHeA+WKVPxFeFK2mgfJ7LC+HXjNvERPWBPIDn0nMhgVSejwYJYcjVmpzTGyF
qts1Jnf6KFkB4krgzPhIq2pILYUJSMUeCe2reEX9Z1gjm2YFeWB9ZWkzP4iOahLi
ayDK5hO2MtNe7qcOgh9IS+gavPzsPrp81hpG0u9JZmG4etD7GSYEntaMpo4j5VPk
spXxy+BJgp3rNaBuKbJX2pDINEy9Upv5kKyPWbpfSEUOfSBt5/pLx3pFKKJ3Xw9F
IFyafc1ScxZWOG5S1P1VENT/8hej67pivuwUL5uEm63i7EYHiFIjWdwvYV4t1Z9j
7aGGdTaASUUp6Cm6nTRLixhDPWcQrb70xjdhlKE1q82CpVtvxw6fWZvlf/AFDq1k
ZJmOPbTkuFbwojhU0Cqg9pF+z6kyDTW3a4jtDRaMwmrQPoNphZa2AUhoNIo8JTnv
Qjctl/I6y6z0uEweamFPIC9OFOnEYVIhadmMKEZu7Hv+W80gVqCEaPKzctOl112R
vresi8vplc+ZoDpvj71YO8+WXcgvZyPOGsrm6K5Wa5r3mBOLDpni7ot6vEoRJpgN
iMjfkV6/y95bilDbnOE+Pr2XyI8EFfJDWcJev7BrUXuWD9sSnrOgF4MPa6pMnAE1
PAjiuQ+G903KB1dBn6lN3SuWZhq38T+/k5nsPRxR4uGalCc9YUjseLN4w8WSR0ZG
l0oA3TWw6jUHWkfxdr5skmr8/tzY2CESj9q+A92GSUURhyZRwP+fc/rMOc4P1+ki
d129Uv4gu/YxD+ZdQCNLl1KR13pjRcPqt8lVx3FnpPvQR8VoNtPWcaiwKjBcuJGs
0zYQoTmASwa7CtGScW/8IxtY57nMlWFR1jpV2dFhV40iw4ymceIHFjdZSIubQmB6
j9/GItalZ2UOzJBnxxZETXY9M4DSgC9WGBzT+47QeoQ/LRq328jUCuKlQ3pshLL4
GWtTQ5eYfWr00UxHnp5kY7TwI7t+0vlpKAEym8nINspj3mcl3sBWhKUlIwvtHmrV
I1xFLVhK2cWBuP6RZMNlNU2vXjJQ2g3DNFj4xmtunwfmV55V+x0s/JjKFlDghaY9
r6enXvlrTfiaZPr2D/VL19baiyaGWK1D5r5d9ZHMjDKb/PeOVtJMBbidgEuLIIoM
euJmrTRsA9inAavHCRgZvy2cjI5c2hvv0sF27JPV1CkFHqPHmzv1OnL7SISLHv0h
Lkmz8rYj+2+Y0Z1mQhpWSUOCajxaKSqxZ+89JhmkrNoxpytCeNol5PSRoSdVXEF5
nJKCL147vj/TQb/bEorkWYEIttx8cqQaI9AdPXMmnDAW1iXcPEeKwaWvXNH8P1iE
6dvTbDFSdjdaLnQbRz49uTaxRmjkkwqdSxHqUR+F1t6IUVADZ5Ugwq0x2Do7vT4Z
MmaZVPZjI/bEI+3mrXdDjzCVaL0EPsnRkA3kyAoSEycRYD8I3wXsB7Z+jWgnqhXo
s8ghv3A7F9KPaKS5xH0Azl6uk7jf3t+vHEtJBSWbGgw7eQUdQHS60ZdM1UdySMCX
TvnObu8b0rFcZwTj2l9m1mHSPgjAXZf+pCFj7kIjxOm98vVekhGi+NCP3fwI/So/
3A2cKq3UfNVDy+WUiKnSnOI4YriLfgptKt40yFA4kG+hElgcl3teAdfSJf7oO0OC
WcylQPrasm9w5zb9k5GhFBaHdQKem8Ir27HLsEQ1AzkVn8A9eKjLbOqKKi1kyqQb
5OuOLnxmQBnhoUN2SL1eYKkk9OAdFAJcK1yMWHX+SjWbMduox4qvtgD36IquV5mb
7AjCoh9jvvOS04jcrG74w8jCKVnVtZMX2idv31yoHHh5uUU+9WRJdNxH/8PbZRAX
K+nZ/SoXghdx1yQQrXpuf43hX1m+6fk2X2EjHTPPTFeYDe7f23+tKVTVurbdxpjm
lT9S2V1onFAxIpo7bwa1gwgml9K2DfZfBvscG8BQA56ak0TSZHFibRheKK8z2J9b
mdr7p/4Ij+v5/M7HMdL+TtGLxtT226IcBIUqSTkYQGbS5Pl2YSYX3bV1wQcqzYtl
3cUl36FE9jz09kWBRVZbD5mznypmZ6cGs7an6gmco/m5NKZxXVQ+1QCckGSF0pBT
HAa2sG9HC25tFaaGvoKhKqO2rfUCk/bK1/gKsk5sy3UptpMOA/DNZXWdV4sUCg5C
Qe1sIgB8RXDH9lnrdEdAmkjfqppUX0LV5/jvs5Dc6cnQAt/ZYr1vy8WYgeQ54Kae
DRJg/6QyNMRCGLt4hgVYgqPFGCEYAAzf5H5eOGQFcZu8cJ/cVoOOYn198OGp4StY
2IRuTmOLZQEzEvrIiYo7VuFMsOvQWyxrXA+f8n44Mz9iBN4CrJTT1LEykPpv8Qeh
VWFUGgHE+qgqiiOyGncPahxg+R15J35QcTIjOMnwPy6c6lxzJs5o3ZLgmnVA4qCC
C7ipfrYNrXcbORjE4zMdGALOl3s8IgAqnp6L+/OKg/kQBXtBe83yxQua/UOex3Yt
rvmY2RKSDoqXOq9IkLwQGH9ogW4jtMs5iYMPwd6SoVkC6T9HAopL3FtVVwv6O3LB
nji2HCtdb57tHPt/py21P2sEU9bip1ZqEx2/U4F+RBSgmoLYFp6Xqr2s3mAij7CZ
np36jFzib7h3aUnt6IgcTswdyr3D+z36tZFO5630/qIvGCG0zDhxECeCKFltt2Bv
VHGPYvVcbmUSPTxy9AG8Lgd/toJax7ej24KwFZ62Q/EdTthzZ1A1XFaJp/pwwGmf
Gx1lA2D3L0Znx+YBP7XHPelA2qLpLpwA1sWJZ0KH6NBz2fQ/QlDRdtQ4IrDTi1nB
hG5HSiKUu8ivjATaPfGE4TKKxJZ9mZuLZ/OMjiPdXY3xL269LfmwsaxcMn900SHg
h6+H57VutLq2ZMUYdS9MPjojH9wpk/2kxqGsE3BjAfy8PXAU+eN+ZEBUy7laXhc+
6/Va4srNRP5n2FLQqNHn9W6cpDGxexPj9PUFqGt9sSBfv6amDKt6eQHCIjJFo1ND
jCbIbXIJcPWDiNwhsLTTzGHeFb2UgX0FPS0u/1zqaE8bjC8AKvXTigvY5x3Uz3XV
OmYcrtp3zR6eCbcSJ/9IlhI7A5dgX05bU80yktlxLjH5efqxxaHkafxGF+DED7Dp
tM4jKMdy/omnTmsUTaUho4Fw0jGFJzRdDo9mFyA922RIq/MxL8eRVR+PZseJDsVV
ballnqFkmsigBJSM6qgl/A502FHd66eY1ngExeBVZIe3IUwadPEU0hBxSUHxCt1E
oh8M8k3AKZ19u75p+GVmo2ovvhQIuY0xjy27PEdVaETTLVMhjDuaCCf7UZSnfsGb
pihmqOqSy8/R1Z6C0Ygosl7CWmsIva84HpG5iakY+kP0sWwa2+oITq4Rf9qW0ArD
qeuKOneFnKAJT1t1DsAa+Rj1USHdaXbj59i2GaWqLNN+okP/zsqRnehYcvFkFWec
a8Nr5STK72gZSdvVOwcCOw/iM0EdQPJSrSm7VKaW6qcPVduWguXiGx7AUnlARVnP
BR/WxWjVgrxdmhf+oC34KAmhgp6FqtKa+JEWzHU3MvHDdbzhgdOviuK3srf/l+mU
67X69dLvgmp+opcX0fHTsh1P5XIuOJuSrQnfZOMEv1547O95rsBihBbkA0p4eC9c
PAHA3R/xxV/86LAqS7j9YNIGAPAsabF5cn6jt9AYTjTwCJgU/5paw0LoD2eQBNGn
WNV6dHksyag97LnltLqfvNmFe+8oGwQyR8FUbc9HiUr9FWxKxHu4ZQqHdtjSRfkO
QvLgKA7hVgSDIg8f1E/nvxykm+CeXurX3f+e47CscKob9tEb4p15Tr/J3CBpEkEh
HWPWuV38iwHuS6Gu6LuPmzaAwReHjd1XZKQAQmzzr3iL4/Glp1gryTVcl6j51pko
dxjqln0eZufMsP1IauWjYA8x53JVsowurVv57k44Ghp2gaxfDvjpHjjZr92aCe4b
vq1s/EjK/EU6RZDJeJRjGcYYxCIWT1xOoF8y+xoJzKieKJGs3H5+CsooKtSs2WQY
085B1q9Q6rtmTmFcx1OljrfTFqGDpgAzrpXuMjuJPaxS8Kdcci7UdIIbftWvmYV/
YC8NowAZtWxfPms7thcBDICdQ9WlhtOv8DFWiauoYUIFtc97bv06OA36g5bkbgAF
Z1VLDUVZ3G8Skp33V2z8jQm/vNh520IIWidkecy+SWIneXDNqPONfda86b+quU7H
qfn/LYn62A9PDXdRJ2QKOc1WmBx0eOqMfDWNm8CQLhNTaWRsi931cQIarM9/T054
/IPFHyb2PC8MJdTaCK0NrAPhx+H7wkvOuT+fzlU5xrshqDEWwTYq7N2ZYvgsLypt
9zXrtB1q2g5mCvulw/4N7bTr0eLq/++NPAvOMNYtGfgO0I2N79FPJizzUmka0V46
DW0cdteTieHQ0FCYpkePcQohlbK8OwCWXCCF9kdOcuC1V5xSkHFEv2nvC94ve64/
qPbGbtnldSU3gsKTIMsIHZCIFxfww5VySPCoLt5cgX69WZUolSikV7Tdi3EifodZ
hWFch8fdUa2HQKVDAOITwDW5CWlDNuYMfrvND+CUHYVOXeMmyRPfSXO8f8m2+bd5
HOX/3/OwrNHnFBByF1Grq6HZf4cWRZWyOVdDjbRds3HesAeF167HaY+cuqgTOR2r
Q7ioQvrrwiBTRA7MIBKHKKveo6Si/vdlb/OJqzYY4dBbFbLdyglpgga5r41wbNfc
zpGUlnzHTDpTOMKWHanjDkfjN/ptS6BvYu4n7pei+xpOFUVAjr1/NRM8ee8i5B5e
h2slzSixz1bTVilmFCfNOyt24RK7558RZgcNVdxW5tsBMIscJvCXBIveKykdmkMn
Wz2quTzSa/IMP0rrnWFsCmR+OATmM0urMamJ6Ej3F58B8oOO2fJ7Mx2EKp6p7nD/
LOogH9ujhYNk4uWdr1AtPy4hS1aYQDZBo0RSuP76U2DYNsiTfKGRl1T/il3/0dT2
apHlT7aDOEd6BMFXskbWcGTL7LeO+PzaDkAmDrOhWYd57Qx2YKiQa6wWyk1QdaZT
CdNEBnPDwCUja5LFGA2iLuJXcvOnY4yMfy0Zldd+bBat3jKTWkWkg7OIVXSZ31Bx
ngzsSAX5L3kBpWeTsZ6tNHUnpcSomW3Ln9vUk1KPUEu5WA9bJCtF8x1D2meUB0Ny
fiMFdE0fUPnyI8AysI7FOBFtwn0vXwD01CZgQRd1ewJ8vBXYZ5YKQ7y51lC065Yz
1w+zhyCYJhH+z/FWcI0rgOu1BAPCLpKW3k5uvwgdZsW2jE0FrsELxsar62dV5Cu8
kghqmh/J1f50/oaX2TEF+2iwNhFUUrRli+0WUkWzhiYiEAq/FRxM3XrpSdp3HY52
PfAW1J+TJpUM/FaUpx/JaztOH2FiMPSVtV+VuBRi6qhH007s1AtyK8xgPQubuLFy
S6tgs59zUk5LO/X0Cu1GxNk7ua8f4/i8jVq/jCuBX+83Nfnv7TZExYaHOJ0xPNMd
+fo4eq7kNFFoOgaprg6WByEkSQIGSVEOZUgAN4D904enKFLZ5ZHxcAX+TCadvJyv
wr6eVrBp90NbNBFtxMbaok77OkDd8T1u9SFvxCesqtl9jQ3sgW0Xj+WNuVpC4X1j
1uySvY5jAcHbrFO/fPe0hXhkVg0d16+UPJrwqZMXsp7BOMyMCuILgCkAsV8bd77i
YFqydRAVxkSUsz9wKUksHLuxEM+HbhmuxF7scroh2wuCmHRnif51JoBk9Y2yHnqw
EhtNtd9avyNSLrZv8BuaRxlJq7fT68H8ft4Q0fDC+2icoyh7hKhZrpU0ddZwd0Aw
vTji2CDd5MDNL02iJ2SMsrayFMUpJddPCanvzdRW5pPgVhoylG/38kuHqPrRc4KH
OyBzBIXzf/v3s7xj1RSyopXRNgQ+9RvBXA7uELmYPQNspuxcx7MqVrM0eAtjNPNU
4GUCpW0X5vy3VMO2OFaQZeiq7goT+AdG6PUL9K+jSmxmF/puB+4FfxtrOq/h2dad
s9RWqNHAjys57plSQ7FMkfutZLUhy3ugqw1qlqmsJsvHdkkEj9V7++80nChZ8Qtu
mR3x6CbS9RuKp7joyaX+2nCm8P3MNl5v3Ti/cY3yvRoQ2fhLgvt220A7ZaI0rIxz
qmZ8fEXg/aga12YdPvPby1way6dI/6FXTXKZPa/6rVxtRfKLz3RGjgsW+WzCMGS7
ENXvmggIsj47+ubhZHk2Mb2fdkkW5oGLTdJkqQq52gxJTpLjt8ywxvWJJFBunF/c
7mmn+VUhf2x8u0Hj/DZOq+PTv7Qamev5yp3MCzZfe4MyEfHMDpzEWQN2RaAQSH8z
jbnBE/MK9139RsI992i0n9p1FogbYd3/GRJvvCSWXdDmxODb4UQfXLtw6zKBGSJ3
we56GdN6nqoGns8T/tPHXAsYiR2dVR+6Ulw7NWrYJzCsfiknSpo4MOwlKseCiVnP
wJwheGsTw9X8PuD19K1bTc3VoqhI5HTVeMKXDyIp5B0s22lY7lJ4i176OkVyTtjW
NoIR7W7TafK9sraWpPL9bGEBqboQPKjiCxE748Ibwjbre2VvD8vzXIOHezikeRqR
zELdamzxcj9S/nELWQtkShrHvxjCPNMlYvwUUvAIMHmYKCrxbfZ4z0CWXQyOAnQd
Ees7Utk4yP92afXQd0HhXo4E8h6sl/lI9I7nhPGqZlbwRy0KwghRnZhEYnowjpQL
xxwjN7/rDVFnGP9RbJqOSqgoyk4zSf8LPd0QhYRYTjuJiXzqdqP6ySlVQzQiiQg9
NaL2xnO1imuv7fJR/+jG9pq20CJ7tfqF/oRQYN7abnsDWvx9X2eRGeizq0LM0s/q
XxHHYcadqB1z/SeY5sczrfo9arHa7faYhb0TdaZZiY991n4CfpoMzpiEpva+grfA
LPspUpe/KdLuDqypQnAp1rp1c1pFG9oaHxH5GlzKs3fW6niHoTDKPsmFUXbmQjGB
tkTgjyJEjzRzz9ZTxC34Mh9TqQ4kxRHvAG7MjK4AhDXE2Ggln1wj9b/2d4jCcXPE
DDh/+Em8nIonH+0VbAB7tETIn9NkTL9osdiLL/lT45a1euVM+rE874aJfurfsJtb
LASaZUPk0jJoMFIxuhy4TklyUHTyohNE5lDHsAV1H5+WAExW36s62aoe9Soe0tXq
+nJph9nwdUmJW7LMnvxTMR82JwVAGAv377gCCyki2RIrDkUAc5j/fQrjd+xjinK5
NvZMqNuMuyRtRgiNeReyEGCqL4mDQmKw/MJSufPo/YeRdMHa4D4LUAbhowKq03Ak
Adevcv4+JSxqXzeqBLTK4YwInVKoijZhXHbif/IRt9OLnpXwHQgVdIzm5bajGfZr
ogZAUhpHx6/nalbky2BB+w6LX0P+5SpgQ0vQhdD+zZFBTA2EAWgMnEloNYRpHGwE
T5Xm4K0nnAzhYrszG/pUaStsdeIM2T2NyLylPh8RRshawZIbaIJQ6L4RbQmEbh9Z
rBGVZy1MEwC16+Np4N51aB++/cehBnJ8dml+QEhKPKpljuVXh6nHxwrYA7J5rYcc
Qcd9nuaxJJVhkdFV3qT2mPcNsR7cmd+xmbO2Pp23AdRcClIUKZ114yGzi20QWAbn
458RRSeRW5uB8HoxzUPA7GzeZC7TIPS78/zDKYXJL3rh21tcHEKpywvxiIqF06Qt
K5yU5dvf7sCENL3udRj0GwikOcPqoigs1ZE82Njf7YQlR8yVRCc2iH1XWftu6tLp
ezlC3CuKsNtXCMA2jjMvae1t3rwRgDcI7L/RL+vzbHPN82qWs+agX/+IMK4zK1dz
LE5ejQLW3ZsYCru/+UYQ2D6upuxW1e7cdW27Y5VhcXgnRnOQeA1ccoZ4aUBCYeOm
jGUAcS0DgSYkI2mEpJbYkVaqYswGU+3Czs435IDuZA+r8hPTRyH9h60/eSJPZ0lu
iUzETmZ42/DuT2SL4Zr4NM4XfnmVhyFZp4CmiAoYRDRDQQACVD91Toel+2L+mcFn
69PmL8EY9pNSh6ON9c5PjvMaaZ5u/eUDUS3yPlBtmfI21yBiE53P/sW9J4Zqpr5v
DMxr2ygMAM0WihL0EmIn5aUFuqBvxEh6TnW8XvDjTsD9pjBP+7qlLQS5wL8NGdPL
he8H30Y8HJcH4g8BMfySmCasuXo8qiHLO7L5dYSya6M9t4wOxLn3qQyk25K8H5nT
k2J+iJrpvhd2puawkgoGcI86TTD7ump7L/z2tZ2wJXKhobFr2w+IdjWwYxH1A/BV
3wY6GsJsvXq5/Y8RorkIc/rdQ+IbU3GIKtnrxXYIu3cU3vrvKsiB2DiEoqo5Fe2l
CunT9Rp2VJxAJzBhlkcmXHfZPQJVzPpOZcJ6zY3hgCDyhNa6lb+E/utQYKDK0MCJ
t4wa6g+Oh2N1KHAVqj6jGE7uu3kebSuvxHxq+QoFXmZwHRAHRbT1TQh+zig5uon/
x4r2EP7dya2v1u3eVlHqiWaR+QrGqCnvaAHoLeDf48Eijfls64A2aSLJXXvgjwU6
o2Cm1FUDB/7URXcx2xC0o3jBZGoqVNOnP2XV3Cphz79AZhYymwMejiZ8/2YjBMxd
bVZvFN714PPzYxqpz6/8cfjD+BledxeywbjuL9rKVK9yYefV86hhpTBpFLCVqsjs
w50XINfQh8pXH/xQ0753QPypO8sJZwtEltFC5flFLViSSzSYSewF0AnoSqlgmsgn
4XH172zPpa/x0RLYrlFmUhZ5cOnLe82BcrdsaqbKV1IX4Oqmt0mYDm7abrUhUPI3
RNEoLCQHv0QnsmXSIKJPkh4SHNdeiexs8SN4MAsJGyhbWeioNRRL3ocDY63/tP6+
5STenHsgAiQTI3fV6t0IGQW0/+Wa+jUB+NgBiSE1qz+p4cL9QrQh8Cmbr5R3FLIi
L3bVIAHpfRsWIvVT7BfVm2z6xMavLnEPvY3dsGhVlqll7oFmyPNYy3WmSV2kOoHq
meNygR92B8zUc7EDl1PHmi/TBQd6lK8prrIsnKdUVValXdIarrRa3kkTMqRoLWBM
xl15ayhs7gztUoGrdOduBiXoo0NsXxxdfekI3OUGLPNOzwFJPpk9DFuSCE7K6Q8p
QXmz150wquctiSFwaiAdFhiVZ9f9IqoO7vFM6Dz7VSr04w5C4GWhCeDqk3xjnrX0
Y/Uyeewhq2GBui1rx3SUK/QE0oNj+GZmkhUIpESpzpSR/uyN1739p4UfS6aXEFkV
dogYLV9QGC8lTRaucKc3Q1vhiXvaFeskcDBvYqdhP8iWlPvdWWKzk4NCaxCFvqbl
k5xLXi/A3Hk8GSg3kelD4tm5+kQCC8SOQQAJ2kFOZga6PyH0mAbB9mogce0kjD7E
n7Lj5sONO+ENjnRsylBRtoQzzgmNB+le65C5Lh8sy/UsQMcLvRGwd5bt2Ii3iCy4
ttg98got4PaLU5tbFb5reCNGQk4CZ2pEgbeQo7D+TRTIOBB18jvLiXTsq+4zAx1T
HRd+Azh8KijryfWzBr6eLS7lP+WxQMfq+VfdVwqn2+VR8awDvHTX/pR6ZRfqWumq
GTbYqOsD+FIKXbY/V7grYrVPVkyIUVyHj4NhKGQlsZchkJp+35jOc5wBD9uxAUPX
tApPNIHwCBn03s2f7ks08rCxsXSPhCONxYvaGZD766+NZ5/KRzTNGz3Ig5X8EVUz
Bb7kyDlaScDwX0gx9uogiTfeZJKrObK6uEici9q/w+XtIYkL+k1bwkX69zE0X9DM
Nqspq6cQl+mLgsxqjJeiAoK7H6NcIs3WmJiahrnIvnkGTG5k8DC/3AbGLLa/xxsO
OzoI+721jkmKEutdJpKzDcc4m0y7cle7RZFp9T0CqBoDFgIk20Ok6pUT0yyGCCZp
On64sdBzFDx7WF9EJUs/PHIZ0tDlb7fTE/w2O5CQQPZZSEBpA68kndqdsgeeBAZG
tHz7tGPL/eJheoA6N2Jpc/yB96QnYmYf25bWrk9J7LgjWCCmgEdEP0lrzradps5Y
XCMBui9zV+4Af8Oj3otGO+FxcC0Qgxp4Brq6QERe8c642E+w1HyvUXdfi/nP+lHg
rDywXxj7hFsEszC2vQVAzRekIAGqv4MhmV+AqNJB7ia34V8ZeWpBYqIVSulYc73Y
A4/iGgT+1iODBkVHZX+1k2eRRCBbUK1O96+WS/XxWZypMntFStEPQSYvSFERdAy7
7ijW9bCsmEKTd1XuFceIMQ3lKjaNnEQ3O4LU1ibtHb7kH6nzGj1gC4Q8aIjnx00B
jrDKCqokbWIgSR9hAYB42hH9t1kqg8hyceBd5/lL4qfhFacJzqhQDEY/+n0Yiohe
68Ui0qKdRUofUV2zz8+PboN90LVEB7q3mYtjJ1k6LUjwPLGnze/OjjPDR4O4Mnem
NtGlaudns2QYZE/Slout52082bE04w0RgzeMMaja3/r1JgIlxBpWBaw7AsKakt4x
81raQZwn3gWejXO4eHcz9AiN4Kv/+ZgSwuSi8fiHEhyMoGRSu4hv9RLq8q/fdEpb
/7dreEIIXsfpVZOGacKuu23a3ymn4btfTzd8T5CJm3UbN/snGMKOxvjqTncEE+cS
Jzy5W2I8vAy1Hf13eKemtyVsrF7jis9BTzq9X31d39XW9znOW9JfH8gvV7um3oU/
H7H2eybJ1NKFDArNVVqWYQ3Xo/K7LGssVOq+mB7ATuRIGWtK41/qQ6ljW5XDhFPz
SqoIrXOUvM0VkrRwHNA6Knc7vTOgPnR06iVG/HZurv2759lvQMBl4MwimP+FVcSn
NgoMexpcbKDiI0TVZ7/r4UPEzoHlf8aBTi0jzWnuU3Ba2kquh/daOD6eBBdPFUzi
fKy1DjR6KFYyAmsMn0cWFpTOetioMyEkbLSXQZDjTpNxuAWdAKkK99p4ZPHOWEsl
BH34I9giFQt3iUbJuzjqg1EFAtupx15k8O5UACtjLuvUWYgRu3yx6pKg+j8vGYCq
zoEFZUEHkWDLBXMFvTq0amwPBNh9eFimT2+YPy9Is3X1K5YBL2/OsXYw/YRwaoKw
8ikE2UT1isphtRnPrhsT73iymEjpU2fsI8blKn7i4+gWPjbGaA34IyhipNfBR2I2
aLXNQ4B2MeV5UPdeYisfhv6aa2r/zMikcuYH/wUc9HdKubH5+4QkuDdJ35qLLFri
aD2PqNXGv0IbJuBwDr3867y2onJ6USUy2GpUCWBTIxd6b5421Ep0njoZsMzvHbAE
NyPTStJ+zPGr55HdUGevwnuiByqVocOR9Zd6Hiv536T1Sisktu/R6YpHr19GQ7F2
zL5sWERfP3Zwj1XtaeiKGaztyp4Rihvyac7dY/E1ri8Z7GJGq3x6yycM/B4R86lT
OrN2I+BCckKix/TeirweX8tDlb5gFabZoUMNb9j6mg/rEMPnRQnyCPYDNw+V7Fug
BqEYM0vhHQAa9Qg1WTT2gu+d8jR+78SqUCoAv1/yV+XSJtG60OYk7mVAw1FZ+Apj
pOL2BB0KEPb7/YYq8+/GcF/Ukt9lLoyxOlCtZYxB5OsqZLialKO8NrXda2EkGMUF
+ENOhGRZwHmRMprMrzmCslR7IUTfpNF1XiJ+U1c9SBLCWWWMuGLQ+twiX4bOyTgF
EXXGJ3rNUR0RnCp7bkRWAg52GMoJ0iWP9UFNWGNBL6M4hKxhPI4bmnN29Dw1rgQ4
lOhTEZIR664tkn+28GnD0NTzlXFVSWwZjA32mUKo7KW2vObScqGCnjZ10GFdMTTE
Ih61dEziE3pJ0+VrO++dYjcyPpi9s7mEOp9rPO/qHQZLPm9iY7hAM8AK5vdP+oV9
IhjianEc8wKQbcZcadqgcKhYCQL8u+poXyvKwivdSleHVXLVzFAGet4pp38AT75p
VYEddinq+EKn29BYOJ6waSUedHihSdPhega/HevKKkyirhAmQNUNgs/LGjYBA6uX
tuOcNOfkh1LLkWzqMi7ldIl2mjHaHLfOEp9+RgweMoPICL2qVs3cYaQtXfZ5b16a
XEagQUaaRtVfjA0CGOCP+N6odm9H8NZSz+8owUvdGNsz5yRfIWBYBoZ1DtyTjtkR
EbAzCLcy7XiZNI+OSHncWcefgzCT9E8cagRR1If4JCzZoXm56Hfogh13Ob5ILvR5
gWHqqtv++iVFriRPI7I3w0NJgbhRLyCjT2lmY72klNVK3XPyxLWL2rlpis7ocRDK
rO/079diB8gvUNDPPnEtknN/nWT3O0UeLEyPeWdy/CzBOlDm7OXwV+zxjFm4LYOK
xRImmuC6Um3GxYh1yu2yXYNjUCFl3P8ZOfsYp6s7CyMw71c1gFWt0EmD5pp+5XWr
OAEKcUNuxZu74XRx/QiSSG38/jlicrQuI0YH4XLtBzWypFXMb5zz0ETr/JK6E/oo
q+0EyHOHTu4zhStYaBriFf3fok+bQlNDeqp0jM/Shft7fVP5TPifw4otF+zJu2Mm
fr5zuk7DTBsFOKyb70gJNrruzpj5CbcRz9TIHpOXwJjA6MPsYsaJia7SBw0kS91I
J4/0C/hW9DCPVVoAGGxsYdPTYyObCiFrgNbc71iR8/MNQjdu2VbxvQjWKmg1SQGD
qC0OOVK7g/RGabTcESLOctUxbfBUlfg56wGELKI5orua2Vtwc3SQLsBPPbzpgjMV
Iqaml4p0mlaFb+uj31XREDxtklwswlGUea3RpHlPWUyL/t3fV0wIJ5mHhW05rlft
PDOthCIyStLRCrMdllXZERR4cCKMcDKAI378F/bB1dIdqgCV73VCD3qFl2A33y5A
0AQoDJiH+Me9Kba0Ye/W+lhxX8c+UxOanzfRwFjwMx1fS2/tkFnELQhQFw/+MKzD
w0DKEcAMREwlet3Lzj3U/EFJC33CipEY0qjZg5De2qCyELRvMASgnHhYZDPS19N6
xQykjhDxPSQ24pFpYgN2V/8yl3Ce8AZEkFMHW7RNoIV9aHZBOTYGjO5N765e9u0K
frP2/0he9C4yLTweDJ9DkfedoZpCFgycnNZWeeb3Au2GgslBztXjtu+fos7fyZcJ
OPiYN9XHq15AJEBTZwwaS1zax8ff6p6JJD3MMTBZbbtZF3Dw8QsCkVKp6tkhMGCN
Ngl7wV/QjYbR/gqPK4bSpOnaasXovnAF4jsqu4LIcFT/VchjZJNU54nkyPVZAKAy
4vcRD/rAE6FMa7VlSHoaGoNxC3hT4U5+6lbq/s8StuSFypuRdR6Dl7Th/c4DWLgj
0+dLIK+0eCMZm0KUp1VPjH8Of9vxaP669Bn4ssWr2PMLnBzGxamH32pNwQEav4Ko
YYEjuCVRlDS79ghr5aKEOkF76NEL9hZldRC3+iPul/+ttKzzppgd+/Kp6NPW8bAQ
h61XTIjyofsLLF9kYA+FgyRrIKaUARSvIEzWXuMLErIzHfvEsLwY5cl19uWvUvlz
1QTokxGrJNUA/SifzI2c4jxsmcnxDbloozghiYnAnul5WDw2Oe0sNq+lNu8NDUeq
bsJK9cCx1j0kEdiBT6bN0Rc1GqqbaRTaeFTIdcPWoiLN7SBnj5dLvKNQWBuGsaSU
K6Zud+RHzuHEpDLdxlbpKoclIkWoIO1PhGZrqt6GHZt5yUvuu3Bwe5JQGlhqXKE0
7ql8C0oaNUZQo+JGB88fZrKvf+nCnpyZm6Wucx5hoeLsLy8NK4NfkKOyoLMXrNsH
M97IGefNdV1DEB3J/JYD2Dv6XKyjDfnQL1VODi04b7bh80qZtGi8zgu5hYE7POu8
+FscEFphCb1kHpoOQc0ey8c3XUH5akqGbLgdczSJhIN4f4GNSy0aZJ/PCDmNwEGH
z1vZhHxrsZuaB5BG55w0lRE3EwliaIGLRHlUpnlb1gUXwF691E9B2uTBTUA9BDUq
GHs3YEsg1VeZhqHnF0WTO/5f57v5+cqhMnmnADy9P9ETdn6h1qrnSiuZl/QS8yPX
Q0AWaNw6gGOqc5uVGrYlt5bDx63AUtEeZzYITfDmxUa28awrNMennDfyaab0heuL
RGr58Xc2174R6jDK9BI4nb8xFT1QnjeZM/uD1FKpKUPakvotUzYEL5CSkh2eyLEM
EVh5XTPNbnsRjHRJsb9cdQPMDJttX+vJDueMuUwd5IbC34fy4RN8ta7b8YYH5f7Q
oD8Qp7LBpVdfkLwb4eJ2lfqIBb+IkRY1VBFHkNxUNadyCRl6Rm2qvo4Ab4CVdYvJ
bNRJS3t9BRJCbgOr4vRSK1ouFTjsBZKuxPqdS4/PrUJgk7HQHuI8BY4uJib51Vvb
0BmutFrnEGv5AUktj3tCFkHxQgkXhUKVD9VUgJh77OJqTrYNlZ3S7lx+JP4jyrjf
jkMpCGZgMXOmlO/ADwoOFyVy8ozH71Onouv+lyuRrcNlr7UbgH/fj/x/xpse708F
t2uSaDYKu+JLDO2BnX/vJIWBJ/1cmE86memsyxxvITVsb1X43fAmTRm2qy2yubqJ
fjBhsK32YoHxY/5ISglsRYc+wg2qoZB4wr2HuqO4QvTkKISt5Xb6AeA+y1HcfbkC
s7KRTGFQKVKYF5jOBTD/JpqwrrZ5g9Yo1mCZVk9V63N6RyhoYann3hkbI8Vyl7oM
1HaYMfiV7UmzSIGzoXHgjukrzU+2VRnLu+nETywtWCa1oAm6NJVGuzKfvzuT7Cxc
libWnAY30lMp4m3bwfT4M/ecud0FTkReyhnh+J5zlpgY+oZ1jYbaqm9kFm1bhrWY
BzXc2iYxhOpNIuun1XSkH7nrMMb/F8pYg6WSLyU9ovd0i6JmoXs3rSUe8vxj+Oh3
ke7Y02c8X44DVCjZz1Kaf9dltuHihBwhG/LhBDqcRXMOu1QkbebcQZxAhpCGxbNQ
PoUwcmsIP+sJZKQ7KcRXvMx0VNVNpOZHrS3Iz6cuO/S9dqGqtOhopbpR1ZUqpuI5
vMOJAWGNAVlhSsut255HqJSYFL3w+mhbf6qRYmY7eBbzJL/bFIr5FQiT0SuUAzMX
p3k/lhjKS81AoMSPtexlq1HZpNKqSZ2I79x3syZJnb+cGoZxpakj1qImQn6nHwot
x9R3l+hhxjXI80hlqfeG2F11mib9rFBHGohKYHP6OzUy5NT5o5SDWAAX49JHBPvi
MSosVQWhARE12smlxU3SJ98z84nevBGSDEZrg0qr9hvVRxf1s8a9VWkBdRCb2gUH
Sh0gCJXgqfyGFs4vuM4XGjtRBt//4RfSQccSYF8pGCMjS5p6Ks7S+SOFhhqOgVm1
0SAXDPYRO9vRSc1tHLQDXgmBZx4p0XAwXeH9ouLCaCN55Yf4VajWPl1RJwIejZFV
h5Qg6wO4gJFNp+75hhmK5ZCLwFxtnAnQgma21iB8lJWL4r91fSREddkWbYhigb26
LKpTzS/hMcYrAsTEEHDH9JXICS39/rouxGKrF2S748nBAfgR2qBPc1XwdVEH/a7P
yQiy0jI1aUJ9yi61IA+w9Ci654Gdm7xxOJupf3tHGtKT59ItsY/G56/T7HM0lqOq
/ds9D+KRTDD+Pb9nCpXEe4y7JQIS2U+A+Qwi2Wh5+MOmNr5xw/YMV3Ti5OgCWqo5
AqK2BWIWDMYD+XPNz0SiP+3eqj6qb77zyEogCWl3UPtWCEY7OvpqOt1KDLtNyAdA
WWyxdJ2UodDgA5eTn5Fx0Mzuk3CpcWYcbmqfdaYC0gGaw6oui0V7s0vicFsTX/1V
7KfIRD0JUuhgOPihdMkfhJl9OHNokzrNfqdmfeEK5PHOf6tWM+SooyBD+oGcHzlc
lL7g6JOV4fwoL7tlNnJSFc8fx0NmCYuiXiQjpxdmKq7U3dDQsEdcz41Fqlktm+4A
Lr/+joCCsaeVcKJe5F1gvaZhn2S24WMjKUrLKcgvMZq89+/RveZmzjTYiVA/XxG4
zaG7BG16PiEfM4H4yPLeADHU/EDHsdKC8tL9fFMc2/5//t1tBEvJ5YFjEIwHasTr
E+w34o9mkwBZ7Zi4HzIX1Jmp1HjqsAIDLL5JbtO30PSkNIss6U0D9dZCeDR2SIqN
yb2UWXFnS1NoyNOWV6KTZ2st0HhrTDLeBKVeTJj0Ec+b3RSGd5I9pds3O/l/wdoj
iy0tNmEeVv4pJMwhC9KHy3V8q9+nKFRj7zY3SUt0vO3B6uWhzyjoLfrmTTdgKgzh
bHuRGfbCPYzx1op1HYlwndwIPoF+CQ5A0b30YTc5GKRPODxoFCjQd7oPz6Lrrq98
pWvd5bIsIrWnOlKT/0fvCzHuhuPFtSZx+BtbYvkrX3w22NnrwQP9q+ANWYHs1KIo
M/1A6xwg+i6v+wlZhe7x5ZG2KTtmKvsx9Nuqnx0ObSdpOlKMb2DBG9x6QInekS8D
IFJCl4my8VCr4hQYcPXj0Ru9TNZr90+IIoQXQiUc+Tk8aF24eHaPlZFYpUBycknE
PNKoc2WiM5smfxlKtjoqelL4Xp8EL91iI1C4HFjPrxwdM41WP+R+WfYgGk23kvCM
veQYiGa9UKmwr87xgnSoXghO44EiiPM4bL/VQXVlgkzPbZY1RtQiLipZKoZ27EJP
fKOpoAmlh3Cj8ja+SXLKQVUSO0GmfbO9LILblgcyL2x5WysAN5frCmzQ9FQ51EHB
hwYWUNLL9bAMgmeJyLwMTml09auZys37WMOyEFuXjNWiSYj5lBcPJ70vu0cdndhe
mlT2QIAFqzh1Xgb/6ue6xOw7ZTbEeLVPYLJXAffqMK7q+oz1l98TkNy4PjGfIZS6
09oGsRfPyupIjmr4/3HyQIGi9IOwjetezfY50w9H5T3kkspyTh4EzXmsd1FKFGwA
vmIlBFG1t3X8X4Vvqz7LCp3LFzr8uFkO5uHUdl7+pMp0EQvCWUaZ4z0S9LSogeYb
w1PSQ99ffY//W+hGlkCdaYuYVdTFksXPX+p4KcLkBat1p9MRTXVQCX6M67zINF6U
r9PJ5rRoHZoBCbh5kj7GBZmfxXcMwiAz7PUw/jF725JNdUNsmRaE1hCYhnZokiOu
ubUdRJtT4OxH4CEuHyTeGG+opUxAoSWl/dg9p3XPj2mVDsJSqZgqOkWAT3T6Nr6k
keUTIwtBRrdRoOUym1LOA06iJsSH/QjgmePNKC865zQ0YN81us/aw2U3qJ401Vmi
lzbLwTdRSCREAfMRWRh1rpiC1l8S8OBdw+l+ja/dynZEolAKIEXBnpjoaEKTQCQ3
O7w3jh3Ad59gjdPpWEZeDX5EW75ivXDgD0OuwJP/gVNBi4J7b7uMJefmbpOVVS0p
QFnK89sWwp/epNEPIGHG6YC1If1D933TZgOKcJizUGcrzzaGeraMl9htbJTBuU6B
WvJPfLYYqLmcaDdkR5t8uShQW/huQoh7T6f0LDvQiXhqYPnN4n49Hd8Ti9Y5E6FX
bD2ecTISrv3cSZflSz8wx0HyUqblxMkAt892vWq8SG92iMyG3zQydhkI8m7Hv4pe
YxgTuBLgqCCptTLDXrWkoF2e27EGGyLle0E64LseeOrakRv56k3lyFO8KX8Gmp7A
EYVV2fuIm1Dn7q2EZvvOSga0CrjKmO119oqAz/jPnV86evC6wFSCV/vDnAnv+bLQ
B+FuGt8XtYxyiQ35PKArO9xXBAwcnMxwc6JO8XdK64hTwAs8bh1I1PD+KP4UjbnO
fpJsIN1+51vymhlNSQXlu/y6ObXU8wq1CotrivPlINHrR0Kci75gc0PmUE1qsC2y
SkZinn0TQOlRdky+VNx7VfjZGznBcwD5arDnd4NEtZ8RWvgXZh9Tr0eYER96XAsX
Wd/2k2a+HxMsVrzVP5bfcrtN8LZTFnivHEwrFxgMuOlDQq7xAlSAXwPgQ3YFlCtH
Sy4UN7qXwXEAQLuZ1sDO1QHPox/3YfVodNnRYq5alVQzD5AI9mFDnNor09BJtG2P
nmOUjbs5hUpP6fgzMvWDRAViNvieYiTj+u/HQxgiKcMxOKMpWGlxBhR5BOQZs53x
VBoAxAGTux6+sK32Wab9z2YwjPUbgbPG0KuuaUzYObM3pVWOACNladUoyY5rxMjQ
uZQUh+TuWNVhNvKJv3D/WZctJvKSQbLYJHFfS2h0w9H5cwtWWa7B6ljzowX0d1Fc
Nl6vgL0B2uw5rfV2MvyBB99A9wtc+Rq9DAAivEnzUBtcBBcwN6d2F2trrW7BhG32
Aw6cOPShc7HIDutguLqO87JMgjjbhgQi/MyziHdqnH5/2nakwzwzUefyPQ8jdH5k
BbNC+sTKdZHY5RI9GSFegqi5Kf3Y90E655hnZzwPbRmTOUKDNICUU49YHbBbTDym
UmpuuZDG7N7mzw7e6ovhCrB97e5srWH7jpNxo9DjkbtSZqNJXLJvOCa1mPCS/aHr
9PyJJ8zF18i+8so5BSpJt1y5UhFQDhaxLa5K97A0hBSLLjTN2lwu6QcLAjRPta8R
cMKN4n41yQtfs4xxqLNlhorpcYqMczUcBwoBbcqwBsf+aF+7tpnUWalDuv5+8BZt
R1DMHyKDwbvjrudPhf7YFkEFiXV8RLp0NdpSlacORjC1c6h8JmSF504+0OLktaeF
5E5VHZBbYZcIVFu9X66yPx4yoCHDIOD7i2qfsoKeYrgIxSfOJb4CmBSGcWP+nQuw
58/8L67l2Y+TYgtXfIN2wrcCbgqjPe3WoFPRpNpBxDqy4u4kkgX+xvEwy4Nu4xHt
sOS90Zc5MTSItZzOED5u3SAGRta4AHVGlspkZZA1nrbCxAW5J74qdby8uPdIkz/7
RFoRYD5ltyjkDTR60FARJSOaWKs87T/oESG3rQSo1y8fj7pFM+Qhy70/RgP5gGzm
KB8t/wpnn9OS3dWsLNd4gwcac1qJgGFl0r4mEotK6Rxyvy9ZHwXTu+cxIiR+lGGU
VAPCAGeKI5vxnpFQuCWi1BVMjM1q0zpEtMxixihiM/RS1bgXWaEtqVrfZM9hHswI
nCrMPlDmJEfuzof3zxtz7WZwqmFxL+GdX4tfigrRB3krRcxpj6k4QdShhqJQOxD0
AHu4cBVM9gOCATa1afP/Cs7mXgKx3pvkZAFTdjkGp86yif/+NrWMEbazkmD6VsML
8LT5dnRWtTzLJeg3DyfWQZ5OpnxOAzei0A+F/ZINyhDYepLYYII/VFGJL/hMOhH7
ZCFw8vDIFlhyMlhvfUdlscFMwv0ac9RTQ3sAftK0tBjnz97/6BCi0Plz1w0prCvk
gOQkUyloTZoF3l+4eiaW3ZP0ubvECKMggYaOwZ4FErFOYKaeO7YjjUuJKKqZOCyf
YQ3ZS8n2gjvRfHVH3couQeZQJ+xI/FACNyopjoX5lnEreLwTN8YH61lQDPXd6Hcb
Xbr2IrKpTZnG5yqg4RQEmAWJVOc6DwxX42rkQ4AZe4PZdZkFvTqNv2XxXLHba5Pw
32PWRFsredc9xnOKJIhPYKR5sxArVNTukCx8vD3fMyei5yz3LEyJfTKuQsxpNULc
dslGuB4VXftQN8qo3+VQwqGcYYlw9K7iAsI/MH6D1cA+LMsS2rfhQ+swSKZVOAjv
R1JosO5ed4ypwnmpXggK8Y/PtBDo+DDzdOehUYVJmGlenWVAbFG251pePYKAaEJi
yWMXhfPQYE4WCcYbHp9Dy8sFgoQgQXNHATj48YanllMkZq8Ss5/N60RDNN0VPe+x
MVi733ehwja7xcdELTISWcUeOyu/W9nEUA64rt074TcokuB6OINEG1/0mwcZfdAo
KC/WxeWcWVagnanp3vN/gJfZHOjLooLIXMbw2mQ4YOwu+msuaaUDjJG1UBks0SdM
P8kx9U2mXtA4jRpcS2rKj+Slf9+iAhT6JzTqMEfeLHyDuVqedYcAX9ENxVU/p5Rt
pjhPIBhJxu04GQhNFZgAQsyXeEAQZ/YzecI3GuiF6a4ppRvFh3WGU1twHrvWPEd6
FJ8yax3FTJBtjh9KfLuoGYMi01a+V4s2cpFQax0WWokkTmh1eMAFNN6fSJdPNrVQ
fyGEiBs5M6TeH+SQmfvfhbbW/skBEM9YRvg7dDOa6NHm7Bc3rke8uZcFTyWwWs0a
S0sQEKFboqrLEX51GKEFVf4PnD0v3d8G+ISHcJt+Z0LPog5iz/TZc3rgdxy0TSFk
Ss/udvfCjI2IDXf+OohAZuLa1KoJP584QBXGf7E1H+qLCY2EUyYRn6ukF3NfdD7O
zFBVh5a+86eqLROhSqBZGuCp2hYaONxnkuACUEqobMxxJKs3+cbISb21MCwxuUZw
E5xakQrtGnPtWEiGGfF9QfyP7AZzyeta9SYSAREizZ+k6j7A5KUy4ygcvDSvxPkY
fFMWooA0Lb7RoO4G0bArY0lxzxUFNC8R4COp6lBdQuy5hjaKW0XIu0E/UcbZ6Be/
1D8nnHbi+81wn3/XO8gZw5RJjvCOCIk4Vxxqi9eHNVInfw8UD2PUYuLcoRjupfGY
8ZAQ+A3+Vk0rjNwQgQePX5nRfYNPSH3LxVBWgBfrh5yxCB4M4DIyAehyiZ6NdT1p
CY7GCQ8BIc6hd0qPdEBmYZZIGZRZXv2KSuZ4kvaa23EsF9chZT3705lB5hYwK6uX
sK1sviWsvyudsykxpJC1EUZpy11zL2+OWG9e8eoeHknULnbkKNKs5Q5dkKxgS/g6
70qHIwB/rLmI/PcquKK8+LcGeQQw1u/yJbNiTGyUr1cWyHlnaiqJF8clC7l8aokr
76Uk6iUaUYxHp1gaaMtHDYDcdoNwEZaTibQcsHixLvcRHrJJebRerZ6hzFRww5gb
tZrbeZISZD3GBa452cV0iC7dbWGsx575uzs+wePooz1SQgKtgHixa5zy4XfWDzOC
tQCFuCOuueuMWB3uUc9X1zTqTa82oRt1yCCuJNpcIgqkbmQxLFZYSkJEVp/O0Ves
G8h9LJU0kW8ypEE07M5T5/uXLKDPJyPFpPguN+rpycITNTJLwaQXU7h6x7W93Yyt
Z98fk2bLP2fSwm083vh7JTjDHaS7yf4Nx5wBK27jxlPHdJYUIQPaiEiQhb201Agg
EbczQLUuB51e7obHilxGYwlMTTrQ56HBqqcTlqnknVHBRXG7w4wwZKEeu/UIYLF8
PYIffFfvpLql851qupW1jZXJFHQJXRh40psJQpUyM6cWpSYhnnlJk4ibIf87IWvd
z5J2bvDt2xW/JvEhormkKqgOCLEMdNrBPiYJVnGdsgKGr8o8cg1gAI9XI4Ayrnm7
x2jqKNptZAwd3emF64NbnqngSkKXbmTZ4qH4TUeUCfBsFepBxyyfb4Tve/hGh2WX
udcMWx9ubIj2RYdDe/rWtn284SCCKdF627ryuc4u33x1AwL7TAHPjieWu5Sawr+W
f761HSgTw8dkBfg3K6N4HntVwKb05cg7YUkluo2UTW/WsjmS2dTOtXbb+0mso4Js
2uoGaEbWmdPDjXU2ubfBhaL5y3vA89XbNX+jJyvDTMIwqMQe41rC7QuRfCKthLMh
cDBzUKYcVlYHQB1gJwQlT3bc+z7Bf19zf7Qowljmnv8JAmk/KsHpn0rDyq6YuQUn
/Rg9VB2/KK6mPKnQ5Q3xmdZYGpnmD/nMTaRu4AKMgtliLLVsD3WM6kPZ/bHdf5At
CVFl3xDISgSEMcFdM/tCHR8476HSGp+NGiQZj/ShxhlBLALV5vhRzfHI2MT0lgYp
rjxCGU5DvODQAO35ELvUBkcLwILHIcFt5761a3EqaTVlPOQjDwH6uw3Lkkd7AUen
MBOijc7s58D7a25HESd7SMvKdGAA7qw+VES79gLnB1zH2QGswduLv/TDdrTbHlMb
NNcJ9OGF7KOrURJV0cuot4v0vguxmgupYxrssiaVGF0hGyVf2OIcWHcMdCx7yZZw
KX0KumCAp3frlU+uHgGbYWublVT/g6ufiL8zkYw0g7Wjjdc6i2TIUj61rcqcq0rK
BmONFZQUYRIthaEPEXGJA67KgHXyhwLcTbxP9TwLURyoN+Ci0up5Bqbs2ob26tt0
X5kLQBuxNgBu1A6IwIXCAB9vorq47quMqj6iocDL2ImKoyMZCQz6n750nTYjE3zS
3msyWYA7rqGYvxG4eJyWw/x8LkaR9bd1aoe2s/lQMY3dGQwj4yLTfA7rv3B/H3UH
jn9isUN6Faxup9hlTU7lqvCfNVaMGHKdruXaQQFliIhxtWAL2a1HtUZhwtkV5y5V
7kxL6UGcNPbcnE63hGzu2YIJI1nBmMP+PexdpVT8AYPa9lWc08srTMkDgcKt+sDC
+6Nc4lCidFhX1bHtT90c55Xq5KHfCFzIWSksjc599bZRMCYKcItSis2SUqd8LfY0
fB30Iieo+AoCR2Z8rYTWdXtMQ3QcieS8NiU1sqrw6t/4+MMRuTtiThyN2mlDSJJW
AyX+C3FlA+gvKY4yPPePQUsHvHdkc4SBvTlMIYy9sF0JQScwpmXqBuUflxLNy6MH
Wut8Uz+XLchi1nJhzmnsgQVnV/lFjfLPI2jR+y82B/izwKF7f5NS2nnJkCe3t7Ba
Bi4OqTgDSJlpqMqCcPljHvlyK/wkPQmafoSAmU+fPOrjCvJbtThkTO+jTD4z7TxU
mJvtKIM/DnVlBGn+pLEmekhBBVEHiISfHu/6kkxgrlu7gDvG/yrqT9ZFcbCtLyd1
z43Q6gRl+9P96RbZHu4RYsEuI+Y7yyWrL8NfyOnYurqJyiIr5vlweXFBFCANGl8s
lcdFQZyHnH04o+E7q5y6reo/yqY6cQ6QrfdzYHGNemqLUv8XTDdknpU5lti3IdVZ
FnNGM40KORhrMJ2FcWSJm+whEEGjOcMd3ngE1t0tVwPS2+5Ho+wq3P0f9ZtbK0xd
YqOVnP6SnfEzeSsAAvV5WVyhDGSvSQEkQku4juIOIWRm3vJFE/r+V6UYaxLttuao
gpPhsPDfG7xW37LG7s14vIs5DD3qbFHnrvIAG4XaljZh2QD9t2M//27ofo+NAcoi
kGFlUw4s4G6o9fKzTeSa04jQMqeRCBIxIB0HT0kAZEg6XPJvvHlp1yStxdww6Zon
r2DC47W9c2UKflLS6GPSUbPndyUODkwIO9L4CwmF3fK87ui8fk2gyrOFrlxrSX/P
3+IuOPT9ppb/tkn9Qr3dzf3JegSm25l/6w6yXTGNZ3dU+oa13EnY4C8gHFwyz2l/
2fEWQAlNk9gkVXyw0UjGCAWyi75eMEMYzt1wm6EtahAM248nIdCDVzAcIY6GQ7uK
zJenJbXYOM4Rhzb30xxwgsa98yBZ7uc62d5gbhUx4ayG8Oh0sJTGCTmSnGLXNXuv
J5ZuTbVRzY76Sq0eXOdnNUi/TmBg0uyxQiDgz3U/ITQ5ZUkgxNujgNI4sdUPzQoR
Y10IKBog5l2d6tE4zYgrz2su04ZoR3jZS61N170RVqYlRYxbxL2kFU537rZfy8MD
uXcvQb8ZeOqH8mCF6K2Kxwh30hPxbIQvT9VxNTCEzhZoKlpvDkoNmgnG0yx68Ncj
hPtWYmFoiQitGhUKQSgW9TMzI3KhwH5w0eRu9kxH1MeT2CzH6RhuGjrnhA08YrZD
8wrvEB5n3Cm39QeEdzV/plv1wvHtppeBCz3OgAxpOKZxCUD0tCZH5GLP6ggO6TE2
erUiUP/0/LIHYwNHLAtC4U8LZt/T+UmFL9GeW5WkCRQb8efBMZS7uOy/y82tXjM8
c33QAE+NZiM5c2oQ92LmL4T3ai9eufd/peW9aX+eNnAx9QW0Sjjw8xVvC7juPmMk
o8sNWuckPI7A7Eis4MMw3dIcCAaxDp4qHwijvgCiokBkdYiqEGZrhEaTk95zlYbU
+CeH+kM8jPxabTk2iQEu2qYysd0NqIoLaAkPH8yT4Dv9tPdWdkYq2xZuI/ZX8H0M
MO4ypcfJuE02ogSjPshQlDOldS8nKqCXiQZ7TiYbPDRiH5PPFZ2KjvuiIJPQeaMk
YfluYmNv9EVdrwk1D4yCjXVzqC9QKoVd/wnYi0yOapZQJ4nqR/hXPI9P4fhGfE7G
Rm5b7SDCm3eLAGhbPi0U1cGpnQ44aCZa8+Hk7ghpxlbIhoC3U5ayWStUHRBiCYiu
EmIE90RtJDD2OEuzuyChI914sFyBmRZ9fxCuwdyH8HCDdE8TO64IRco7CnjXSMqR
Ymg34rMAvugWIpmLq4U4q81Z0GF/kLF68fywgBnyWslqFHkdejb8hTtlYqtQHEtW
JmlcBnOinUIDUBSYYyI3Rw6F0+z+yPNgUtuDyCesUUcT+M8OTBAeM7J3z5dvWiva
q42cQmQYvNv3h6WPkXPDYfFcH9rdMOhsNkaunln/M0H97OuAH2BxTh7sSpCdg/Ul
mO82TkrzNNt3EefJwfQApXV+af5GZx0izfeQoqSlw65nZwn0TTE/lLwe8bKZG+5W
LRcd3VxzAXxnSURu9bJQu/5C5odBCNaBba69vF5/wkK1qrJjFU1DmKe3YuMMQEab
crsAe2E7m1FDk+114em0cW6vLFdXIwDRosr4z8Fi6kD8TwEFfCyEjEZXFZg1oZQW
VEgb6yWZpLnFnyWdTMB1VCQMwh7VcWiwh2Zu4oAeu7t6w7X0BtDPkgr/BesjhDB8
3nCrbsHoBpIjOY7hhZ8EPfbgjTmA/3PEng16HV4jNt5m4uHKR0IZfAGT3ypwRhYj
qe4Jx021xPs7mwu0Fb5hfIJM0tUCYhBjDbfHhVVtueBLFLjANCm8HYkEBZhfGAoA
YG9LuFI7mSo6mZMCS9gY81vjYwU1Dm2OGDVxCOJsT79rjhdbxWwa1sHpXMwTW05k
cWbzHoj1/3+u72I/qF4VOXQY43EV1mrSPdONArn0AZAGbITP+8qVUhKin1tP1w9j
jddLdrru84dj5MSzchAXoA9/5TwWVaLsu1h2+W1ahry0rS9G6EujTUmsw9d0Mkm0
rsdfasRls/2RMjZRqbZyak4YM4CIMsKVOOyCIvgH5Yn+3nHHBhuMC7ubDaz8gw1L
531ukYRQcN3LocK0M2fYMZ3LPb79LkwAZ86eIirsbhUctYGcqYJHJw0TpmEmK9Hh
OQEvC08Msq3WiihwSq2Qf990WHjdSGrQjkGGLtIfsvP4KxH3yuaQdygnjkR44R7x
har12sM1K6bz0dtMXgi1VVuOEuLmyrdP80eq8ed/gyYlZV5ceP7gt/xsYGYtYP1u
iwQ5JYAhCX1PqR0f3QqVfQxt0qM/GwTSEpNNU7XfMJhLtm2QXGjTogPt7ry7AH2V
EHf1MwvOkvId1UOi9Mx/Lyc3FE25I6DObN2ow2UqEm/ztOKp+PUthQvGYMxQ1b+K
h/QTaznVsa+5Nql4zeGq8c2MAca1g4eNDhhe+kzHgX5JQt9tdLuHsNEC1HkeaZ6/
LWI1UkOUc90oHlgzGkVs2ykFjkudTXhtlPEDbd1SOZuu3bhW/wWBxfZHp49k8lmM
Hczvhe0VJQPcrL+lNT8nI9nYYl83bFJDt2VM3UbFoTGqmNLM7Uu4HZNYsFZcNzBH
6+OJfePwT4OQM42qc+8LweiZkyfuVlde6bMtHx0kYahXDc2O7xyKlx5Q8oWNuMsD
fFsmSBYez3wyLPvyHwPQqYhh7XJU4+SFBGIPYwV/iq9Rz0hLEXnoS1/hlxXc/13i
cx4e0IMpcNu+QqXXDeO79nVuqXi/ZUNWEKxFMoAdqd0QYjmOwTUcyvbv6zLcQEIG
NFU8bPs9sOsLIkJm2oEWwJIqzO2EUji8VFVmrh89FgGq2poff9g0MoDCi53uF+Tm
Mi+Lm7ydNgZSEc0t7SK1VExUfmqLbWB0wWSlUEYfZ1WSSHU9imd4J2g0aCsZ9YYj
39st0/QBkiUSBd3SZUE4P78KAUbmlDq+XPLBDJtwdNedoEJ2myME0sxbByiqO1dG
Nu+ZiCjFapyK6aBX8njAbdkWXAvgXDiJWhtxu/L2Usy0lBqRFdlmAJVxp0aL6kKX
R91PWF0qMxBOqB5Ux1w8UY+I1DvokKNMr/ypDsoO9v59kzTNQe1mSE2jVPqJDJzH
2/UXdv74ZRT62miE4WQp6zUV52D/eohjYmUt17XuEFepLrRaILBcEEyEkgrU0XCE
bEohhyn2/5hdXQ6+m0pzKdolmVUHowao1pZwsSZctcYcn/hI3gB8pLdWw4Ygk7wg
/QMz6r+VTfABNs3aMR85SSwMYHQgxZ2glvis/OsaP8ojlm7xj17Qf6c/pzR6AwXu
T6yHFEoQsw9NwRdoWgydG/+PQ1ILTSAzfvPufzvkTXKD4m2ZAp/ihrgmfWZNKvDU
caUovtoo76tykardZH9H6dJswbNKGy9SCuEZnT/qe04IYKIuOPr+gdJn3eB1sfsg
oLyiFdYg2k8RjBL+RAhgFiKZLHahi1my1tUZZkj6jZAo7VjPOw1vo4Hz7BJT5Wbc
xgTDPoode8EmviaHe1X+jSzriU6V3reI/ralaJtWNtE2zdCVMUk/WQy0FsQQYQw2
0PUUjL0IEk7fbXn0cV4fSwGlJ8mymEZBHHscDNSfo61EYBGH0VrdfXQj61lT85Zt
ohREuS5MlhpK7TkVw/cQP3VK7fCxVaIkSdhGhekiqpflQTyW2JAwsKjfYcRNIif0
YLK0uoPmPOTiMowYploQNaUgsI0J+tcj3BlCpkJcdnJzbJNv9IDbJ72NhIsGZw3I
kZcZAHuRDEd9uW6hSifmXVRVkIHXy8ig7O3Zb5/CEP5/47J1SVhPVFEjJHhh1qw9
P/oXCIdpmAelnzGMXqF4WF6QXdrgAGSPK88DkxsBW+6A2YtkU03J8b5CpHQyMA9K
rx/3gPR06Pj2KGYtGhWrcLbK15n5SoUqSyIe5EBUSpmjxcJFr558St3tV76KAm8/
+ftyBcwONLQqFo8urJGnteMlwxyqowU30XosgpqOg2zCiSEmhKRwSwG87T7WlYLg
jkaWwBlB0swfThj5cyHL6vfiiN1piknzJHNaIXkAdr38kSMhOVBOkzmiJO5w8yEf
R7AQculNqsHvkcDI697yM7Sa9QT2GB1QzafvrXifEIPFhPTeg6Rpq2sDbYpUbktM
PU9aIhKbALLNGLePyIUdGZISKbBqrrcDUiUik9BE1fUywTX5AOBSUk1QIoVdEpyB
2dkdxYNs4FNTL2g0MXowEXHqDbUGJKlZyMG10GkIPanclG6MSOyimTOmtQy61ezx
B0C0Kl/p/pseNOhhbu/GL5KrsdiiSBrKpQMxKfkW7KUpB34p1j+rvVkdoAuBMru3
OZhh3uPUs3zYSdWpxbM2WE1gN+dM7JiF3QWSR8l4flPgYOX9R6IvqtMa1xmJpVJ6
cfSwmNevv4Y7Te4JLNl3TXcJy1kvSoEFs5F6EY/PGm5fWXAj37n3WFQ0zXr0mzXx
Bqn8ounvJUBmARnN2mNizZGWsRvP6wD73PgGPrsmwAMXABiQzFue51uaV7zbr5Qo
lvsswke95eNYPV4Rirml+7H5fvV9HMXwdlyjnxfVHTubls6QpANuTh54++XRLgm0
2SQswRF3eii2e9eIgjPzHPLEjxXg8z1GAni9ob+tf0d1eqExunItHh/mzowtioL8
V8o+Cc4ohyttBgKHV4Tsftmf/KIHxBLiENSuAik6FR9h1RQKeGlxTP3PlilQRNsO
tRKf0VjLfVwLMeyXfAaa8doQ2SRPXL68NV4EugVN6BD+1oUkM9EvdlVumi8udOeF
HmxNHMJidKx6nNjziCLkmZieZ2AQudkuI5nPbB7eTLRZ/VEWQJW0YuEvZHhzTCUu
CoLiMHMcQq/zfLXHm/IxlMg9OEauz4Tc66x2O4gAvbyTaFqXgHtHMFTuR+8r++F2
SUjpEvjh6nlTK2RYGrvcnBbkqk8jqMA/mK9RxaoshJDsxtrYgpspoQrxlAlGmjVc
QiWb2FILcTXBcp8Afgw8j8Fbyt0bGt4eNT3O57ZWrgIaPhZCRKAIohjsPzDrY5kl
nSn23SirK9RFYVs8AYXFVcnIeXmHLkZn/Cq2m5jPe+6GQkKhnmB4dPMLq3Uv2/V8
CucPEXinAQEMeGBrYky+wZxWpxwU0yMj/YMYemDEVh0MOP3JyccYFv/7FLiPRNDL
XkzleeSwQ3YpIr/DtiPZ2w6H/DMhFxZb/nwqYScSvC3fhju9X+m5w77C1lTHvmWi
pX4c7E71xq13VCy2UGAHJs+cOjDum8nrftg/DVdUjB6HkbUu4DFKCQpylfeu7Lnl
bmeXR96e49GF546ngsjGl4O+GMNGLWP+3yga4b4IViQTNKZxGxHzCPQeJQJ1rWUZ
9cOZlIwKmaGjcInsAQb+C5Sv8Zlh+9gtNGv4ZDfl3JxBcJPa7NZR1dCJ85BaQmYM
ity05xuj74vTzZXmVEsuE+O2DeFBM8wsiT37RdQ216ZAJpbqerssVS/u+In6lh2H
/mty2zWkQL/3B3UpSooF8KByuUIS19oLDv7Ms/Vh8wGVkxA9iW/UE9hhgZ72Ml1p
aIoG1GGuZE/xTWkyVbWj2x9WoGWhubSVvwlyg/UQLOedV10nGAJB5iDHJ4hiLduL
vwbEMIbsxTeDjmagv8jWfyk0/DC+Nz/ftPu6b7fEytO/rYMqRNDe7Ib1DzfEeOP/
aUq6/m9V+rEGe/NgQYIctLsrCGrFu/JdLs9PHDQosz7ynO2bIDSDqBglHq+PHdxI
b5DRSRn3kVe2gu3BSCL0Bh6dXZugCEKCCKXy65G5rIG8biD4fmmTcJNwud1HuCUY
1PUg0L+S70TEPvhhXlZZFdHP3QIHBcirf5KXlkXSUPslMxzHeXpYGL/jX9V3fLma
T3o5v/YgFXvCdQG7LnIA5Pk0isnlsXs7QB38Uf+YynmTqotzNDJPDBE3G5CnxoZ5
6usSRNVVKx3vpslpAL68qlDrOBepGWUQbQHGi/lqpbdiH40GUb7Xj7fRkv2tZZdn
5isBHzIHzWwFbGJAFBG8bgqfwsZ1xnYyiZ5KkZMtsFmDd2JlcKeAMsMKMHCmnRAg
c66TebwNeNV8KdDIHeGa6fJA9swyQoKGqXvft8kfI9dY85P9JUibVmOpwKYXS3Pq
ik4PyXhEMWgmqsAjbcYzQDpOpGVlQsgDVu+hKiPUgC0URPxApTp5Gl8H8ZpaXvur
uvVTKnhMegMRImmHkzxiie9bJXx6irogvoVZhVHaTDdnBNXM1lJw+dAGrNZmJZVI
rjzCiL8k7deM0uDn2QiyHkt5XMqmiDl+SQgYcn8+emrL6bWmaza4mFoMuaeWBSZP
096V1xO5mT3UcTzETNqk2F3JbpInhSl5rzwsjqXj99NumOTPgmvKADu3OrJwUU9I
zq2AL1cFW1dgsCZFZj/Z3gTSRmm/hiz2H0mw8LlAd+/Pc7vYQb2Ko9h5bvzWr4jA
ty1VMsa7yob73tHdM3JYPqmB5hO/DojIe1vdGlJoWCreu1/ReeF9IFkGrTNW8ZtK
6PEPUzs/O7UPyR2bi938Cx3KlSzXNooo0JusDGibYf/avM0kEpkPHm8sl/L8xFVN
7kOJ2ldDgKiZZ1AxzWFJBkgkkordoAIq/Ig+0W/EXvC8PYEmR8XcWJhimh4c3fTX
0WN+WcVMg/d011Rj6QqjGuJstHvQcaj35mYoGe2M8B8klk/UeXqIWIojgnJ7pf6z
mLh+7r260XI/bEt4tXKcGHo2oDQUqg5bXGKmZVfX34RskYLfcvrGMo6YvSn/UlId
rSekoyBuXg1yN7yBOTGcO0sxYfb+k04fQnPAZJ3nIgrZeqX6ePokwkhKZd2fv4Bv
j4nopyE9QGxZZiUkaoKJN9GiGj4sJc15/y7Vh/BAaVzzl38ukJ87KcHMBMNd57+X
i/ytfIwSc8W2ArvIqMH40tC/LUJsc4J+plS/B835ZXv8aJ74dqhYqLwRbp2DByw8
XMNH6inCsVu3n55uCbMFR6k1+78EN/imhDYv+stoPudNeNmXZ6EBj478zhsbcDZo
QBdKFizEb7EPF1QiCBanzsSEmeaTskJbTYTzDWgPl6Zn4IwAk8jb8jCEdHllkc/W
jj/qUVUseTFGBmbSP6DOxd/q3ybjdWRkbhF2yIeoARqf3shLPNAFZniSieZAbTJf
wAV4xy2ef74QWTBW/QOpSDsJh6q0pgFGmYiee4m1OB8MshRUf+rpa6msCdqoqqKG
4+48zuSRM5H4TmsnktoJ3uTprs0+lDVL3c1EaUn9vxUMnR8bPmnxEofPPmHiDW2J
fYfQ3TLoNgbifVU/BrKN/YioPAFduEC8z+UL0NnyScYoxZRVRwdFi2Gjo1qk3YWP
EtACDdAmn4dadTWllrVWoac7P5dwQVKI/4L7w4rQ968GLVVjjP/Ea4bDs47XjZiP
PhRt9Ey80Jb1qFXYPDunpRBnxOm0p8HgLEhYhWZyx5L6Pt+uciPr1t8sR9tqhy/d
AVw+p4Z/QXYK6ChNtTeILMvtegmw5PCaLP/x8hhceIAQp4TL6x0cXbPYTkFSBMQz
qzcYacJ3TwJ4KjfJFLlvkS6p9TOiUBTeBJufjCSMmiZuxjm/uaNwwk2nCQd8Bv8S
rjJyIEYeC42mGiPf19M4qVu9ZFnUx/njMDQ13ELHVDpJTfNpgfROQ8V+s6oKv9yh
/3MVwaKELaT3S4LhLEdpOX1GTOSRo14ldgVGhnF4XJdsGoDq38EiEk/h16TQlm7i
qvz5dnD0cSkUy8/C++TMLSASmsrgP3Ip7RbX+W7CPHWybjvkFMOVk/75S2aBnVdP
8J9mC8Zl3w6XvG+UnwKoWdG1hVeo2uHKum3GZKd1mk3mvQNY/lvt1qeTdO2BoPzU
G7C7CJFQawZv9DfJtpCQNQv3W2eofXJ8Ood2/mtJWMUOaw5fmwU3j8xc+2CvuknO
ClxdqNOZ1AtsHn2iShAy/aqhi4p9Y+TGETK+vwCqhjASmUCh+fKxNRiuPqerERRQ
ZsPZELl5BIaArk2lhqClxkGD62mTwPE1yZrmTjffGE1HcVlZs2sUuTm4A0BjrESP
i9YqORR4J6Vr3ZcRYrmdkt4srKv5blykI5JOKMSrTjE+RxYoSZWYzP8yUKoOFoFY
SBTq6TF+5f4VP8OW8qGTB7lpULSNBFBgMfoH075aTyeX9CzpGYZ2YP3sZ7RnlQ5E
tbGZtSzVj1QfGbT3MEGHpS8t6BVI6Z/FIQZiSX9WORX3UsENqFEjuSQ5ZZtaCMlF
PpAidzfK/UdXOtw9NPSKH7dzxDrKY4Wm3PqR3qZvZFHaMJCW3NoPvK01ajXtEMti
z2Upcm82DaWQgD+KdaOhlGic7lFng8C1CR64Lnxkk8QbK1txVS5lzUNY1vMZBrZx
vyExCzMpapX/5xemrrHdKiprH7Y3ukJ1u+3x20hXSRHhGkx+DqK4vV8fzMuetFP/
qGK+v/ODA/tA/6HbbBgcEKXQHsMHJEO57iCQWFtIH9gAM8sZxVToGwyW9yVsS0x4
0jtww+FKTZp1zbh/vW60IeZ8+LhtkdwdTSXWyDwIcB8o1edNCCfYLk1LfMXHonP5
g8YVfGAvKld/6LnmSk42O2fAdNjEEaVr/AL9Hv4kXl3dPbXb/eJGymO5tmQGIgwR
oqOcAobEgrns+X2LlMfvfFLOkVbOm7FdwKPLwp/+PqdSCqAbANJqyAI83rzHAkbu
vjQIka7SYUb8YwX5g93hPdfzS2TFtLQH76mXp1NnTp9JZHCbxM+GijO+z6BatP9J
591vatFxohroGzjRjJkbiLnvJ/naP3WCC6prB46OMYVmNaU2xoQ0iGAePrQdr3Tz
JMYQQPF6IoNLYT53gD8kI6aoGE/jswvDb0ddwNjgcv0Xs7KDUxuNbu/m9ok1qPSm
W9ktUTzVZC/wsihav8qLs1B2F7HOiFxMACikrCy+/jC4mG/jjxllwIg/7aChRhZ5
BvXsI00Ot6ZBzSxEEc5ROuWPlD+R36auGsqx+PreKMkTP9kJv8JtZvLdthMQa7+o
7xQY42FtOcXzp/zMNumxOfwVPdHH0h8a5rNB/nAkwE13BH3dMZ0RbBY3MF5DqFD/
lDAql117AKcg/qlOhcCPW5uJoa6RS3cDtLVQFy9XO0J7x1wNuZYMAvjhh6/cPWGm
fihqIaTaxXnlAJJ7IaBXFunPl99vKFNbWWMZX3uW454t0Fv7knrc2PAcnNMJi9po
+EClIYoYmC4RS8RFaL2P744/wR4H+LNKuFPJ/VW+W5ATAn2cMm1VWo2Phwo05eSO
X1aFeD2KbGqX/U5VJzLLIlCM+dzR51TC0cmBJG+BHnnYt9Lk1Mxbx9yu5mY02vKK
kTasTBADMjKWUU1zRlWS0hHnVYsdlVwswJ+GVJYMqQLG/YMrM1/TQjg3DqZ6LnyE
9tBkmen4RPkYH6EyHpGkWOBbraxg1ab/AHRv6aOY63McC5hHW8yp/7kk0bqtshi6
qm+C6bsAZnIr/Cm+VFm9C+KnwYeKaG3wZOotl7472igk5cwvrav5Y1tBbvhiHE6O
RGKBFClEkziYT5W4IF/pMM8/Hvwy9DGeAqwtMOvN10tLN/hmER8abem6mL67H7pW
mjv9DjxhYvKSr/KyKY+dfWm3losppmAGz+UtI13KDZBfhGGi0r+2VOL40OSVHlLP
HaAzsZ+P3x5I6AvpZ2bXRSON7mjjMrHS4xtu9OnILV5dZHD8lQwM6/mXUF5etKzj
qqYjpmDSzlljymnPsf7Ie0rXWdHKe/Wsi2QeRCS6Lt+KVO1gQVcct87fin+DFk03
bYIA+wGDgCGQhPz8Nh1/dfBmYhyVeIZvl+5uQroWuTQmtBpsqz+89ziA8CkkWvgg
EmgzhatBMQ6PDXDRvhA6kxSUHH93muBnh8vnhd8Z+H3m1cKp+JXXtkf7EzoOXdp+
AcqapuyKY1cmXZW5CfWDe16QpzqJCgdOwBM2tMkVyAyOrNhvIrmIN1ptg5Q9B3e2
Y50e+BJ28ok2NF4U8PosWRcWo3EntzBagnWjZEy9lgehWaaRmX/+fhdU6Yw3hVQC
xTYIsBmVHN3Yh1Ylv8iDkY/HNfO/GliG6Wv8FDWyTXT5Ik7QflTdnsK1qIk/H6tQ
kDIE8WkNqgG8bt9R1bxAJ5v0YoWSe3P6pD8RxiNjx8iUDN3CGxfMIBw92GlH4lEm
7W3DFmveOXdgnxqU0oyhkPGM0Yc+97FJFjfUDxepH+2C/ENydBJtBW1tAjrUEx34
lN54sObrgBb/uPQ9gTDpeb0twPkcBlxsqsR55G/yRp1/HTOgivDcHO8pvWwisQmW
dy/wMzhs5Lm7nUSdriyrpNqUSgDlYtAwNHkKJao30gAUJ8PlHGojR7gteKhTfvJW
NXl8rF7Oj/owzVEnXJCZByDZWWrjKWzZmjlZF+9QVw+4yUdL+QV+6b/ZNkPvMp9l
htbFPcQga44JyJWdwht/h9sDETSsgjvtBTWZ6FentN+Oi0LgYinuswcyvrKPZ0LM
VCeBEipD6dLTPxFiYTbuTlryYS8XNm6NKbw2Yh8aXmx33m/IAXgHbpUWgcl86/HR
MYTeEdYhIXvnP8Bc1KR6DtHnfyrBJXWJzLwwEyeEkfL++y9JHR767IdI4d5mRHfz
3+Sb90lZLt3cJSqQpPxb12kyEwXyNkL8ncu4hpp6VPe2+sKvNGBTXfsxrB8wDggz
bIUgpNm7vNyF8/rrcTAKIMor2yCd56u1ewhpbqoglepYpaCKUPp5TkmUOFuzhzYf
qHl0mglwfkKQilYajiGtCbhOX1rrKiUgYXxJ0D65gpTM6Uwb7nnWlYAN36wEgy0D
qrAJ8fnBE+SK4thngkLOC2wR4g7YP6TqijfaoFi4arurwAiYw06p8u0p7zV9clS9
6yfhvpNvRPzT0azYHTPYLZ+mNDTszkhS8+8VzF+Y6wjmmdW4PxzQjpPbYabowIPf
V4iU2FR1YhJAC94c4MhuebN4FrLgjpulYSXezN8C5O1O2Q9+kjZqi6Rhwoa/JYQi
ppJLIFvQWh6LQQZjsMaK6taKQokuWgMODSbfhTswFg9E0CuUel9r2+kQgBEFPewY
NSPrf4bZH4OLkONBOf7MKGaHacOb3rwZNxiPNCQmfIdGcISqm8z4OVgkbobbEoXM
7PdB4/QgvkTgCC0sULyDeZnfjnKddw/mQTAFkUi2PJTfqZ7IrX2QD2UEg8JnbeE9
70mNN4tu2YUeiQQaqKPmoaq82n/owtyVtqfhlEw3Gq186wdJPkbBL+P+a3xvwDl4
tY/mz7mdSuykGEJY+IwrLy890QVJasIwouPbez4AYLGylofBVEiWypmg+zEvYKtv
nxEBo8Eja0Wtm0pdbd3DgAXJtgA25IOG5bOOSHTyKatN2yv5K4y+XSSV7M+HpWHX
He0yQJDh8IHIRPz4j3eISPxMKg+/3q33uoTY1nR0ZIYGeA657omzgzUAk87/Kwv2
rYSMQDJ7KgsX3JI748JNax6FZYOOd+s1gpj3RuhbgvDRuCCOdLfKnz6Cgy/Nf7+I
YVN4zJyayW696k+qUzk9WKOFIrwR8n+ze+Lzv7L7GUGRYx6nykzR+gv4Ba1bf8cF
LEQp3ZePhFmME4H/VQXIqR0i6dgc/PsEQ36R2gm9GD5KCxz2OhbmkrGdRXMGFjJR
yzn6r0tpePqUYdQxhM+v7JZpqzw/GAkFtTq+QnD5V1yuiJ/kE856iwO3WDHMTTsO
s23KaNKVZdCWg6v1iLaimwq+VVJoKeg/jbqOa9tnBSMIKWrCswnW05VQT6ddmrsw
6BlemLnn4CXyyeczGKYXpMigyoB4voULFnxXVzfMo4bH2flMtNK+PJzOryiPdO4a
wm0yF9+uCZwJeqywjjNVyBu8TFoo1c5RXobUR+FZE2QwQXIMFoDaGb1JOXp3G8CC
UPDYX+47Ll4trWpJT0tgmhjqPT42k1wZAEQNnbV1eUnVTUQS0LDbFL2Z5ckDDrTF
yZg+myudp5qGLcFw07VVIyA0pyqVBl5nj8Y0IGbvMqjn2w1/5SXDC/9VBNsTdriO
bXYBwLtaWTXovCLHXxo3xHZrPLSPZyAPMCJui39vZUUSGzWKSvLqRHeqtF70fLYA
22UavgGylsDplgfM6w4jgH8qxYeV2Y89ihpMO/o925wUrSZ4ylgqorqmRFWbGFu1
v1VPUvv/ofG4/GNkeFrDurYKovBhu/q6P9RlDAtH7IbXYfZn6CnoG1N0sdCx68AB
RpV7C26xiVY+vWF5oz3sNwzXHzYekXhq3BbyUcd5rWX28LrJAIWLpAq2Hq7TgsUR
I8XFgdwFWIq/Op1c2jT4eQkvz8CYP2jItxXT527uVX/dH6TKZwty1w4heN7TXJ2O
rWANyFj9fZ8phsSKGo1vR9pYJDDhZxczvuTQSlP0QBg6R2rIj16ncbqQjQd9rdW6
kWEGlqicntDtU3IkX0EN8fmM1tB8QKYS5vCy+mOOJJahUs/RAHqluVxsEqdQ5Ho8
DIQ9CgwZlOXhTgVydqyAQI2zpGhTdWF7jCM0aVis9idizzV9EALiHkdKpIcM2VSh
0w8USwuT2MiZY62l1XHKYbXCEZezFicviC7tPN3LTLUvPA2PEyIbItqPoQtcoBjj
+c6htaWAXNzwRRyn9Jhbq7J/A40DRQ47zAAnEms8bufTOhmd+CGoJZ0yEpO4Eo5e
x4GJfJU6Gdjj2H2F5KBP+uDyvRRPJJfxSQaPA/Psd9zXVSTemBL5eZkJBA6pOMD/
JWyjpFhFsMq9jmFtD1NltPS1UifLCEJ4G0sa2lP2p3UFX/qfgiZTse7XJKW3Z56b
WMfkVh6FPznw4OzT90AXL6kwn/3UpSAquuo91CAGC8E1FAsExt7wvMbjkOfN/IDj
B2Vlbu/zmvjfnCY96hzmmwEVnjRjYk6u3tl2gQ5OcX/LfTNpBOBwjHVYUNGHoukY
3b3ZPT7ODbmWrsq1mFJ9kLqqHp+FkrhdAAjvqgbQw6hP8MB/HcJ/r60tsipYB4w+
aqPZkNtEY4S4v+M3tIUgEdLStiSlbTTKe47WTaGPy1bzXd9//ZyKZKivl4piFnu1
xzRutu2ktCjfiXRmqEVqdhQRd+X7+HgpkAiFZUe9B9BB4X2Pm/j4BJ0qY5nnINAM
3jt3msOufggYvZZeJyjXXwM1LsQroj/n75jk7G6nl26zlFuBA5GIBsdU/8pHVi7U
lgnD1glfdigLK5iuPnKsMQXi3eVfDiyLNDeOkAjfE0yBkCtLcau6utz1/Uhi5gLA
1WjFZZnlb9eqEb0p2MygaUrK386Z7UcC8+G146gjgQDnqTgI2CQzKeCe6CgPWG+p
cJwdqL+0suPxgVZ1U/8tXoe9CRQHtMBmgUIJAUcdAOeBqLDZa/gkA/eatt0h2S0F
jaTFEYIQ1lqmyXWgsz9mS3feNrk1GO92ZuNU2982uO/GAxJdRlLwlj4DP5rXJPkp
Q/XWFuZ6qsviqisbZRmUO5AXELdPg9PL1Cjyza44rSwvtvRvb4fp1d3GkxSEo4Qm
YOuLatkUdKnAVfO0YLA5O0DIYD5nQF8TAVNLe8ezGBwog+lkNsBws4LHpe02FOlI
7GTS5MaS8k3Wok+AmbFy3zaSgByUxG+dO+Z1hlbFtwC+D2O/UJdkZBw87vb/cZh+
XFpHEdiiVAFYhvFUMuF/3HpRR9GLMbKhVw7KlYWuCSu7IuQ2lfhNvbmfQD9lPxxG
UCKwgKz3aLRbYIFWqFOEQZiYALw7ZzlGSvn0y3kdY0YhbF1ciosx4YDq4j49zzFG
BmGhbtLB2qgX0utyk8OMZERoVgz7LYWhEWTnYdVG9l+8gxgSf55eJGDnyWXS8oPG
52T2lJgxJl64S1CT+1XIiib+bGcZXyn0UeBrx0Q4zKSwrwQw3nmEtd4F1UtWwKR1
7SOb/+3lZzj3F0HzkUoF4tjyZfJbvh1GzjRs+adN7G0hE8SNre9ZHuK8j5lYM+AF
kvMwDIQINWo+86LlsESNwbrrl4J/+K+LLGDZ7ZZdWwCcMklix0G43z6tdoe7neKj
cF4Far3E1kixe4ZTzBmvqb3InxRF7+dmTYVQNZOzdykIWJiFpY7s30JjxgreFbpA
NH0W+RG95JnX919rHuGGHUk9I5o2ccjzHYaV6xKvtJ8kUuLy8Qo5m0WzCzQ+ysFl
vmZR5A9rEo3FKiXx4+op430wNXNZFZ4wB88ZzhAY9q8QsHfAIPDAXT3wyARLda/g
a4/r0DC9GDYl5LYxFu3LUn6fyOAbq5Zx11GI8n8lDXZRR8EeUSivWYIeC/Qq7njN
dyyp3n0duuwNm0oPQqcRHUkFJW+hKsqCUkE0B0Le3H82y1c1w90Mi5nbMKGzQN+D
9LDNMp6Kdrjb4ZwvtmhKZqFTovS1uF9yh0exp1SRm0bakSzsAV2lwytxmbq+DACA
OVJUjYTwb5vyeOobIY4R+j+u3uLj4JTxqCctmoOd482zOLD9ITyk7d8fo0OffEVr
D5ILtDzIPP+xMThwRBcrOvea5EIE7npNjV2t/4RJIo6DeGeOMmVCM/ibSv35yQhG
PZAT/KXsga9sAXrzHEsjy3cIdJIi6rrXfICjbSQg7nasjK9D+FHK6GPNu8TnOM2c
HqKdfLQLl7jh/0NnS2fHu2ogZCsOU6BYI6hpldIHhWUypMm8d0CSwdx8D57wMTJQ
hpw/epWysvZaggm3j8+zWHYpq/Sbf75vSHcKCiecP2LBqTGnxlPydqrqLUIOSJto
VH13Xsm4U7fbaAYjg8marBQr+C6jRZMcK+nB1N7kNnXMTmS0tIL2LvW5dmtzx3ha
2sbhr249szcyJawYrldxaP3CDHYoYsbrAz7DYfbRIEAz+JOsnSBu+PQS6478stqd
4mKQAJZ3G1jLJrKcnVGWlzPv8RP9DUjeZhcO3yckZV7JatXxOvh1cYsNyYrwnu3h
9lQzF+6hR3h59oD6v4QwP6U0lwJpAYzhdVkjKWDqeyg+AhJ5ks7AUhA2EbKApfO5
r3RzsB7WMrfJ7orugEPeWpV/7bXdN9rc6axKKS0p9RqPsOG7f7Q3V8tBrf3NHLeB
bo9KqBXPvSaBMdWpjq4x+y6ZY908qBqZTyhlIQucXxjNvYuICz+BEgNF68Whjc8j
mu8Pzf+DJqCj5RWPg4C+7ZZRHqicIuKqmJm2tMS8ffRJBkFzl6mKzyRQ3pkV3mIU
r6K/2Md8nMU+yKsZNA77aQzK84I/ykOE6GGxxtvp/xvZ3pDoqnDebcAxH6KaijLn
ccge/C2thS2229T5rzwsSUWlFm9N743dbAa4YD8R9wnCsaLYIJRqq4Rbj2AB+VzD
ql2T427DBfmnNU46TvRovgblYKA5r+lrTmXfYaol9RmP4dCF1g5hN3O86Vjwf1NS
kNbmFUmFvVq8XgxsnZ2QhzVYBS0VE3HB/1x3bS1JeEaXD4wkLz0OVoDVNkD8YIL4
xzHjdNZpLC0X86QA0QJgio/D0xA1g2d+HHJuP64JRrs6zdIeLFe/Jz0ojkzxEKRc
DtuAi64So6/uAO+pj6v6674F2UBQE/kULpQsVy9svKAulFZCqfYjg0s+eafpe1Nr
7Yo+lC2CWqbxfiDvMy8or1yI7kzybrYIu1VWGF1JK22prwPkIbpLcgfTKfvPIXNw
lYn/WqW1Oin1v5JOMeroDFUzLRjsHrvU6IaM+x9HSmFktC6GO/UhNC6doO+rpc94
8kjzh2elgggRFe3pp22hGpGIpVREnmTC33n/PWEC4MIrXzI5LUDCJdAPiIWqaDxQ
f6eMvE+AfD3EiZ3+CKxrfaGSYdiQyX78hWmCSf7mqfwDcVL7pJetzW2tlah5bEuo
VJ/9MeertcoOHmVMRptfq7lnn/CFmBXx3P5OwOyh2wPQP4xzoyuZ2nlqZ5Rj6Oxp
RuYuDB4g6GAZ4Mc5CryXrNV0Jjegi/gc9pnJTYxkGIXY4rv7asludOeln5f74AaJ
n+0umJwnxwScWy9Q6xihh9MFJbkyG3j1+J/C8J/SF5eOc2Ymd9wHVTps2SU4viCy
wUQWaSPnmBo9cFwx63DmP+ofkOSeYEp6nlzf4hzb0Exo75o+lpOnV+QYZeISDSpr
kTwpSrWqJpsZXwo8adV8mzSVF59oSqYLUphURe0dQ+nNB0nDKtE6JWr2EOFjY+oO
fbd4DNBKzTSMxArGO3Xo3z+Ri2oJipDEGh1awvfvYBO7jsUbKU3aIzDmh1B9IO/P
DjriNdSqJ5xW0qr6m+P6TLZSEdIGfwx3Rt74J4+LqvNCivyTzOdHPNOWX15xslt6
/NFyAHr2o7zRze8WNq4z3paG0K3IYYSEIEEcRbhN65TWIA7HM4n/hq9jSryeDrag
1z9C8RFEW3HgqtVimcVzsjG9DeqEWJgdFUwRnJBy2xpVJIAc1RNHcCPtij4QMIDI
j32rQ1yBMAVKzT/q1z7Np4AtC3ACX6BsJIOf13QkhEA3cXz/6QX8S+JCcyO/j0yb
0pBINqR+1VkyGCXdMa1No2kIJztgr3+XdzSOA7rGAoh5BlgwvTQ8p5ZXGxLdwg7K
et/zFlnaJGJjXjIt9MY/IrsYFqtYHr8VQ1l75CFeW/sXltGPdhfcOkMI/RQy0v/Q
/IcGU7vQjnXjWUc0HVtEdEOqH7HM5Yy/kTbxNZDBabJ3MNbCTy3aR4TD6ijfTTu6
f6v75WoT4SXw7PHoTejIvPQzlutOGsK8sL9G/8PMo0s8Jz10hni0lm0M4ky2TnrH
5cIS1HWGfF4gJ6+oq8TS6BLexCWyBmYTUwCxSuibVbMJavuEiPg3JfO4/wtP7ngr
T6sfNr9p1r7lYEe5jpFHKKnpqM9il2lJ5eXNZMgk4Ye2+z9PB1/wWCMT6Lnu2l2L
4XkxvEgX+9IGEYW12S7EhCLA9Ya+R/bJgHI0Gg5vJ3ZUnngJBgO1LhQoDpxSy2P0
0oja4EoS63N8tGiU27Sg69SMhePyF9umgUf46kV5ANzOFM80F/Q/kH9aNJccwM31
XroQI4ALzH6kFGFqYVqGdcd9T3r1qjmF6j1AaqIXWB2bmeWqjO2zNF6F3Uu6oWUI
rDnFgbwjnjBlX/Tjp2LuuvMJJSTNflzyurCSIWErQvI1N7QxcaQe01DcZXyIzHtJ
Fdn6+Ph5MrVUMnSu7B++a27nJvspwoh4fSHHO8t4lCJvqaDHrExcgYaNxb82fdOI
jk59b8Lj1cWGqYP7oUe/EySLVwbYeGQJPn69KFjqxh5dBj+fDxCNCShyzxUgNtVy
nn6jfXAcKifx8PHkAINKE85gWPwsXWOVsu9xz9TF4/2wpE5WhTn1fp4WBz1d/8rB
ErpzyM46h85aY0QJ6eLzguxsfpQf2+R6/yvNAxdVVxNGSfhATQA0iSxVErI2JJwB
PBUMJpu7lC74YJbhW2KRZAC4R+umgxzzyCRyPM7eFbscpc82EkPmUVsbDs7Quxnq
CnbUINqV+lsUUqzOsBPzh1xn+PF2Yd++WVUVD1QS7mM4Aj+/aNMOtQPm/6SbdcGW
yD0mg2M3bCYuoLQbZO37M22v9Sf+H/TAUhabFNpg4HBtIScftLEtcrb8RWqB+Gsb
zO8EbLlXPCZwSEJew/r+1i0NLU0CM879HyOTDKsQD07zmXTNjnE/PbwjmqVAUk90
KClzJGiy/J/zvVmKqGT7AfFPO13mt85NxPzK8/p8YXFe1Q7vqMzQUJQYpy48jAkS
DLf9/sAwd/Vthnw6XFkp6v6VmTjFx/AKYFWvcQKgtZumvbJPtAqAnv0foNIGVtmU
yTwWm5JE0+I0ItWF86Ul/2BRS3/ovy7xr8RjiQz6pecimYuwnfty6zepjZgPEbH+
lUMFhZ5+7INbX09nH6Mow7AhlTH8xOxcuRwRLNAHXYn9LgDEf/VdedFJuJAZjxNr
/R6wU95zp5Q2ysLaELF4S5ryvl17M0d8x+IMLH3f7xkXm8zHRzYT0VEKwqWifKkC
aVFuTZGOBZugbXEBNQGEp+twoOdz4SmXVjg5mh7t0FlLO+y0PMJnTwdyzizt7xW1
IsvCkD/FImQod2Joo8imab2idss3qkky4CGFFjpXH4Ptqe+2NVs2DpM1/Ho7vK5W
gTtqXEEdUFX8G8tRbKsybkVJg0WqLGMhSHR3fJPIwaNw47iQAEBUGIiYTMotZ6Ui
k+8NU2OzsSZTde0ePz+Apcm7jEi97EqOBI5sbNPKhAk0PEl2VFRd9zCnsbSk+cpP
p9wQ/ATutOHkucfmu9WnRfbZI0PwwQS6oOFD+FK9/oNkbCXrFjy/nvJK/sWCML+4
RoQLEvAzRLzEZR5k75FE8IR4MptVSBYeABb6oytNYaipTWey1pONhljyvY9el0CT
bkYGk0BdrDIgSpnkpiROoV/i7J5z0HIlN8jct9J9s757vMZ0k99yrSuwuS5vQqNb
Ec6GM5MI19OYZuGguo+GGpnJRkV/wKhQrNpDib0Rm7614fAoFEyctBC6omzEFCpR
5nWCXtlMdhM5kitrIVLI+yEIyfHkPplwGIkmmsB0xKxzFrgkl8bBri5VAC3Lp3dG
2ynVIdFSx3/+9reioDL6OJN5UEaMId+H5RstuLEVwBY4xrlNrCn3VrLHLy6WK1OP
pHUoRqPGAOgHdCV4ER5S0au5oRKcRei99z8atkofgc9cKLfYO6xB/jWGLyCNKNUU
08FrlCNSw96R+b25s1+k1mz33rN8uiLhhqlcluGEWx6VhyudhsSKGIZGuvl1LEjc
KpDLO1RpsiXqrQqS/VG5t026DL/OCyjLLxNjX9NXVPNicHz8xV0ydpI4Bf+NJDHu
FmIqaaQDSvcz4Jni6h7Bww3VKJ8sx0fvsqkEkOajO0CXuQHNs8zaN39TUxxO+sVn
DHJCUyfC7MRk1wHkms7p+wGtDLP/MDnekEK1zBFoXtDd1ik6VDEj4CGbBwWeO8Pf
2xro4lKSnq1wKVimykuhdU5lxjExny1l/jviqY58rbhKXFFLr4x+XCrUldwXCIdy
aTF9K+CwOmDlV+I5icBobKq2aEkz9tC/PMAUkEe080NUhM6voTz+JAVMlS6lmIMx
REcBS7jBHMiks8XvuKs7rPbpIJ5wQfrDSLloxO42TQsZEI3k7odNn7sFit8fhDEl
Jz+JXvdLnuzQfRJPtxxgBkUXTk48jc7EC07sAKA/g0u2XuthblZTfRKIUW7BgS25
QC5MvpldePlppmWsUjj61ggfsJ5uDlaG92bteN6XYGPRVBbz5VKqdwMN6LZ9zvgB
ufWLHDSn3GoT+YGNOnb4gU8vYM4fDLRa0rDSd8YcpdX0ri8is9uRo3vz84KoTryJ
4WSlh3N0OUFkE3uCGq8b0ugV3yalWcL2kEAA4DJuh8QQGFiHXxIJDBOvBnVXkCMP
+Bpab81JLh5SWD2CMuuoEmHfkAW2s4RRyiBG8uORUGHzDkN53cATvWnNe4zNFxzT
qKsOuWffuWKpfGpxqOZsw7s2rfirIUqkBKZdd8m5ioWORneeKwN1kZKG6bxCHPCI
Y+IYdg1yH2dnEDJROWaiSWlA4I9oZJOo/rZY9AVKTqZW+8M1v4bhNM2NGs3f7Gaj
KapFd4L116KhHtIxTUvbrPCZ2d7GPYE7SDI7hUy3Rg5m71s2JOAXQmYBm6sAx73T
37PINX7Hk5lvWg24vf74lXNjCtftDwwdaiM4inEQv80TeSHJSOo5Pna/afNznsun
VzeR+ITcZTPMsnQWWsapb4HZVE70kbl8CozAOM5FnEyAHF9m1U8JdMJtcj2T0edE
uyh/nsCfUjh6Eg8sCxl/gON09MyU1g8ebEi7fFjRwwmnX/Qbvc5GPpFZKBnfhum8
7BASUcrZzTjR1ZYBphbjbyrrrEuuyqTDu9z+Eoj516lOcjOH4VWG1xnlNmqVyCX2
+NgCJO/PHPv3mCt6zOQNbMtb1KtI/+dGVmz7iFOk2qD+hHfh/ow01vE32mOHtN19
cxTW2k1V348DEPa4R8GozxZBGw23yxh8yIbJh3hMIEyxZRVoUva9snKIRKVK40pm
NwbRuMGHEJ1tjO5U524rwPoFeWXh2NtZowlFfDbeDCyIyVAg9CwqrctByWYF9EXd
4+FoiEUvtx/GcnMVq/UzR0Cd0/gwfA++tSpcXVMbKi4OotidBo0tVLhQ4e23z77P
RfnKIi8NWg38s5Z3kQsD7k9g0Qc69E+TGMEnE6I4MDCC2Ik184xzjWtaQ8kPtmBr
x9scjenUzpoiYybg59jCzrjW1NRSlt6hOBgwNNALMNM9A6TzxUUJtRJV+5KATUvK
Kxh9JwbtIEyxB/cLjv/vedtlDajPFrIj3WorpYkUV/sc77twlY3aMwt1dBct4EF6
sBz1oAggSjI59k6V3O6gIaGzcBL3jTBmSiY9J+hmbxkXdp4ONDLZGdn0VXoNqMEX
5500Y6dOfo7NbuJXlPqZ2+SG0d1c93Hp51idrDdlmRy9UCOfYqBpcs4X1o6JikrA
3hqzmF5WyBLSt1xqIyjmAVFKoJIifAohJId+bKDxiFQ+hsDPHfgSKiGia+vUce2t
stpMLR8PXQne2tg6ssbJXN4AhWnURW0jB2w0Ke9mdLzshMalN4B5zIWKgQG53h+X
NkhpcrAHXpdqJob5sEaH6KPmwJbkdgM/TEIo/wPTX+sJceOqP9+Nes5CNu/AzJ11
vQMM+G0NvG37c4QoURumioY/g27i9flFactJfWb8dbzb4QP1ZO87qvsTI592b7SQ
J7XHTWM8527ywxvcVt0gtmfapodAl51Z8bINargG/8IavGBLVpFFen8DpcahmZw7
NvVpKrMZ7pdO9ncjJQ3AQAu0On4vA01uRlezTwey6l83eZRiYHLEEY8aNzRB13OG
a+bfLGOKxdfarEFyKJyLL8ht0yis2aB4GxI9YxSpHRU6lFeCseJ8QbEFFFs8EYAy
qym3yxnDsvDTOaRtfKlMLsmcChhF+/BqOMtMv0aSUmlsf4SdzotKreNSY0VEsX2D
Nw82+05WtIM81Eift5ncaoome9v6f/qusgJ+j2MuhHSULipsJdZyAqHOMdhXVipD
55RSIvWlGLak5SthjtF7BSVOG55YfjfZs/OxW+iIa84bDNaHm6e9yZb8/7aBc5G0
BkYLcyfxxIuGZaFO/aX9KiERRLpqe9YpGrywwadjnVwFUAJjs+RZJ/xXglJTr+NM
eniI6XEUORKuMkP6tkImEhqBaYP6MTkj1CENbDpHwNtnhgdWDJQzxurCEeROtWs0
8FkvZuoVtmA/mL6TWX3vL3qbqvrGTz/LasMuG1vXzX5ki7GqO3I6/T7gKKFJ+jcc
1I2aDL9m0023V1N2jRssoBt/oAl6rDbP7eSpeV4L4/XDkSXlq97CHAapMpl11xc+
HTTvPQOpDErg/s0R7MY+P2gDFgi30rNjirhqiRRYjDBZpDl9/Xb1fOOJA/f83SuM
TULT/P3I6dbGVhE+qQO0IpvkKbwyA0Nr1Nr9f7Z3HsVz3vq/WYUlSx/9vf5GX0qe
K2oJMWBWIqXE3h71rwWPrWW5Q6v7IEGt37S8lGZG3w4GbUwgmysF/ir3/cV8k+3D
tKPkaQBlR96Qn/EBIUXm8w201cm+9yqStdUo112Okxn0mNUbXLY8SPs/ZApz+Aor
CQxKzhnprDKwihmmjtQWx/cZeXUMG9sKx6zneoZXOu96tYC39mW/BuLORemyRZHC
59L1gwLFdx2cDyaH5gvuZaButXMDYxFJdPEfzHpZsdv+Lpgx/ghXSXpoHlLg32D1
ZbZA2aRSleSU/YqlPvRw1IcPR8dye4mdxVwcby7hkZsXSkYQnmRohOMjHA36u+vd
hh4Gqb4X2A2uqXAhHUcYfHyCceyV59Wn2yGNFl34FCgBzE8WEhYoJrSv7WbH8LhL
Ia1vIjIbZmpu8wClvgr+6HguWoK5VvsiwWDx6S9R6NKkXFN6By9F4BnAQspi3qxm
DpEtSJ3nV7xcbmTPD9Du/R5UPsmf4JfFVCiNwcc0v089U1V60X/E+LNWlD+40OPo
jUelWoJg/D+KMvrQ92cgiruvTBFv5n7y1cSsD1J4NplWa6Kst5xbUOrJxCk91sTc
mZ8AgSVAfkxsLYMgkm3h1x1g3QuqCE3XwOL4HYNtMG/u2S4Gi94JXAU2W2jq7+fR
DfD0JbkEhr9cXXy2blmrdDSKVUjYpeI2PBuO1FvmjP733z/1jUR/l/FYn79toz0e
ZywDWn8JWo7ziYCOppwEq/xuXLwf3RjXjt4e6gGL+CHl6oIWGjzB34rlDSDwgvjj
Q8S3NsfLny7qwfSLLgqHqMjJxdAAMWQpVJMrNmyxCe80hCCizZ9J1D47ZReEnLzF
An2ULPhUgUCPjwXG5bHk9lYEcIgNqotFadWbpKcuK6yxEOWcDtKHoVd2WOSUm1la
XE9+mYi5Oyiq92uW13Tll6xihydMlXvpyyk6R5nqnwJ3OKsnKGLB/Wb6boVgZAig
Aix2Q2RyGAoCNSOyksLTLAVAPOjtP/gWj9SLTZB0qWIbKhcfBan0d+rVBE3QC2P5
Ut1SW7HydqL0dUTrFilhJfIfCYxQuZipI+iK/pEQWtb22IaQ1VR2p91U0xK/OGF3
csZDu6TVKmQyY7Q7sW2LJadQDuTuFEy4zy4Y7co3NugGfap0GQb3Qe3ayvzY4F7T
D8T9NlcpOxaGuk/nrj2Pl3eEe/eR1C53+3Zo/7kYP76l5Haph1St/VHB3lQeTt0k
nU2n6yId610i+HjTCfL76uSdY81d/Oy8nJICLribTVQSML++325MDAf6AnMGu+cp
c1ROwRu1YfxZtTbRXqZIlaDK9oOrg6pT/zKmsR70QX8LOUpTV2yhys9tJIUm64rN
5Uik2uPiZCR5uUWVse7TwfY9eQL5j5aQtWdrDQYDIzcZYhjVF6AXLPAHKRjIXMFj
P8d8DtNvmKcqqISopRa/jLrsmE6Z7jGIYgG5MpiXeRDigCQZpZj+JlqWnbEGQTfA
B1SErrgBG5Hyb0ZN3ZzCx8dK5y/Av5MdEGKFdP/8qYjjXdifSsnGdsHGWwAC/GPe
8/ydudp6eO/mJQA1bCXzvHVPNH8lfGUki/m9T3go274yecd6JUjnvs/sJ6wVZHY6
NMUsYSk1eGOrk2hI7pZTpJXrCS6H6VXzw2qZW3+hPrr25XxWeE9j52iF3VlcOBoX
FtTdVMAiwaohduCnkUB/AbDm2IxMjV0Mj2kKktptrD1CQVAQ4NL2rea6nDDCP5ai
nN2sjfXDpymCo+1qzZviInEZIJ7Imd3Ea5gbdsGKOIgSJxnAmhsZqObgJjFoIPMV
w70pHrP211hAVhcrtqCKcj3bnkmXBA3kMNBlt8J1dzEVPo0R4NKVrcCOob30oq0d
NRzeLZMNtpb1YTxYhN0s04O00B1PNGBq4yIPJTCZYG06bCewlvZhCGqvtgYFo+sy
zm6A4yV9AUWREAnNl5vTw4CYm5m+xUWDID9QbjGniwz+wiImro0O/TgtNwMOeBh6
GQ/kd9a0Lgnt/EWJXCMBgs9y4UnYLQOix0T4f7/993OlGOdtPzzz4dspmkysVO27
QTzLLwTjbxwvPTDCWUgTwjp90QQlfsofrFyJQwczUH7LJjiLpU6eV9xXmCkTj49X
QAm4jvRtZIK60sGhge7d4foY854kZ+KEAhCNHWHb2bXNzh5pBV3DQ9kTxEi1mU1N
xY7D13CmW03oEgaZrFLxiUHtHso5XJmt3td7VGh2v/SAXnXs/ivNlzBQEdrRKMgD
+moV4AdOU7+jc7SORwIql4+LfLe6OFmuicZ/xSqZZUBz89qZqRHAKc2/X6y13Dn4
ZmsUS2aXCIVhMZuTfpzqkXdRpo55kMweLfdwcrB6eP6KbCSC46SyHnr3SnZWZFCF
ng+f4w152cDhlQCB7mc7Ius5OFDA1lRk5GX7pwADdZdw2DrNWl5xAL6JRvpkKLrM
QtYZZ25ehQNltwU971wOB8fbAWsLBl6FMEhVfDa+S9+NF0EbBguXhWc34syDAcxd
mH/Lr2jWqrzOSdDhFHLWSqlpOvHSMkP8Ln0PDDsw/kiPRrVp2ZkVHZTu9V8yYySK
rpy4qdtXH3ogMCXvL1ehXHyyS7XOBaRP/zvYy5PGDiekv5GAR+IePlvf7zkprjgt
AMlpoGcklDQoB1JkLyvyu6fmGttIWyJX9xwJyxkL4sXFZUoEyymHdqxxxuN4bRoX
pBWZJyr7qsWT7D0IqBSlQ8VwKckROkr8z0hBLvzS9OqtmI3uq1YNktj3AdI20tIi
zyo71QbZvf6A4kFow8R+HauE0FXx23UP5zvaIBB2wQ61vKe5YPsJ5SC2pbkLMBOi
NeK0qOGdXdBHjwR7Hi3XzEl/pJLxb+9E6v64e2/0divGVBIoULpxTH5ekv3PX0f8
FkCeViD03E02vGhA1Z8/Jn9t5d9RVigpsfeA4ZC0J77quFHupMjjkXtQHL4ofWOh
4r2knpu2MjhT82diXYs0Gxal4U2HZ+dIuFawby7bKToszoRd1uJZ+g7KVSZco9g7
lF4Z4ub3pDMe8mDsF9az6FTCZih1Z2ptAk+OwWAfSXnFA5oDtz1WkNyhfYFusYl4
cA1bQ09ClDTjAKaqN+uy3JOUNxFZX370HSGq8vGQjt3IcdIDea5vo0RF7t2FDSOU
fVE7rKztwcd4mSOwPlkwWcQmcFOanl6MUWJf2QemAAMrv1dYCL8hniNs2AhsG2ET
DmvLIkLiZwuA0F1WM+k/E84SZ956SWTfp+BGtOeqcueDHx7dEUarnBqY2B5XD0GN
4SCi2Ugm90q47k62OnIW9e44nQ2VkuMqKhpANuoLl2UfbyUb3TjbqYzByTvUkEp+
pndMRwX2iVr2j8JeFqa6mAyDZNQJMi2vLHASc00HMwif5OkhcUuArPEkrfnoE/94
dLn9aJkC4/vgn+9ymruPQI/wZCPpeXondxF/Sqgk6Qb2qWfxluu9H1OisviFqGJ9
/w4B7g9uZHSPiQ82VKl21JKHGHPED9aYida9bFWDBq7GbCQeYFSNzkCmQrKPvl5Z
pZia6bIqyQ/wSOMafqpKLk34sGxO+bqzlBYtAZ7WYLx0JR54f02RRkmzOS6tcc9m
L5HXrX3r7XQQ+lYkbaq9TSmLp+JG2DIh6yybX70nJ02OOrAqDE84mWqbUkLkY5rf
JAIb/MKOgAC4YEPucJkM+lx2zwKju8CUG7engu40uwbh2l0EnDxoWfLWWa8EPDAE
8kqtshIYObfFf0/IaslKgKHRO7JfcqK+ywq2JFcFJdf1uqcDDmSRmarR0xAf0ZPL
t0G4KOSnZXeDgdk7W4ZZpaHBvgeqUgrkgzuhyv2FWBMCvugQeBs73xhfE4rkpXDt
pg0u8yD5U6VErf72OxPF7lyFtg0BXGzpdNidjJzy1pK7LsZGUny9p37WlRA01z1j
zmC+STVHz2+ZaC6JQbwDY2OZGld5y1HjBqwgugpo6d2PV+4fV0yMmgYJqFpt6Qj3
i2wHLCML20GmVi2KN1DWH2QfDgQky0d0MaFxchd8hrebEi/b+RSLSv+jwa4v82Co
+iUFGluBUBZcl4zLaDM25ObZjzDeA4m8nSTa2WK2L4Zod+XY13pzaCmR8Ma0l7RT
1i9BbjXi+g++j9sDzhteqqAe7cQgXI9u5nh2Njgm9SbnGR7YSI4aF19oYrg+BJ3r
3/MLd0UoY20w7aEZ/35mkNrKg9K2hIhtXf19jUZt4HzrtqZ005DaaUEas5cUgAaR
6QL2Q3X+9FYXlTEEpL7V8r0wcgGIXSCv12B1VyEKPWqzJNwqUPdJ/VCKYRYUk25L
kSaU9c5kW1p/CxSyienc0m/B6oyzidH/nsCmpgUFhiI+5/ghd0TKnrrEKqzXXZz6
iXKMR74fZ7+gxzbiwekswEvsDwV/T25Q2xRaqmShXFFgZhLVnE3LmZTxjSEfs7T/
W898soxYEn61eVEq563uJyNGe1tWWjfC3yoKj1/6LVgurJ4hr1yDy5vNdoEMs7pK
b2l8pSpdam8fHxnAAjMYn86q2D0qBe2NmUfVOl8/jYZZXGUKZQgKnE8IT8kGA+zo
GnWSsjrmlWhpeJwJcPypJ56fYX07PC7UY1nClTSv+/ZsDyWQdnzoRx0Wm7sB8QiP
X7GRrEk9jHtNbmq9BKRHdm/hB8aScFXkhXCfqDo8JE6JmB9+ZT0d1reiNUDLjK0k
qQQEW6dOtDpOfzA2pzfeuUDASJic0M8dRJI6x0vH4q9PRxoOQiH4lEoGg4u2kCJ0
iiOL0AIzfWXMW0D7ITqBRnAqR0jmg4fSJ83iqirkqmyWEYlSRlRGPCJG3wf8ixau
0Slb/C7XT5GNCrEZvuC/xGmb3Gz0qpkP3MXVLNYGFadn5Wmmz0Ab/TAY05HL5P/P
K1y5vYkqam5otKWnfv1Y1Cq36hfCe9xjLyGbkypPXIRXLkEKFNEfEyPYmrOaKDFE
t75YDl2RzRrNsceQBNlmOebrV+Ys7DeuNlEx+mkePAgEKjvMogh2JwfPm7dLLx4L
CpDp+4WCpzjHBtWeixLwGyzd840LWijjmGTPfvNEiRkOac5Tt1GrPsusPOPlxQEI
RVnh3Z97C9Anoi9rJR0CEWKM/MErnXseEEuc6fXStOCRZu/49HjpnsusYZYKI7R8
/0ivCA/TKEzbdnt4oSnBtNjOymiI/M58pyauaKsdRdGe605qjUa3Agdd3KJxyt1X
UpferCMysXatehfTSGmx6z72IwqIzuzIAKJJ7uq6OwVaLyYHLnnhF5aCmdk7a1i6
mAbTVrDN1/SiL54KGC5n7iHRJr1vlb3BiWQe6CauaoheeOSWtAfwxTVG56TdIV05
Uw6QojWaeh0lRGIjQzCjDF7BrHEGlGjUD/XU0IZ4jxfbko47pGBBz0FnKNl21iYq
pyiMyoVU7UfVUWXihx3NPps4UUPtBrMBYdbo3opD72lvcud1EXXQippUeZ2MvrCX
VpXYupnAMIc0cj13hCtt8Ue1ztVFLMSf9QmHJ9PhZujKx5XTB42Yn0Tw9KK7MwMj
ECQFWcAGDpO1531uHgyegeAacPvCT7teCtsK2J3j2Al9F3pvcb7k16ITCm2xfgrG
R4EqUb4zNamnEo8Bzh2XiCbjyCQENaLSUt3TF8wQclwCQxt92Ko4CAlx1mSsSlrL
j4ylsQ/xPj9X2scUlaJxNTPC7bFZWNAR88+7YOuy/VraNAa0bgC0HpGTYfxOiorq
bUKpXoTHNDykFsXxFPLRApjEvtyQN2B36q3i86/K5Bxg7d98IudHukcnNZz6Pe4P
JKaK8kSb5LoVOaBteTy2U7YoUXzHgL/cCE9K2mYd/RFql+wrwUeMB+X49SPAu5MO
29pQWPQN5AVsTVXdwa5kAlPWr416ZvtroKy4sXKJtgTNoXlUe672A7GqVraQ6iUw
F+mxPc5Cd162qKYNOp0PnvrEudUgzNHHUNt8OQw7yVnZTaVlm3ZJn2bPAezgJ5bm
5HUbLxGBwlG3cq2ekegw61ZGWeZ55b9k+03Blr5DqIAVpssUh/TrwZFivH6bKOIT
BdvexLGhVMWQ/zd4YwnDS14p6AC3eFJDNt1h5D6QSRukeuU4g/BJiB6Hr1HaokLD
0HgCfZMbgDfvlU4xW6WOt3YTnI0Q87Tj82OgxtHJRNsJs03/ivuxLnVTc+p8VK24
PcG3X50MCErMaFFayuUMjsPwkdJ1k7xbFvhG7WagEyw38KFNfqly23lex966cYUL
K0+f4Rv+EFPCYvHchVJr9XrJ3ypVU9UQ7Srfep1oZJacDJElfwbBXkzHOAGs0EDv
SSk64PS1AMX2zEp9H57QttmHHMWZLfN62RgOMOtohRePYO+o4mgYe5aNCbDBfjhU
brjXIBb+bEJLg/Fp/B7oKzumzKo1pzFbzIEfCWxyQshWFIvRpku1fRiP7F0jPhsb
sa6vE5KcUEHTFlIqo7Hl4/hQzG6WlfTUOh/dZJv+EX3WiH+UDBd9Zn5McbOoOTTQ
hfYY9DaFjao8SyY2CQAWhMQdXh8t1a4iDgy1k+wyuxeh7nqjx3NS/icpolFfgBTZ
KXzoMPJabLGlAATqwF0uEmCar3jklOviQYPuP6tPXwF6doMQtle0mocWqm1LcDYG
34mtlgB02T7hyac3Z3u/BwJ86VAd2MJO8m18y98gXg7ZOwU5JbUzyr+ceyhTBjb4
fA3lRjT4n/NXkMQObM6LRJQvb73/1eSS4hOxy+M2gsYUX2Xc1RGX+rtAyWYzmBgP
Cxd913DLbfE0eywGNEGPmNKSr1ptDjDfTuN1yqD3H20X8iCKHX5VxsyeX8rGkCLS
F6yOmDjJita2pamHyf1BHq9v5egr9sCwEku4fYpKaA6h3NkiHhe5EjEwjkTc140H
aWMmF7UesjdQjQHaMt2tBZgY2Ltj8QDZfZMV/x0jzlOwypCRUO1Lw+VRb/JRPVAv
iQIKXGZcjWGzvR8rlqbSRy8t7FuZxODf+O7QSWWnoOg3//vzy1vIhOf8c+oYWEBz
HIVPrRKVSh4qF56GcPn/hp40Xp/1nm9aBMfki04maxzJ7PrTIVEfTvyyf6ANVmyG
zlhFGaQUaJPzp0vQrQxbSWY3FYhV6IFYDTtv+hP34BGnm8DEg1X/Om21YNMvTN6p
KUF2/GXzfa8bMvdNgc5h9cd+G6WTLmJTAoKTLxj+vcMmQSPYJRiRy57kLm5YXwFA
PhbBovHMpzXVbKkFv4XYx00egyt1/L1wZ4AFwmt9UlB6vcdX9GTTxaespobEdzBm
8wK0TL/EZdt4PcZTtlBuZE2vhbTOxOERfADvMO369YZRRK1wNKK7cZhsVXaMlxvO
aVb1e/+SjKOK4HVrCCqcVl/YVO4IpElLEZHmfPyeAQYk5hgN6fyT+XGKwfvmiGm9
enZwKI7vZhZZXaC2I2mdBSaScVzhwpVJDYZDeT99+S3Csh7T3NZzUJ6223wKV843
JRqeWzAls5au4K5D2kxVEfNH03kYBvpxYfJje765sqg7yDG/QM7GWEXl4aEmVg13
FyLenNBgYM0X226fyhleqZwbG4UZ6DED15t8c1Yz4FwOO7T/c8F5Azy3LBXH2A2B
d2Dt7rGinZLEhRF0w4F2WHEcAHH3JzlsYyqxBNkx3DzZznBhwqkYJgAkVQGdE0kH
QJUOzhpzAKUFRXWR8hP5GH33jg06D5fuXuwxJrwBTWKRGRINhvv5Hf6B9g2pNOIX
+lBqKCEUscZN0PnPbLVgxQyQS/Stf6bffHLauLzOmN49pBWn4ud5Q2fQmwDo8cua
VXghccilV5lcjYbc5dAyU4wPjRD0wbgmlilaLEhRtml9dAvAC9ZZLIcPLfDdMaIl
SQ9w9gwcL9YroDs1Kh7Y1ulnPRCr/ABzc4sbbypyZve8mI0yGEaqWBD1tmzcVdMD
l51kAJNvD16dxHJ2VXSiBxsDGY0rQJ8Dko0RQklfZ3MYGvgHGC1gDTBdUg/GuoIS
Sdi390OrMXPJwb/os4SoNigvtzFwkXzHIvN61gnvmCfri8pF+CgA3/zuMjr5S/Tr
Ocote2+1/CzAN4zQJsgfCzJDL092OSEXsKodzZunBEujLonatQdcZAcRe7dV3K/H
42YQRWHqy5WBiuUSiTKOxyX+J/ARxMgEt7SR8q2tlj9HciEhi+VD69vTlSW+50F9
SDLrSCzqmUZRqeEaoqQEFAxhrdUGZXEtBE1TkPxc0WszLA+umuTiLiXOFvsLbgue
YY8DHvLVR8pJq8Lomq6uH5gd6AnG4Ljk/il9p4AbU/Dox7C/nkJWr6m94HadBtqY
sbdV/rJA34xzyf6wPo3SEP/rztCuYY5ZlEf6zh/MwB3ACQmnYrW3IXpjw2pooDhi
6dbbKtWIAxAjWgYpjA7EnPylemNVF0LysBpcvcSDUSrAEquRU5q6UdkrNpntYq4m
RxDY2vBVtsw+jLjh2Q8uI69fZRurAVI3YMbl/cWjVzhazfKXFuCywyjyiyiDK65n
1Vtu83S/LW3tmLFHvcdeTtrNSKSgjBxBcXoadqBRed5NK+k1Xzz7X6AG70c7GXlN
uW3oVu1Fv7FAtzEALCMxNxB0jNLVCfSW95LQt75mzJWQ90TLHQLP6MR1EbRT6kwz
Ce9zI5H7ucgEBniBaFXuzrWaWfXb6xTqAdZp4jzqYWBdDv4o6ZaOuYAU7QoPLvcB
EIjbWHHNDkwqGqCrbmb9OWXDl5w6VuFsMskYOPbkkW5nRLP4oHGmYIMkEJ7f6Izs
JsVRvYEsR6oMcpxcY6916Sdhku+e0QpUmDlykT/b849ZA2fJrFV7nW26jq5vxBzY
yWyYbbtIBtNNYnpukSIkDtk0GSts7kcMuvhwmuWWvulBKyhpFMXOJ/5S8/cQNwxl
QfRTZYDx8qydQUJcDWbxVcVH1UydVsY7r5qwV9CRYfT4lUYuoZi7kQHeWbI8hCeI
akvjaZCePq5DygB5LkLXANyL9WE8dw3qFRwXPus9a51n7jNrfimGpkDr0jQ6tRxd
JkPAbueHvULulkELp7BFwhqXM3X/5/pRSWW7qWt4HokFhSMAZKwtd0Kx+02a94Tn
YDELx6k4v+mkuw/EY0EhLXTPJxjDIuhaPa5AeVJX9Ra2iaxo3ynJe/gTR+znUn+L
gxOMYXjtzxZLrUNdCFawXK/wBI2URwijRbGzuesaJNYgDyIWaUDjVDRvCJFuqYfG
zSlul3mgSSUrAd5Jsi2KAyfx/b10j92HvoSaMa2+Wnqi9qt6ai9UWBGje3UTEW6S
2Khlc81xdBJh930dYnHbDoJUXRzHGlO+jvy+GrUxDEazvbBmDrggcu42ht9kLhtw
fVqGSQqyC5ZNQUNhUzLjHIC20LGux7wuiz1mV6ZeYpy4m8Dw5eTPoGDQ/x3Fv/SY
7jbVoj7oz1pLxs6yvMWdwMSTxZhqb+ArmPhwuTxhVmHGQxECsR/+LGJuvoI5hY+4
H8nb6NMffuXGGLZZHNQNMlAtC9Nq22AXurIHwLDrAIvTDIpEP48S7lL8to9sGTf8
LQZPt24VeBnfo2tnf/YVP7V58ajJe7ZV6e2TmHq1Wh7B41IL8Iy4eNlTKWdzMTjn
w8nMTX1YDOQuVM44P1G5LYqxVvYZg2AqgUxDwhSfBbA/z/9W8Q3QPf0zy/LZy5Rt
HHaDVCWMzRTz8raUx861+Z9OgmBj0O76GZDNElTXnO5jxnr+1LnOK612dYGnPPeg
C+9zfN+PjAtDQmnZhql8WsH6xSwYltsHJvDLwmj1Ps0VBosCzfoDMXDAZNWpW76S
LhsPOIaPW6ZK0IDsxJI4ByLL+9LxfaZonWZjNgAXkr3kv0tXrMSM2Iugjvh7jvoB
nIV8o92KU+65fwS6nYZAQ8Gwup0rzrbHDP6qXB5VqlkbSbYX4v70XlxBgkcL0Hl2
/Y0KxQZNimrMykFiFCWcRgfwPlM5BNzIOLTYGXG6dPV1oVKfBF1I5g6z79CisGq+
/zxOq5yC8L9CZONC5rWBS9kpukx3xPid56sQqPoFDextnV/9zRqib63XuJiXDBgU
pcn0rPsJzkUqtO16err1U/sfTIjhq/k5Zsj2KQHv/xWWNJonUuiQjLydKKOC5pHJ
74KyRNLNv+wTQniI6Ic6WK1Kux3yASNhnD7bhCiwDUzk36PgnuaqMlQ+uLVQky8P
QB81O9TGlPZ/5cyTnlkbkrbVzJqMLkrAPYfF1MT6Ildv+vygqPk0rWq01sjLiHuy
uAmPCVk87JBlOR3JyVCo/hClcN0gdENytxGCtz5o0RfV2PmZ/+j6TfXsRk3nAZBZ
J1cXK9i/2LhFsxEWsoBF5vsjou2ko67SdG8dzsT/RQ4v4Z3xopjxfozLP9dwThtQ
oEJD09LKvRM1XFRTkDUotHf3q5RVF6lYdSA1nHaSqxfpZHvhKmneis2gFxIiVrqR
v8MsHGrwcqUptbnH6p2br9JJtbmxZURb/WT15thZ/Mch8hVxVxOf+cO9UpBPW64r
007UxvM3ted+5Ui0D3AHeOHvUGXsBBWQVo5+1BuA2mUBMrujmfrTTAcThXULlkkc
bvr2wwXkpEEUxeJP5/t165EXfbNJ8QktDDFkHwa5mL3dgFh/J9M93DNpacmv4jB2
LAk9nrWuAuP1uK+o9gpYcfjyR3rnY8kHmcKWNj0vuZmThSern7n6m57p21gpSAci
F1huP75SJFBuslcmZ2J6vXDOy6KxJ4WQRFXiL9B1fJtBr8JxGktjlf70DYCDWhfU
afDQz+Gf1k514Ps74qHO5nhXD+G93y4Jj0LBzgUU6//nRNhBNww9uTh7br/a2YRs
/oeaV1L6Gr1DbRu+hjQf0rd9dUHQnANQpXxWk5AbGeaPkw4qhcKtLdpqSxIRm+vz
qC4TUJZ4FPZOFuUm5TyoiEaJyl7GuJrbr48tE123fA0qe5ywmsXEbit9PiPThaKX
SSd5hQjHyS16BrxNB5VQkgwg3yXz5q8Zsx1I3Hu/hQl+lind9xrbDGiIjZWHMlFo
7G26+H2AEq05ArLQsJGfLpUH00NBhPOt56oLgpppffGX/0QfQqT1W1nnLplzkXRK
ag5tgWa2jvwQzZAtUGS1ur0pP2YWJndC2gZbMkP3XI9RVOmDl62H5XGWEUwIa5mQ
diGaEEtAwSjNub4mvETaTk+0gD8+FkfP1Z3qg7sn6LpV1sakW27QSuuXy+jF3q1Z
1DIJ7o3z6AHhdxp8KohTyXg5rCCDY+x/Y/kg1l+b62ENBR+nwbFZhKuX/MRs7LJ4
FQ7hEi9Zq6vdRh2+CTU0ZZcCz+l2I8W5qrfUC8tWn1VM+dBJqTYKNMT5YkO8MiQY
yAhtyBXEuuTkKVC/TGxsjsMYwWwS0BrCUUl4OXGn5adoteEqhGGm0Zavsow20PJF
dLsYKpe65qNij+K0yWBJTkX0w5w44oUXar6ZBFLvVSJSoOnfDS3o8xCROywMWj4W
hqJzMYl+BFQWquSyaheEUi9uifiH1+bkwqMlxUmn2KueTRMs/+9MDkAKsaWbNvQS
BQDrQ7e5+H/D5Mgwjy+/q/WH4LuJMRO/5QjtQ+w0/6o5LtSkT+2wBGy8v516DHb1
whXlL1c65AxNUCKgUgmBilade/Qt58BWAPdg6OXE7TIXeuUgoLnJ9AXDdkoORb+L
98g8HwqJD2Pk3zysc5hA8lcksY85PBmlB8HwviBYqNifEcDlYIYo0TamSHrjZATE
v7XuY3rsib192VgOj8NBMcEoRZ41iMv8Mw8Qtn9MnQ60wR4Kz6Q3rliK7xQh82Sc
618Bq6v5uBY+thcDeEYhXT22tmQkYorlAegQN5AptnAHjKFgm1HW4QHCwkQVa/8T
nur1qyf1Mt5uCkIFh10pRlld+cGSHRtdlr6jXaLnWQDgxok7I8K0/o3Fscd5UdF8
9FnvqTU/Al4Bq18v07GvxJAcDR9X0DYw7ctuXek8kIGr9Vp+QDPEjw2u9a9opmH2
XYei5+Roxojq8ouafn55x7uOArzwaotDRkU0gfd5vf3OBzCvHZcYPVIVyaYGE3ZR
xT7zf31S8AW9l/AIK5vEmtUoltz4bmuBR8M5UFNxtE/NSAT/yPgJSns8iykwaFdC
kOWVExGiHvWMYNOpZ7O5rH5UbKUOg4BFRkqX3VuvyE3xam2l83e2GmQAB+RyMMJE
Gra/Yhw0rUc6b/aGSkrKt2deOyLn6Fp3FdefBQ525KOKyeB4nHIZzghE7UCy+/pV
3b17a4AEFFqYJNbsXF2/UVkea6RLn55rkUZ52Okosgt8a1Zeth4xFz0D31QgEJlo
7roZeIGWtRaqjtw1TtF45IcWr0ZYjPKPv+fJyULqafhAo325WCHohxPLSjRb5bqJ
ae1GD4jWzgT4v2Y1/wmUPJ/gdzEqI883GCO3pT2esqqQNP7iF3xQ1O/OIbAWUm5t
4fNsKCtxdyEWPCf3WWdmbcWZog/syDiuzuqq73SmEVHNIXmpKgsmyD8hd0mFw9Yv
GFIAHrusumXuTScY5itUIGLjGPK4r8kIV39l4+/pAO2sak97+fqfSKBowzwKLjCq
6a51qiN69V25ApwjFRSPZD7rbICCNbjlZWjpxP+hxMMQpdbrD/JLWrZg+QpRjiiW
S1iwq+DrVDFLilUVBxhCS+yy0s4cxGgVa6NBxYIT3CTWLJbIckDUUNNJ96gVD+vB
AoJRqsAXk+XWH9bD6r6RPSYwAD32TYK0ha8kxFmOXREsw8wqWZyBS4JN6TBiM30X
x8TyFT93LpT7oaEXAErCyD98WKcE1/k1BZ7HrUPZUhzgkay2hWCOEa175FvCr10I
jTwHVx0TsKqcXtyB7aLH8UF6Nap3bgFA+TgmMb2VhG9qu8DNXi65sSwlXwFmfro1
4nomfS0slPD/1YQGPna/qiLMECH3xIKhcjtQlmfehQVebuF21LNe7h1ZKNqb5CFd
3QECywFbnSUmUNiHI4OiSWXFtXLe2CSGfynMMXmQGzMUQ7P9bUkuBFC5jSRQnDyX
gTwlYJ1Kl375wFcWEY/jNRtMASm1Xf2ZSoiUtgvhoOhdhD9uCcsvdhonVyWmtO86
ipUL9PyOr5p3iyeCAoVt1pLUrRuUfV5EIwnaKty6spJWtHToA/lcfeq8r7LS0vhG
ZYshGKMNM/5U5S+ANgzky1oABmZ+341/RZxCRnQW4mSWgNpKSCF9z9Sv/CCQfsiz
xb0GjhslV4d+FMIbamgwluKGTyZDDwFMIwnDSvq/Twh1hpssNozSqz2WY5Y76Wn3
rvWUyiS2oDbGH1B6wMN20Tsgzg6ft14dKp1a5/SURs00Ow9O1/j+R/KiIZOTKX5X
h3liCDIcqZn/Jb88QI30lX07YGFH2PZEy2TwSHcgIDqhMiJopCxqPbEO7wiOv9YN
j/7g/efdD9gai2h4zIFwyG09yJO4zTs3hoQx8opEvaBQNuXOgeMMMnEAECMCtda6
Xge+DhGTQIFdMHhDS1V6pdEEO65OpBtQ9xrRWn+jwfogj681j5Sh14WAyhNrwVD5
a/9xQlTldkUqYqfRKlc2HP/pRaoPJSg3ONyk8lDgVVUl0PG8pXuVl7/d6cC22qXt
auGag2brbZWThGampilvZGFuU8w5RVHTjx3o4QEvwAkrBcTp2Nmj9pTOP0Zu6z8m
s5fTNpHc7HF8jv3bm0BGbbbkhVy8EZgh2pxJNSw62euVlu2uTQe4wdsuJ98ygB51
cU8oOflUTFWVR5LTpnB1w2O03TJrL2fAW6znhUvvPLge0QbgvWPkwEZw/26Uxp64
+TbkZRACvuqAos89rSPughhJrf5KpPbjA02orIe5YGf+PXbLYPuKrDu1K944/mBl
atzKn6mtzrasLwodhESrowTwhkfjePqcrBkiQQ7n+JFGKlWJdmmk1XwFi+5bOWGJ
IzeiYlxPeyj0ZXY7h3E7lQ6o8dg8M2uxKS1fwJ41u2dfonkOVv6lBGzSoPV5gWhQ
lYF4s4QHiDEaiCQtG1zMb8otS+hZ2UxQUnVeBMM65+IC5RXWn3kpgtABBjeTL1/p
42YL5pCcpnMX3GxEtVFyw6cCM0D60THgvsbprFr1m1oo68M2V092c8CcJCgw/oGg
wbhtsP8rIDvdD8EaAgBwWVL1dB1oOqR2a2RPmp2uduySh3o9ccGFBt7FSlvkh6sk
P1v4EuUMMQ2OTMyi+7KMzHeSXSCbpiUu+5LcY68MAlMBYX1MIJ3TpXJ5dfOIXndR
Okvn0H7bEf+m2DeKK+iwiuWo3Tg1FNLnYiLFwwOchvJ2xubHSRN2YFo6uDi2qILS
KwO4XcOz9ghVDdTnVonOkORYwvxMHQQZhJdSWvIlZIPQfIJGgA0AqyoL7KIv5ADD
x9krumkl5QkFOw3u5feMiDKCpM0017X/AWojb1+WqUxvdCOWzBpFG4BF5yYJZBLf
YQBUvne3NTkzv8zgriPocVVPNwkGFCdMoQtUQUTEKo62bIaCqs380o4L5twCIfag
wq+I4SJq0mKxILpVasfs41KGaXW749H0qGnGdgieg9O8D1qYgs0vQ8Py4fnCzprT
mAGoc6M4rZG9V53TXjbmbNtSnRDgxYrbD7nTPB5jv/ba8ouQ3rWmJZND9sQrzcQi
/VKWHuDeDK2SsucBh8HYuBnRnj9BTgXrVAAMclJt5yY37x9adiG/ahM8PsnO2J8P
oZNZAURTWPelLDPvH22hkTGf6p38t7hJjzDR/PN/PNfJwiOewCGFhW5MGVKkvomZ
OIBmB+zmw+/BcPu3+VvumzmjU0yvIql2e3edJDI99TpGHA49jhMOIbUzH/NuFsx9
5ks+BC9aCay+otIOEJM7JeIRYD5QQ4GGMIu1+wU2pTyITa/E/Ts6/HvMYcc/PB3i
F2qdroKCyyDNV+5/U/RasqOfKYefUWRJS0lm/dZCwAPA4QNLBymeokFKJnHtuJCh
fdRQ44a0bnaoqlBR3azNlw7P2aXpEWdcpWx7GiXJtNAxOsJ12Qw97M3O721TEacG
Wh7vtb/dPOtp7yGSzjblWd/Ka/OmlUTSNBppnBf9mjOsMJ2mZ7F8Gj7ib1hqYcu5
Mq/XeTdazJwksNx7DDlQy1cTXyiYWb8py1Th/P0Nm+QONDFhOHEUMXBhZa7SLYIG
8G+GGKkRSTkzAA0l8vcc/eOAiaNzXER/cuOoYheyFaTjRxsXG/eVUCK5bTzzQTT3
GwXxr5wBwDLK05Rnj9pGQVroB2SViQrbOk/t8I0/9b9oFgJEYP1hdqaip9O8GeX+
+s5QJI9DV3woZC9vaAnKpYIaU/XcbacULOYWDxbozkvuCdn3CWsmIWrkW6fk26xD
41aeKbsNPv3a1mccUfyyaxSrSvBtygT9aBpRjFH97D+mh+Tjc5pe8YPgxlj5jzf/
Le34fQSIfx7Wn1nq0DNpxgiY0Xoo9rfU35XR+Jvsb1miyyt6yLDx4at5gZXHMa4t
GEV9p40nKJbizYJQUIs7SVkiZl9xKalcJNyCfJyE+IiIjf5Kf5sU1T7HFmLCwA7f
tz7vUgGhBlEBKC/n/c9N1qWBtB3tGg01UIzApaNRRj6tSus6lySQuneN/mdbSh3w
Zh4ivYUeoKXiJ1HVUfX+tDfTq5nuOnwFd5DK2V8kyuCY2UEYsmo0KoFkMJcDjuhR
d0R0gRssNeU+oR/UL4pZfFiFc43hf2oQHmysvUNXKHAGECg3IQ3naG/SLOpSL0RE
ymkN2zlYC/3I3J8SEcqHAdFD/AfKhWVEs0zGTJuaTsucbcOTyg7r0sJAaeY5eF7I
BAajWlzh6tB76T6aMdxfe8l5fFdhSDh+mADAkpOMhsCvKI7NncCCcEsl+6er0ONi
gXtardcXMif02pT5ppcY+PITwFLkJdb0vd0TYyVzjtP/xdHLBmVpVr+Sq3SWUGBG
se6qYewHKI6z5Cp0/Dr6FYmy7w9jmT/GzZ5Uw+j2heJ8kKUjZVi8eoooVFT1B4hu
6D5vQWyRk+62gmKeyD1QhpMGAzcnbXTZWDC8vzxhsnk56h4NNJa9rIvynQztZzWv
+jQhsyjfe7bcChFu1s3s/RBgA3R1j0KGORvnIc8tusx7ADmF1bWLXgDtdG079//t
hOOwUKK4alf1Olxj0axnjqDibrPG8If4avkLkInexrQrW6W0QSGfbFUQhAkf7P2F
A2U1FVzUM14s7OwCezTuIVPU/6ekI1EodUis9fkbvkt9cxIcwiQF0dtMtEgzK+qA
2QMsTWyZb6HHy3CGe5f3+3mRS4ub/bl9uq2DqAHV43GMQblTwBLX/YZw2uzyt2TC
FpVIR6A04LOutcTOtMGABBYmoOQItgF4dGbLFi9619J13G02DZ0MRIqKcaEet/cn
HEDWLi0+4PFB3cniDu9nk0PLJ3EnPqv5mTb9YLVusvNOz0Eo7e6LRm6J5l19+0Dy
m/mNQ9cG97wpYGHNUMdXGLBCiZB4c0XbGaYe2RVHWdutyhQ1ruqK9M7eYKxOwX9S
jjbz3mczQLgWb6hhmefmqXhq1IerzVu6IxJ6x0vOl2h9kNsvRXfCV5FCvbfwElQh
Ox6NygIBvmyRSYF1aIKOQ6W6ZJEpwLKZb8Z3uKXA24qbnDi1klZxDWw57iCQ9nGO
8R4vCdRuPQsjH7SC6SzCeKb/0+z3ZjswA5hQ45LRKRYxQBtd5uwX/TtFEH8QbMPn
Mm0JduMBIdq0K/ntVemUlqHuWeEtRNizUkcQo1iDNa8aOzR2VTlQLfz3pAyV1KUU
hTs3LIBekot2gONDICjDiMXLCbjC0DT5lC//gjYUImL9MnW0c4ijODLzf7Em8cej
xroew7XQzcJfa+ROH4WDtzW/dG6SzQWBvce1zMyQaaApUCJxJDQnqmLxCUIBJ5Ky
MWflzuLWi1AdgB/O+gzUnl3MF7s4j0kkw7qV44gpmz535nk6XhJwo7zY9t7Z58VG
6OQNnyuZUjiTm8EYQimYkVx2sKsTk3P0OFrQuDpD8eAB1l063kErcalj+kOOLOpX
kOlgydEJTBGt9faOK78PoDsX1sov8Xu2bhysuerf+Y/n+tscJpwyEZuBMQ+s0JiY
RRqcxHNJnCqiLn3xTNXHha33d9gc9DwQC6BeF0W6bDZtXmfR1WgLLEbCuP61MHsI
dFWJh5q5SYmhVScgFoC7cI5zPmyjGTd2ufccSvkyBLCFc7XrHaJ7eDeGc9pvb0ET
qLRvDjb9EbrzqC/uqDHra9W8s5mhQN9E1jCGhzuAuyvzYaepP3bM5hWQZNDSWLPK
sTGAvukKo2564kDkE3jr1lcGRHIfWDX/LBHLsP5xS3gK7WMb7RqT5HmrRgDGk/6K
SB+cYGerKU5siqajkFnVOvoZmh6wsSTc60TRu+Gj0lo/p9Avso9m0UuZ4MI+NKoc
h6wqgGbdKz/PA8ZhIkVKVIhGIEKu78kqSbXYZEBkEISFQ6VsOEoeL7u8TB2yRoT/
XO0ihCkGyAF7atCPRuLuV59Dq87GPGEzy2XJlxcAZTaqmADgDErZd/9MgrkM+eHq
Hzizg69YV/9n+PXpL7eHl/y0dD12nxy1MZqXQ1G6y/gNnWbfpMF8IAnq56+9swic
FV1vMJ4LIvPmD20h0inJl8hmnePROk/u84GNp7MNyUxEamiBdINEsTKGyXv/7s0h
Yey31BVlGU2HrTXVqwZLNL36YOM2T1kY9SWq161GYdSErIJKk6U+VBg3mmvnhlF/
tOzUkWMkEhtFsv5gD2s4BfNhZPFs6Mg0Wdd11Hx9Gwpq1YAAYFxCjy6pPIVAvFj+
p42qp3QIwHjz2JrST/2CwaiFWjAqA4LCJJo+sbG00qt9sZSlXC/uXwGpib6TgUWo
ShdUYt7qdIMso7T4M76AiFS0JEsjMQHgbWakM+uT1cdOmRvRlj2OrjCoFlRH7qQl
bunUpnVSOD0raCq9z44BRMILzYkhDt+a106KwtFkkWxYlmuVlq6iQAQpaWkWNe96
Rcu0i0/THsSzIG6fAeoTprFBe9YYebc/J0Yxv/uzab3mwezVse3gvazaCfqrqNy/
sunoNYGpTy8rWTnAQiXwjNItkIM4XQq3UuCetjQfKeyCGfHjnxaBlDTa0ZvpAox0
8Pwk0NIXtqaQOjeLCIze8ph+FDKdHNXctuCHgp/6zXSUmbnXAG0SKCFoRABDXPft
ahXzO/9sLSba6AANOTTqnoxmSL3HHdU8PqW2JuxOC0gqmBlHFDi/gdlTKWcuQCcJ
RRm9wMW+r5zfvVIhTcZcLqc95CgoN7Q0KsqmLkjqifHXPT4+xJ4jn9qnPnTXp44j
/wQHidWqRm5XG9bCjU2POL2tYIjlwkepOfIWN0K1FAxGhHe24tynRzbVPyAuFrB3
AYqdYQmH3s2ZSYVnJu0IAetsNg/jcVl8v32aopU/O0wLnDWHZaponeXgvAwkql79
dJKOnITqyrHE1vR4G/DpzuPsjhc0br2JDfYq6T43K4K/lSfUSoZXPtR/vq00CLUx
BmDVEgSQNM94mLb9HOazDHXpEv7NP1e22z0jr0mpPl0Js1jeAN6OgCnXH7PIbQ/3
VuXBoFeNgvtIKlXSsFHVXb9bQ+s9B3bbQoMT/SrWLa+twQhtYsN3VqMUN+FFO/kk
66m+egTkr9jIFNTC0F8FxSKhhxVanV/r5XnD7CNvWmtl5bg60uIrn2w6eaLF+dG8
eMM84udNK82lSPxkLAcUTCWTpbTK2siqE25rk9Xz9O22CwYyleYRhWjs7cmg+ePH
RPtuLoOwboqzNNmo4hbA+d5VBdoHnqQaDEJNp5OQccbVGpKYOc1R21iRhVb9SZzU
2W9V6kYPZXp2VY7VzfDm0y+Elf2c/+7FhVOMVbKYuTo1Ezf4AXGk8UQ+R15rTApl
UgB6OEASu+A61UTDqeiBDDlpblq57PEqujX5JpFDwljxG9DjhEg5mbKvLe1xN77u
lbcK0aqZqazdxDDAnt7b01SYg1pctp71ez7/xMMc/BUViRux9Lc2KoVk6e4WmJIK
dnFeMbw5eVSGQ3vBe/n9o9Srw2IAAbaUYtxLuoe1YBuPa8nfGRpai479P6mkO2yf
HvjGfXRKOr6USsZBgY7hE1/FesU97kTPhA8yr2VQoUY4pIAanOThzjIYgFcQbaZw
FyhYTPT16EmyoOFKYPWQeS/ZpTS9ItgS9wrsW94wMMRsU/ynL0tJtnzeMJvRPmIv
bMxroBwEKUCXkFgHDy8bsMb86T8KJIOhfvIG3kbJjGz7IK/umgZtPAquo5qEkJhw
odrx6Mq1kxZgWhSi4arWwpoCh62cqrmzZWc2fyDgQbBgU0SXrO07NcEG3c0L/UbZ
oKQQaUclwNifMe40O7kOvo7BlRDLxgHHQ7gslialJyLTGXw7shKdUPkP+xap+a5c
8fTK7mCd8YK8XQ9/DdNakkWJ6MZsoDvQ2rR8xRsUF49OEGiioZBcE8Y31zNDVHPu
90zC+K17seENJWwb7049UbHEdXK+bod/vpnnvhpA5rHUnUgabaN5eM6G8yt+Esy/
qKCwzUTN1bJPKqlDfTsqbUG/9Y7JzEn4+bUpEkjypRlwzMeap88rFArjaTGE/+Uj
EUZKxXVjxd1kDtCijyYSPVtrPG85e1PQGNnUB+7Ees7AhhAsvlyWRoEj0Sv60hR7
MiVREe+zv9JXzy9cqPocsYrGNqu9Qln6xB3aTowNYb9gnwepfqci5N/qLtvL1+MK
NRzZOnTg+rvuTydtgLPnk4ykTKPpPPACXoh2V3e2Tc0Ut8NpG0XmlE2+NfjTIqLK
mrB1DtkTM+1eI8SVcIHt0XvUcpSkBfI+5hqyiwBofJbeXOmxa4oaCEP4ScbybE/T
ZQtuC9EvpiwM3W8HbKqOdIvvX18n8p/ccHQjLxFGEPhbkJ3wBTyGofFHyEsRpt2K
hEox0Jg/nco/3CikCSPZ0sEG2NQaDkYELIf5EckAvxlAVc5T1HlfQCKtsRySitWX
TGWaZB8O4dvRsPpRxLaGK5p5L5443RlbhL9F/S3KyjVjc1hEuqx5L8PcrZ3gkRU4
Y9pQE8UNmvFjBo/6yXgb5CP7RjwGNH3JwEi1+AEfKfbHZw0ZFJLpd/FFL5jjWZyF
64sUTNfj+1Xp5oSQF2NZBCQavEGhW4PeNTS4U0jzQUZgwWIsEX+Vpszi5toBzH+7
hXPcfqyuA935nEqCXkzJ/vXMvfMwSTHqbW1iPyG+w1D8XlvPpWeN0aCRuq/LDR/4
zfzRQqc6Ag5ToRu1eBUONSJ43i0yKsTQxhn22gV2+O6A2SQ7tauJd+ydxudoSpSz
M45ViPOyOY77WckLq1gxXHGBrXDBmdulK76ADSMJAVFCTrWhZpEWG5JLQ+GoAFxP
i/dRrQDQks0J1ZDYZQwLkz682MB0siMXwiOu/6nG4Fc/9Omg+QOg/7QBcKG3mxYC
dI6wd9DZ6JCb90eYlYenWWF1+Y275jVGscAnJOmNgYjxWYytf1C6fozdehBjgHb5
4CzrvzEzUOAnvsrdYltU67MXmcbBqqxU7FT+uu2hU6BxAdi02xqmVXWGjFFwX6//
7Uqk6+04eVP4/n8s0Oew3N2f5vEojmNa9nmWYOGRcX2i3RmjPRSbq2ujX7MSAwDj
5nEhrCERi/VKOJuQs2d1vsLoDXMJRcywI49hlXSo7SnOTobUbeQ0c6FZaR0HzBYb
iH5iJtYMjyTGcNf/j/QHMqWUdzLfiBmO9bq5WD0l63GYtDr9IPi2UUYZ+bPQC0jM
qVhhcjyI8tg2ea/QpZOXAGWgEleKFnr1ilBHYhjlPpbKIOeRfbmViCbxOWdikce0
gWjdBmVIezir6KP1FofCWbSfgCNe/o/ABNeMxSyF4PJmMVj/lMiGUpOZa6NW/vph
1chrm1uG7q9hdoKGEbqaqvPSVB/uTP1pgJDf5kj5FHvX15bhs72JNSvdfjdZvxr0
545Qfj8UNHiK4c4lSch6jYkHmo4HxeSTZe4Ub1wBFdPLdB1fTFQmUCcQdJ7FOIae
J1syGytvJyZXJG2ECZxyUBF5Eq35WknzfU4Xc30uP9z87mBT/c5+yj9PTifrwTKl
Yh/6swbp2EcEjZSee/btMudC0YdXBaODbQ23v5vIQqpcsqogu4JUzPfzFkzLNjtV
YWTg9xgF96s6ntfPBptY+7uOShROmTu6EUPdUNIu2QWkC5OArwhp0eTJ6yjiat+l
2NJNauK/fAZVm+MySMn9BW00Jlr9mzg3RmuRAGgUamczsUJG+Uedlfm7wBnF5skZ
WV5a1cA+n+Y8V9vI96Xy+6zXG9bGLFjav2gqgQm56xDN+bULD7mh1nmu9cFOIN5Y
hS+v7odKIhqjEJUs7zXdAeQ1JZNgs4CP71bWN9+8n9mtnXFzs4xDuc6DHDB+lhMl
7OxVkd1wDZsCvQNb/ZMhOROQxy7SqQgl6nIu/oxN+ZsHwqPweVhbWWGp+sMf9HPf
SLLiHTOEu+YT8Asy6y2gIpwU+urFpMAdLqteEpIqYjsGmm6abhQAO85qD7Wfb6e3
71oF+G/ZqXrv7mPKN/tGF9UqsHGtr0Vx5A7J1yOWZhSDerWkB08oLfkA2Rdwiz/F
BIoLaDFBe78sr5I+MjPvHdJaaidHaHrSs/FMJkD/sMC94S3R/89AeIO8xAHeFYQo
b20clGT1bl/TrFyaybGrQNu29X+6anOeRM3pU1zLEEi9tBhvnoO4NZ5OLNoEtB6H
GtC0m/fSTc8kdxvSnZZEPf0nyVQRjGiplLl41wL6CWv6ao1uRH+pBjr0XQEB8E3C
bfcejt1zm61VbZ0X0NinU/uiHLPHvbaJK9qUvdFXtDtcdh5wWkd8a6yIreBEkFlY
/YpvZZzNpVzKqMypi0vqV4KPRs0NAmKJM1FE2eb/h8QZEmjczGFjEe18gYd9ByCT
A/D9O0JW87gc1NYwNgdQyrqKUm6aDCrvpC9pXT+CfHdh/BQLLv6IbzX2lVt6heCA
Clx85cMYaU9x5H8om7JpnILysM4QD+aKs0kfIlJb7NE5qNipKqPx/cU07L9YCcbN
YSnAPaCl+q/FoDktYTawQxI/lALBR0X7ExEevFQf+MJcVWq1zj70/l0HolS24lMQ
oc+kXpyGSIarWWsEqKn/ORUB9jiQerhqYvFM/vXTPyLisiOspDF5lB3nIFuCU6vT
jShy8sTJdzCmcV3KvgoDEW/lYrA/MBeVq2qi8mjbiMvRlj7kytWzXy7xma9X52ff
+2Yxe24vFt7jTBofOyAfsH7TCj3R8ewb5tI2SSAdqfiTuex6r/5nb4gnaKId/HUy
KQPnGUs/Lo4XJ/oyKXvKrAx8PMeoIRCnJB6d5ZT03a0SIlpu41zhG7cV08Ci22lU
yqUffoejXCuBtpCIcLZh87uGAiiMpVAVwlH+eHhakUU2bcMctpAFjO1O42Kk1WaU
wGF6y8GguYqAH2ybWP8VfdM5KFuRJwqudQzcGFRopXje1hVzAxJH00BdcPy7P9rJ
gCR1fNVff3BLCaAaspgIJ3CIMFTLY8k9oabdJPoSUFIPcr1kau1qiuUn6UWw+rBx
z4xWUOGydZJNJSLSwsy16VbVNdZKETZX64aWlSD8EyJGJ5cWnE6ceJ4VAsXxoafh
h76NpZRFjJ7nrniF/Ed6Vs0vUFOGDEVoBL2R4ATf+9FjAqDjWryzZRJDNYaaYUgF
SHi8OlkYZV1AoYZH1KFAtdE/E34O+bRAY9iMHGjso7l7Wl9ykdVEbxSK1v3UNQQN
wrvVcSpZYJi0KBrU6xOBeCKeURyNUUtPpU5niO21uyrjc7OnLrwqIYeAHUUiBJyq
eDBLa9Ob/y8XXULL/gsMLew6mWDt1Pz13BCUeeSDVvWjdyR2tilZv7At0cnquL+W
xhi1xo37HytanRV7gy7CSnS3AW+RASLftaSgyWP/6Xjs+NStghytaxg48+tRQ3Y3
SBgpk/Y7mhxt90parpE+Rf3kzD1rjgM4JDdXTC8rkAqUvI5DunQ7/e/PowLTNF0T
EWSRbzQB1F/6e+QSHmIzURm20ZDnVgquONkCfGGYFMrmR9FAEhNUrtqajON/xxJe
l2K4Ct6tR5GdVNZeQ/Q1M3A8v1c/WTfDT77BFo1JC8UCmRwH02YJ/K5FNON91Aok
d2IntS7eIhuPWjU+twqFQ5kTgoS8d0ZwxqkV2fhHtl7s4AGlW7x7mc0gI8OUbx/b
tre5Yi/hFbToZbgaUaidWG/JdCXerdi9CHN470+LquW+WtCTnqKIfWL4QQnoxtWi
+3C+Y9+xmg1V5ht1sR3K+7cR0na831my5CEA36RMO/BZLRUALxtnRLIPGrlTLaVx
+KBhEIu111SPLyZnmi0PuiJfgXbHdfSVmLWOABBCZZ1FF1H6ja89hsuh5nOSd2p3
mg02rIQQA6e+omSrhTUfoRIkQkHMYbCGXpO0+cLcxw+l35GjmL7gRpFGnHap6cfg
eWmoy+WHH0l3Lqnr8idtvfIzO8MTo1N8Pe0F8Go34I8JoFEYeBl6n7UlJTkxE7hH
THvfdMND9PSmyriCpxQhA+g2baAhCGYO1l7yuKOZt5eQt3ZZVAVyBFBEG/D8TjoF
XFO/3cN6LozmYANkdgAzJmu9d/vIFiSN9qS96r80OBqPvy5FY8N5GKSptHDK7/ot
VYD8K51Iq4VYs30YmIgrSWOJy1+/UBUT/z/ddBKB7FUw+umIrCHQnFLv4/rIQzov
X+JUNfOtJ+JXAyHKo8taddQcnCQbbyjUtLRyXTEM9fd1faknS4XB94OFMFXn7C8/
RPHWUliVnIR8s5ML9kY04QlRzoBK0ttQH6fDMRGiDAZO4z1u9cUAOzvpgdYI/MTs
2onlAPGs+A14ZRtO2Q0qCu1NsKTZy7ED8z7K0atDPGMEy8htAJm3aem+gHUQ/Yk/
bt0Vrs1eq3Q4PA9mc6zgk7SMt8o3S0CaYBeHh5QOmT1oS6EjT4lnZ5BvcuJUe55G
PRSDnazhImUIVKiid4hvd1NVuu5PqSO1u/a4hm8AR4XuAVdgnJFURL7J+jhtT3/x
REi3rWvAugSoHuDP6+MUeWhRSvAEJFiMNVu96tNB/e86Ij5G+Ep3y2JCPe/HaUtF
Sguh7+7Jz4G5VR+ovyj7rxyEvpTRigGXYjJcwLJGwXnVOIpwJzey2c/VF3N6b4JE
hMx/+PkG8uKlcZLBDGYo9XddnBGVboMK9YxCmLOUR3UgtCwCKBTRa7lQRTldlGci
W4EsAMBkWfE/YesgECN/4TZLs4ivnTzwC3a4KPFeFu5c7GE/aFSevPV5njgYzsIp
usVkEo9tpOjdlBL2MeoRseZeothAyfvEujf2TFABDqsNY2oxQk2yKeUfFYiLyCc6
Kh62n4JcDqcv60h7GvMy2US4LQj4jKOVUvaS33zryRkZ4dp1DQGIXp1S5hQNNo0b
U3KaRWXma5a3x/1kuteVbinBEfZJ3NTnhsq8CkgXuYK8LDRY39D+N7enWr70PT+S
eYc7TT0jayz+3CMnc6Rg90ipIVX2BSpuIxk+5lbIgvYhVbxChF7gmtY4RjkQVG2N
T1G8Nh37FWPHY2aPzd3LzYg21mIkvRYUqF4ysqc9qnFx1nenBugD74TRGrUwAiwi
p5vnfZOEYu2vE7vCy9b76K0kAF38pp1WvHn6lQjT1ZtsNz5NyQN+pvIUFC0NgE3H
CoE/YpQ72Z90JnzxFV+gybWjJqlQXTTvNlp/qaTY+8MiMyAKs0/3k6X1O//FTKA9
mO16YLu8yxTAS9M9bHvxn3uBsJiUEMtQGnNisWCG7I0/d7HzQi4TkS3z9Xrfluws
rzBmchgDSVVXd199DJBgkmWvGJPUqMZSzP+oRVPQARNpbvedeJRCHV2/V4nvk7vZ
ovHTUjnoM3tfN0ux0/V2l8YXV+M2P6Wfh5o8gxEA3ZRAqknRm6X0ynHu97IuPTR9
coU78jGhIQlRvlUcNWj0pJRxNrVYzvYU6lXko2hIQf273ddE/y/0BR4LGj/kCEhy
9ti9sVw5guFwGMGPRKm339PIPRq2SuJpsB1+PiG1BZblSSW91PWf5liKxdXcWMEv
NEmV+J44tRE8kiMKVnTrm2oxzyWo9G4p2ZKlhEuV31t84sla4e5a/BfKv7Jf9mhT
ZbbPi9UHB/IwlOrZ6eHtvtb5SILwBb90P6xSuph1ZljptOiRTaoxXBBvVUIqmWeo
8G3Bxf5SbPWmVEc4284+1LSjuVrT3CuXxdBxwdmp99QXC1YSMWRvYU8rUXUlt/Ma
zPmUU0SUsUGBVolWJy7DR+JlNlN8dLG+54Nma4NTt1xnFCuxoblcw5s4PB3z0sJm
WuMMcZ4v4WUWu6pYIn3g4H7YEW88xoCbk1Hha/qy3wf2v1dWclliZjoBLTCWBCae
IDADM0Ksxa5NCjejsYJ8eFuNX7GTRhrx/Y7+PKPwDXNF6bqQ0wRnFiwQ0Oi5Jn70
mBBxN6VqWVn22915gqBFL0Cr3UxB7fOM7GomNvlOeJ91VJiz8kc+CeiL9I7p0A3L
hIgpa6bazUm64daa9EvplDQwsZaWKSNjjblLBp2sNhHhVJcq11ndXYIyURtIwm/4
wXpU67AgW8R+HpJPjelcnPtfsE5hTNfBd9KErEzwb72erYUtOcgF+cZuG4PRM5jp
IFr+tD1jwZpLzVOofnw++nANGrbVBGo1Am+qwxBBgDm3rvhXu5SrcbxsWu9S+NG2
g8z7t5ulRRDDEH8l2qs22t1ePBRUKX4ws6fcb3/YyckYCtERtaXQPk0HVjxLBq0u
tVr3ZtPZKGZJAKQMEP/Yv6GnnWLVMC0wwiRL0rAImQ+wgfyZBy4fURQefeAHsJaW
jG3bc9ffuoKLhZrKmUgKAge1MRP4x6cBgE2l9dsrmFQ6OwFQDhls/wiDsKlQFavm
RtFOEqGcC6jdGkeq9SE03JtTjTcKFLVuAyaMkwxvXtIgCpH5OyW4rRkmqgYlxg0i
KJBzDofI8TKSKJQQIsNH5U0tR9vL9L7M2F5dzLsMa3K2nkjD9/I2bFxyee5dP0Ep
QnyN9Mz0llCPLZA4/rZ1RZXg7dpXssvJQolIKCbnu82kXiiqNCgum3SQgHIYClSY
2btuqhB/Wy/L5F0nuHt+xNy2xX6lFVH/vlBZ2M6u/gi4MYuAIUFzYSryoKiIo2ZU
57WrRMldQ7aU+cjGzT4s9zgaym9Ac+r+4ixz+sWsQ0yltZ/atyRv45tc5uU+8Uhq
LajELUJhysEsk9VOEQZZ+HQ8mINzVQJOT7SjJIv3gtNjxBg/5Juh9K5+/Lz8BNj+
BofuaSP6QpiLU53o6W29qFuIYCxV4VqPNB0KvQuPDR0pdSaDmOZTqpG9IDxCmpTO
ctFKQWiPkJ8JOsZ7CqVF9RnaMlEcV1dC/FU8+DxZUyz+UiwqY6ZfF8fXrBJgToQ8
2L4YNO6YidSgCY9Sw0tsUMzq5ib09KmXCfkBzzDJcTWo7URa0SJzK4RyXdQLvvEd
tACzY4C8LYBJzT/fzxUxQ7avdvUbVLHHBpwjlpVMkzl6vv2h0flwe1o9bDc6dqlD
BGGmZpejCw2aMa7FM/PrKomWiK4dN7Nzf6JIYUYK1hL5U63vvUGeQo7Ln5KKLwqY
aTlobnCcejdwnT6Ty88sKmRdXzMTOzgdxrBfWLRoEs5dKIGa/HCuJBMHNcJjMtGl
G5EjmtBv4ABhshf+Q++lHXEi1Hy85MYV6eHGKwLFpyWdWsF+hzWbCyoicV5eGMhR
O0ymNxX0jRIHzKYrjx1rxnpDnxtFFCZ5a6oZvTLYyHtp/HsauVy4scSbZl+aZDw1
kCP5Cb6vIyoUDeNsAxU4U4hDwvOIZf47VPFSVivgluhUnbWud2BW0EoRKQwTY68M
A9BYKuwdAsE/aEJ7Vl47vfWchVEchvslHRexVVGn8Ev3e8a127nEc1i7nVUV6AM+
JhmDzpvM8oWuHduAXHPbJDWR2anQhGcgrUARj1saUD5Rgi99C9zzyU8PInn0gzel
6JAZIVQBqwGZYogNdvnJmNfFZ4WLbgYksDhVBTnFTrlGQ6VrEXZP4TSgxh0slACa
CSUG4d2c1PZs0JspEvxdfyRcCZpJ1Yu6MLH/NBekGirzWDWpnBeSep8gjveyI/Bi
Ken/9z7jfOA90qqI5eXJvoUeEnDxvJqC7bVeB5UHvt+b2tM4bs5e+ZaVxQeorpzn
yno2Bec5PrrxSyDXNlrC0tuDy09vytm2mVQCJtmDa+FOID5r+10F9QfJ6qoOpLzE
1EorcoqWHQMWI1MqZKUN0+Z6g/IDxvG/raPGDidwKK6mKaDK8aEvm6up8qbAzK1m
B+gbFeILViCc8TCHjC/4VPP+/6mICnoPS0H1afUeFKldcJ6Cjn3uqCX47+QD0LFl
+TcWB3wIJVTbmmz+h+yddQemN+SBiNt8jPxxPC359M7Pnyrow2n6uWpFjfFeLlk3
jAgQmPoA/HaIeqwEeqkIbFYDK/CeF54zeYEme0YiBWDHf4tcRTVDWtgWCdY/ty2F
zSMCsTjaudVzTS+5BMCA+q/66nfGEG8ZgUPMPrOs1rNROxHE12q2RUI4ERnw1nJ6
1iBdoOj5N2pyrHtjokHOszK1Urc6sGw28TKBb/AJ76fmtqzF8faY9UAGgDd39GKz
y7eY7GkdK30SIangKQcgKOYkrS59r17F2uMPr3SDAtruQUp0R6DthtBfXH46g7pQ
0KnwYCR8LZAnjF6Fn5xjHGxOSVwihSHE68NH8lBxrZyTbY/55LJarQAedEPIz0Yr
E9qVuUiFvP35Z5JcsrfmAtIy+OES64lx+3mvLSq/R0TJN44vRoi8Y7fr4uTOq9Jy
5n44yDuQvi4dSAKCfIATI/dK+3pYcwiwV/3EUaRbYzv0kTDJyeRObNDTIoIQbPt6
EcO0LzRhEmiB32iQYNWpY8X+xvvu+MccXNzBpndOFRX8q4awpS9OIZJxw1s23Esf
U1ImphdHedpFvWvzZGRXN3yeVMQh577Bm5rjyS+20gT+8FE+DmJDYixpfIIspnp2
32E0HqmQp5FBgBXgms+NCceJStqjJFYvpdy81yurx5nQETqJlbc17xeL8X7RnQCE
U31y4b2nPj1q1sH/99yZeJ++S/jK4SA3+OnfOz3NhBcPP/ZInoDucQgB2Q1zISGf
7cwJGkLS+spdipIfKzqjKIF9LpXHwBGbxYhvYrmOHzayo6BDBO1i43wD22FANKOQ
YGsFIKcDZ3y4PsvRTLy53DJOqWJgoM3m1l2bfvCqEjl541KPYYeQhVwWPHWHVbEC
dUbSdbgl5LmFx5V+VZoEXwMAymXI3xzDmbeT4Sn0rMKsZHoGM2IaVp2ZUnC6E6RW
IKb54G5qViakfFPzwThTgZ6guD4bighRPGLkv3ZipmszNu0SRHToyL/DP7WuqJUH
Jh/Z+up5a2sEsDHSH0XYQbp7x1tRCNCaFMEBHcyYq75kEbLQuS4XTVtoYkvIZ6KN
QBWcEHKqX7PR9IJVMttgETTg/qQ3zdcOAhrI0o7ysyjJrZbWKPm10bV+W+X1IEgP
4vEtkRYpelOlZONEjPyjcfjc6dc/FEGmydmEDJorhDIz1t/atxvcr7ujG/GeHfba
5ntoKLvflbpDAAbSjLO42B7g/yjjdFFWPUTUk/IfYKp527n5jRMJc+matdbL7kAD
GiSIzmjPgBxJYFoJW8OBUZBuH6Watp1US4vPHa6gGWN0PpEm/Wugxqq5GUiWnnW+
mVn5tmF+ylpGJBCUEksTfzJI1NLbantrFEh2bOGsDPrvThWZl6Cjyy7YpRZdLpA6
5Y3p61bIS7btoWsOgdCBO/6f+0Lk6VJYce8P2E1c60dKCHUcUtvP66UQiHs5h5UO
a9tcfGL2Hz5skIuz3hBwIA9NmPJwi3UnvfLV3MGMy/IaGu1ok0Y6QLgYA2bzcbv1
9jco0we2bi5xd1ol4qdUFyR1dr7aB1ltsGRXvpKUANpBFwMVsa9+1c3jyI14q7od
LyaDe7nuRSvj/Yrg1zZLM9o9HVwTg+HjSxkYRN5jRiE5yV+rxoNSvHHw1LxhnaJ5
OMLLyBDlExwJ6MSudi7qXBmtUOXWaJI42uS9dMK6AGaMj0qfqwyke3DEqVnc4Hqu
OdSrN17g4Vprk6cVFdx5v6NlfFQ4J3Jh3T8envbBoiE3mJasdqfJWahD7nO+QoaX
kqAgCWxJ4L8Sh8PIhZhG9DG2xCh1GB2+TzV19JIdzGgiAiiNCaTw+Yoc5m9LjtCw
RTdQC+HVXWYoFUJ/33tp0vAY3OgwoQPreDwAFi+9OvVE66nuQwhgV7updCwTEiMr
EFR7brvC3UEhkIiNbWASfgdu6z0yPlFsWiGb0vnD6A4SEnZDhVKqEJud2XYxXUBD
+QIT9zcufMqXK3xum5mavGYa+R0XV9oBLwOQC5moF2IoHMuiBCdWEhpgQ75rxsqG
F0SI7vwiH4COUFP+PqY6dtj+vjaokC03gPa/qtZyIi9D8n8GkwCxF9P60+Sd5mWp
orAj7ZddOwBMrD6whWmXLKjSxwnE2DfONuFGySDDIb8QSs3wNxXH1podKDZ7EWmd
0rVELagGK8rR090iB4uCKQVOjbE3G2CHPcHRM5+roiWFqSbruiowgXKA7O09O4Fk
Ka/W5ADUgdTqsdqp9xJSyBU63ssTiTviKiuQzqbp/NfESxttoXB9JxQpdteE3Bhj
s8P7bUht48ZBFBpTgHlZZhYULz6s9dIA6CJuyhlRV9Bzg7Qkw4uuZKAaudCAGL2r
XXKKZbfmGmMvuUo80J3PYT/EpMeAhtzKgB4B/T13GF3RAiU12FPtvbfpzuGANVBy
8uYmYE+H6yhwZoDm8dKa0E91YWRMfyWU6+50FYsWug8UK6Yh9LPcihmwpzJ5byxV
nunzH3KiEz1Z8kXKrF0IWAKyiAOQ15ucww1iktEkZWQiV5dOl9k005J2+sJh4oJW
plIqgZ7za+FT6mKe9dYP4lcrnGB1PNRFKzX2rZaJN228iN9IkUpC1/I/RlLE3nGM
PE4BcMEf62xtLqdZVWHJzKH7o+L1PNDJku7kJyBdOb26r/EdFrBsZAeT4XLrWUHI
6gcwbVsaI81e+7C9incdQv18YJKyGJAbEjBB10cBB5gj0ewSvdZxytQwMeu75+iX
A+PZzpijDHkvlXOQUwF+E2rAuJ7vfiDDtXaWC6FKhGZSf6b8jIAan2oOsDqKk8qk
7j7K58dp8sw298uDyMuUzCj9PucZkiu9hSeN+2WRtknxZ95irVnr2R3aB06NP87X
qJRap74L2lV5AUKCmymMOi54H/T/MembqVy+jt6VML8bmyDvkqaqHbuJpngWl9+G
GJdSDU0BJZBGtIK83YATEC1pIB5GBvHD5LjKbWAnmRPYdDNLTv48ipndCsxy0DN5
NxogbyrAxipWvyOHKjpUg0xVSvOk3ApKNo0OvETfaGDkmtF0U5NMCPEA5inj9/B5
i8y7tuGVG/em5ut/GwHFPUZeVgFsYqNlFibdmqdIwF7SGb1zZbK8JI/metjwuc72
TZaEIF6Jvq1cAnSnFEM44Fy6KyCiTJ8s3edTUIsBLz/geU6fG2hEyXy40pQmHeIx
ImLZ69ne+a6UGULlW2IBiVdnFO00rA2t2uZywWCMOxc1peYTwzB0jCoAmMTBFu0l
wTlobM4BwshoFO88bBR+4Uz2RdbGC9ddHjFQekZaC6k7kZ3v76o7IYgXIczU9b0l
VVjGM3QAkWOd+twtN1PvlzFCVa5k4dnq9ctGGExarbQxrl/KjBYcHG/Wr6tEWuhr
lg31bNrLqTCQzmW804hI0MRp5e9KFs016pnZW9ngc6pSaqIQiKiJk076tc2Mhoty
w3Ya7uALczr1GWnhXujbPguLSmuGv/j2GFMKMCKaXyNozMNjfPVyl1dh7pkbGQEI
8f5DaXrObq+uepQL9CUXCXEtY//GdA0pRQkhRtZ+T/wcICJPdIDMUoopOI9Owi1c
p7vHUSzXOMV10KvOJzgJxaMG4mEvmSLhin3RS2ITQ9A1fMVIxnUb7a8UsYxfhgZ2
/BAc/uM0a1VjeesaCOANzdw9pRY1k23jf7Vf8CrpCH1DHxPK3JxoHDC0RZk8VTLT
bOiicFWihgTTSGRyAT9ep/iy0LGlf1CJDnSpwK8mSwczNnEccgduY6WZA8slzFmx
jOwUudDunjPyyIY8ZPuvDCz0CrVbOo8gbiWwMw5lzLX3OxIL8KvhHwnWydh7LfrX
Svt99mFdU1/tJrvtQUm1kAU5bpqOq0PRp9ZrfmE98JiUK7KZBOm6BmI+iP402Jeu
bgVFQ8m95X8jmuxWcNy736nQKHGhQ6JPRehbf0O5kisonSeNKWih1Nn0LrP7plwR
uQjTpeGZBBjS++wuWIUcYYFax8H5yLbBeHVfU0ErfcQT5J6/pLs706LfXIFdTDoN
wef0fjZ4+sZGLWSJlDK2O8Es6s1QDs7MW0oQN3jPlhXE1z0JJS/TI+4Cyo1hgbfd
XS2QsNbqJKu4VFA6CqkUtZLol6v2V7HflXtaZ7bGmTbJGLxRKZUalnCULT8wkSEI
/I8uUWx3cG8Hk1WYC/cfC13nk0u+SBFD0bWJCUC4wc6RaNQ6NdRltxtVv1rlHN46
3BhthqaF89DZOMnDOZjGZSe+CLO3TksXTpTrrgL9On5tRzR831sO3053QBOieHtS
gAn6EHzZwsRz5H94G8SLiF/hC1SLWahaq7VdNMom0snDmhtN92sTEGvZ/ln2hYva
e3wZ6+OPF8cjOr3oZl3lrMx+X3/MrxcWXLnp8DgE+Ro0lWV0vEeVmCe5/mndYc3/
JczRKzAqP4VNkki2ajdJhlTYZ+g6BS14FTwoYVgj2jlmcLV1vp1aabOJT5npDG6K
piPRNZ0UtPLSwbEN8V+UBDuIwt6qbAUAEI1/VP0rimHTXLCk6VF/IaMIKRRulRg+
spaGglWa8Jzw3JJNjNkX3uR7AjzsKJBXsP5iiLcZmFOqVpkV5G0WPG42MPmy391t
5MVIXNcmgzL8gmuwWMAegbFWdTiJyxHiF9v3qao4EyWGN74IZ4JotEaxd+rzpNXl
VZ16UH5G/CNVfWLpnXuh5gfPRo3jY+yfzfaRz9JjovM71/PaA6gjLAVDKcHsn/Sv
ndcjpWEKQwqYmMeG0pXSQBTRaeC6zxsf2ap7NghrxNsoM2Aj0wKVPbBhfS7q5o8y
5TXx3mvFzK5oFLWkhXQmfJdbCw5wkWsAAwQueVW5k2Y6MfmkvhkyFCUQNquDLQCB
Ra8hQFbe7dIa106KoinyLYIrXzxWOoFrVigNyqEzghZ/iiSpichQoy6MjLtLAVr7
jL5txKKXPqiMJAAG0aQMbPV85RNJjbNEI55/5JwkmYf+vFxtqNIh9aVEdIz/dMb2
30bAV8YUCS2iJNEmxs+DYHVuybVj539MbbQPARbTFoPpEFUemwkuYPywmlXQB86m
up/RR12El/h69J4VsdoXb4x5qVkjqV+u4AsRJuwoJikoWRZ2pElfXIenvw8mdl+3
FR8PPl9Ob1UjZUHApjAm3PocRyMHy4VLGKWwQRJo1K25Crhc4rk0dPZwM1k2wV0x
UEJ9dyGy2XY2EiAIqEYL0iRl3o94chcG1CWYdJgVogyh2UaKxJi9oKPboIMdUeU1
P5M1s+TaGNx4hVJRQZK/wTIePpFA22Jn8xz9rgwJHVy45Lv5v+tBBHjyIXdjIyFQ
2sVtvMJ1rJQyOblgOaTHcCgJDQThN8p9TiSIz3JcBwiIop8B1//6fXStDZMAM16O
48ODUOEsIYTOgaTGEvPlp+P2CwndV3ivfi9Ar+jFT6y8HdDn0jKE9dhY4INDKsnZ
JY6oK2DnJQqYKlArvSC01eKycx95Xkr0AB/sxflaVv3EcJ4JNDoM8M+h9Do/XT2+
5PhEMfc0MIL7hYGru5tCpOAqivfotUPzCUeDpgM1kvXdaEyAOL/8YgfOoHCqqEor
yOZFVsevJ6iDiocmtAcCbndqbOPJfxdDoqnc2EmhSIepg88BFm+DetqQ4nvRC9I5
n5bT1+gVoX7z7gqYZJZtbDVRC6nILYFKJj/01sg57+EnYyxSiwM/k/XUVL6wx1kd
rKHB4N5A3jOKLCnS6q01hxBUFx3DYu2uchz83HCtCC4v9gLD92PFYaZUCwvZC4cv
s1dtoPAMSUVch1qBHEWbWyfpnqnNW4AGfbzfQK92ad00u5W5xBdIlMfnkhSvNdRy
K0Q937yY+nfLZyMHxIxvJLENxi1CS4klQtwi8+jCiClDLz2bZxSMtRkJ2HTwM2Zb
f0/DNwRFnOdjY72MZ27++bxoJr+pHcwA7QA2aULbp4C249ZE41x73dG65ZDP5g6z
bZzC8xfiAKEKoQr+QNIfrWYetp+2bbbaGNaPn80869bLiOEYOeJwto2dKVHASa10
TLCLz+m30F8cUXJdCnnet3bEgD/y/q0+IUxzlAWD/myjiSJS2QhqAawri3dvLFtq
Vp8ZOcbo5liXFkB6/KrbSOV01SxDbnYfhopDKU85aroaUqaAkg7n6yEwKaNlUcCE
ZLteAKv/zF5/d1ueU7BpNiVAtnzc38PEqQqmmcj6i0LiIiomhUm1JRkW/2z0NrQm
Xz4Hxux+VYKdXBiyOrpQd44/PH0eGv0nosOErLN3YMMmaOWFPrJjEOZRBzMHPWyM
36FX5SW8pNcHl5IVIV0g8nbF9onHY7GxeG3V8Nw9jkJq+J7VwAJaPHPGK0m15E+h
mZXU7y2R+/FmqxmSqVVt/yZDjDmYNJ7TsTOwNFQKFicXqpjhtkTRX756FL1WsEGo
l9oM3bGYMUGIIUgiFgzEszATdmctNztBoQkGcXCxzoLYAKM0mdpZpihiZtLdKGKZ
5JsJW+DapXsLGnCa3hfxO+XaLhu2zEPvw8H45pTZwSMQQ9ILDOUPAIHKaVvHTUCx
i+vdICbC2YirGtwFvTiEvTuDqP62zN7FedDBc4yefH3TZaijskwFk7JlKmFzcgRV
19c4RHpJY+mPu8mq/Gl5nium/A4b/Cgg2k8G9LImDxpI5gz/SU/WRWmBf4RIZq44
7unWKvsc1JWpC2Yr2bFMjWMRn4xSbhhMsMWATuQebgk9wqR2g/zVgxACPlVKwUvN
K0Sf7nqBblkN/OHtfK3VgQgPo52eMmuqEbEn3n72Z+Xf1DAm2YzOZ9SmghEqTStP
8P8fU8Ikkxk+xCJnVq/zI6cpwLc38PkqY6G8LfJMAx3RmHsXvRLJhHTMvlVBeJwV
hUKXe4rxO28h2x8xy0gmlFghajaAVFnU3C202YVvl9n51xpKX6jUiVZbrG4UXyqu
ZaOec1A0Brrt+dK/jp856cuxo/1MnoWoN9XGNlQVWgAV1oiC6ZY91eOfXm5yJCPj
KjfhlWPmDqkNKmAEvLanANTk1CVJ0odJmkERuf0nNE8oYhG90E4loc8/A6C5qixx
Dv5myF9ELKBTLYOblpq+CcNbFSV5ZXjlkD17LmF3G2brMU1gV502uxVji98RNBul
FNsSgWNS1h/DjzqHWnpKLycoiDY+aRgjGZzINk0sO2QrqHOx1PKW5BuTFiao1sU+
E6tUaivJKCuKdPVV5yWI2/UjAw/VQ0hjlSXP7RfzvNQ1Ov4YrjzEyG7i98yipNnW
LBRC2GMmek/9nBNaAkGncQlg1MUVh5mjVzK+AqI4XQ7FEYGD00tF0/O9asBn546K
gbH7RgvAoDutU9uWdFSRqa23bjkxHbn98AUhJtp7IBv/+3IgXiOvYjtxQZ3zbRMT
J16QWnxQSFpLe0aNJLZwPLLR56wuI9s9oBtkhi5Acz/Lxl1mDjUywAP5R7hXgUcv
4EKxXSw6P4bteRf7n7gAPAC3WfT14NFyqZpxPTSFDBGgVNxBq3BW9EFnYJPOJkhL
P8cE4HMx4hjN1OGzg9Inbg3dDrcaReODUvS16olI80fi0WhYFac0YqVC9crTAAJB
ur8mYvDocrBRI7FrzcHshuN6yhGsHt4/X2K71Oo/3UaYVlJMtb5A9N9WamB8rC6v
t336cxAAQ5q2zt982G1hyFrwzYHH1fjdsmT45PCwlXpWf6rnydwSLNkZdsbzhGzW
VQ0JxquDMaA/BNZS3bvl/aT7kWdvGZ+p8gqNN4+YoEdMWzaFDMsRxvkNMgNDIINu
/7JN4GGSAaUOuVXQFvaPYb9p1RvqU+wYJB6Ck32Yt79n/rkbY/ZMGDp12TS4zVAm
HcMyY2q1FmwppXL8g2d6mhH2jTyXFWhTNsrfIKn5l/tONLGz0M4YtoEfgVl5Q+cN
ZPlevX3thbtNYclWjAvaNgKbo2GRD6XMA/Soj2VJYVCd46cQEaW3SKWPWjJo9oAd
X0jc/BT5UAUi4MRVVZeFnDPKVKweBhK5lW2b0BKY00zuqVQUCmlp+Yz0mqPHdUvD
05wlLi6hbKXpq+Prg7XCM+VJdfEwVZgW2iuez731vZ2ohdt+tQsY8MrTirX8/Wps
o11EbXewO1Z4UOQLDnt3/PAK1JpQHVJBdVOfhDZq3tdNghth2MW823YrYVDPH2zS
gXPbK7zNsT5XnhvxO4afmkajQMN6RQu1OK3086aTLfcJR25ghnKptzKQ2Mdnx0Gj
KHAgsF7ld4QcVIvAvcodPueoEAVu2SOCGHcOwU+Ir9+GDv9wTS2Zma39XNWg76ni
L8UEygjiMzXsXZmBpYOxHW+wWZwQoPLIE4IfxKVAcRMjcXFmjmHMDhik5yxfrT9J
34F2kaiLx9itb9igpeMgK21mJ7QKzYg/BptnAlS0O0j9Dmf8a4NrfRyRwQTg/7o6
w/ggJRDIA/r+4vc5yd2yZK3Setb4oT94xaCenwxRSqudNe0jQQ4hMANGwlQ/U6/i
r3NSCfDqpr8p+NHSdujTrQrC5RYokuRujyGvZ8asVJLPLCllG2A1/1g1SaNtjs1J
Qz7I2LTzVW3uilYZgdCZQ9wH1D9dArtYbO9FUfeBNH3dezNxdwfzC40xeYc6bIVe
/Twv2lHGD90uG8Shb7N3v2esSucc5tgrC8+h++jEXX6NpDJu+/g1CsjSiKSzZfl9
jK4OD/D9Mndia9CMvR5L3+eez1piaAI3qIIYPeEoLWbjcw40Gky5kVAsdRkl/Y/z
aQqc2yieNjTeCqjKpT0X5H7OdOwudv+TbYrQtwrrbmpJ9dZ100FV8/0Mv9sBw5qo
Mvff+efyG5I5BouCGTrHoUzSFPNObZ4Er28J6N4yZImZpqfH2krTsb4s6mIFZ8ML
wL+M8KcRf2QVqqGTbmoiWPeSAEE5piPq46r6zQZ8grQH3Z5vXn8n3qx1OG588sMi
Z25YzX/QFLP8qlj1Tc0VW3xcJVi1LZyfWvWlbfhvTIYvfwcN8XTnl3h9HLO/ax3A
iuOsMo1pE1O2Ok0A9GILV+F8BW5BDgbNrQF4HmA+XTrm+UCGeZx9108jChLy7o5P
3OcjoLhm4iah5vNTrz3eJUSrlU9cCyvZFl6Cd3UwyQtwcCJzdMuSDWErwqTGp1Uc
voc4IjWslXRFbRQZkatTHL8zYGlUOJGyWdwNNRuahQpSYjPWrp0yIPTXvf4mQmSb
IxcMOvVSokD8dr7tm5BkJXR9wxRJHhFI629AuGFvG74CcBiCD0yOAxLTUnJSN9vH
OhsPr0wz8UCd9riLbeHybyjDQyeoltodfAri4cnRqNdR0CLJc+KRMx1tbylDWCLU
udkcqLQit7JAcIJ7ni8ZoSLmKW3s3/snA90iWOzFQE6SHLFF76rscMmSbarussY1
/eppN9x8qUk5BaU9sgDc6VG2LmtMvo5UZOKaMDWqFSMpJxneAF0A+N29YbMhhPGu
v2x2mVVFdEoQj+uq8DPXUbaKj8gnfmEiUi3nt8xKCXQWdLqKM0GiDk0h2nCoui4Z
WEi95x2WgkUH5Gb9f074ORlAFRaFF6H38HykkwWBrsyycWoJOqqvJXz0SLEv53h4
9r4dEfCTwftG+sNSJuXP+3tFPGTZRzJ+7k+s0jmBipf8BDJg2hBSD2LSaix5a7+h
xNgWaUlq/Ly8IwKL+PhR4waytudohfyK0EltcQKXTx7ne6ngeXWT3ufSEJnT9Av8
p8iUEJN/ysEwoByYyfCbi43liHyxHV670aj9GrGDMDOmF0YqlmQnOdw3tWkn/YfB
kyEOhM7fbc6toeM/8xjy5xnail9KQbkBhgy2OGhYcIz8Ju4/JuMvBIxsvDyVfVyh
JKvdiUdjhmP4vGDnMmVBNvKVbBNKFYYfJSIerLBH9q+s2BZlI19+0q8CdcSm51yZ
5P73XDCMNK0o4TpV4HriH850V1yElUj4gVSeJ91ZeCtWNhXLjALjt0Zobue3nbTk
2Wy2wrHp2zPxq3r9xLMbQ1NURrnP1Jr9yLNd1her/qfTAmhS2fn6EF4s++0Q1eBi
kA8H5kGmPqR0Z3G35DikkVIYOXWQfZzH7N9l8Ttt0yWwbFJTvbyE+pSnRJeiXuMo
TFcxOqYHNiYJlQL1IRywgnqSgiSj9fjVtpYFzoJxNXn6tuVmUQRql1tJ+wnB9Mbt
nlWv7oLEBJgvPwLMZ7frKARp+I7aJxXAI4SpRpdxnZz9mZvohGkECWeUUkI6Q/jj
aoUNB6qTjipVlsnuD3ic5dVUoSXIIO/3u+qNQqpYZUN3QI6SggtDfTqT/LX6lhCd
rcGxBZXzkJ2d+ARSExQPMgoHY7UzYyt58Zft4Wl524nmPUqWuAG800wU+4zPRb2I
uQ3jfVipDLEYWe77E3JoPkf/rC9JtvM/6CPwS3lfwL28/Z4qh9jEzJKuGrJ0ySvh
wgCaXK2w8y8XPjojBo5LdQFgLMcO9PZAsdi8s9vAQPNeDyR/ILbSuq7FomanVvjR
mIZY2w2O9/9/ItAKTKLAs6U/lZASYZEzBXXMxUH5mxSOelHSO8hU1XZSnDrX2Jks
Elv9eB48NT/K/cBC20/g0WzzkZDlBFr02e6pB1edz0q2BwO7oOEvdnGia1+FYtWn
9Wl+QqeqhNa/upT//VpGx/byWoE52aZbNmS9sN3UQECdvSNFzVb0Rjg03elq7+t4
kjJKxZDzR9Wd6i/cPXefQ1Mgp48AIZ8sl4k3T77uvip1r6WnEKSSVvdKP8NGqWxp
Eae6nt7oLUdXdg+w98CTGpZ45o4OwWNnVkjfiXTBCsNTYOJDypQFE2VWDAqrfgDB
TSln+nRRpga5voYdUH/zk9bMwGYKUmIr6HjUr2speVny+/xbMRdeHa7C6Ngze0B6
7JuZnB2YuO8FkRi7WO7Jf+R54XBOWZIwRjUMhZUaa0ds3BxfQw+ozBruBcPWOwfm
uEhBB/rAXRR5S/W+6fmy/pFM7nxOED8I0WFcHi54cC0YABVnQ1BgpPvpoStBSBCq
60XaHbVVh3Vb+9xciZIRH+fNCqguZiKFx4XNLrZQLUxHa5D80V12CHuMLmiR82DZ
zSdRr3VDSNfHFCXt6n631RXJ4Un+hCd1qIx9J0nX0LYYh4VVwjGgbDuRSdU7oNxq
VK0Ynl3vPdVIYx5xlsADRcJ4QtV+QdefTMRKHKtxC776GDD9ya7WyrVD7UOFENCj
T8w6ClTtXhpaULltyVg9NQGIN3W7jiqyY0PZaQ2U3d/DGpRwrFnq71pomSPBg67M
6Li/d2brS+DxXt61lcqIjlDmzcE0JNSPnQMY7f64oJ4ctXZ2rtAggVHAlTL/bt7o
niVQgf99L5ytB6obkXvBx+9tu7kcecRmepOU3ZEiTe4cj7gZ1v2v/gjYnqAngR+3
r1Vy5o/+w8xkHPhICHDPOEY0dlYW3wlwIekoaQCk6RD/u4e2kCt6RyAGh/K7j0NP
KHE+5Csn5M1KutlLp3UshG5b9oNAtPnRsPg/R78bWhYeOe6lG5aB2QIKYA/Pqrdf
qz8za1C/GN46EgyLQORrWIcuseDPh+SoBIzI06V8nb21kktdtuZV8laUgrAEX1Yr
ckOgiuaflmqvQjLOmAOoJA3KRNA2lHF1WgaJg9qnNxHzCNSazfBPA9NzJIbSxfIi
o5wbLP5guMlKA5CPuEBOk2QpJD0nGMNzbkfIq/UfkWZLwdFMXZeBTJvfYDhWUgkx
4RAcN9irT3hEgNrws+EkS0XyfNlkrYMHr+CrkrsAWK1gM43bKalEvQB3+vAaPtrU
rnURu0QIH0MYTv2U2gblNU0F0GuE8dT8mGaUHeaJiU3HB4wEJWK28/plggUl8xFx
iH56ygXrugufj09F/IUS6QtZ3oe/5wbHQlt0qwBtrn0TBwjqT5BN+bNfpXQPcStE
OHMFJSc852bcZOgy5pCxP5zl3KUpKDfI9jHGV/ud39N7rkZ4lihDnHV9MAmoPkjV
085z90xLunRIaxq0CUs1S7ga2qdngsvlzuBDs+1t5/bsR3OkXcgiZsssEYeUNav2
EBBmyfInKYw5/q/TzKkQITCwkbYiTv3esSXZ1JMhXwy2W7wHxcA4T7JhGvdzAPhn
RByxHEDcy70I3gJzQZ4yDNUZ/ENzA3Mg3MUuI5Z9luKFjjuv6Q6VwPzR4VuVUReP
cE/9yfBLqt0Bf58DgWa91BEXgOO7jGHip+EIoqZ7+cnmFnmAl+TQRVg9dsAzL2vy
8oFMAGM/zsgJTX8a8RuQ5EMimskil5BdZahUkJG2qLygdlU2SU+zi3rx7rl9vm21
M7dRE7UYv4WC7HhqV9OTYKbNwHQe3NhhuaneaOJxk26GsZHJiK2wUHqqfx5T2TDA
KoDAQjTCNzZNI8ElJd2a86KirFq8+k0JVd2MgT5tEGAAmlXH78UfVc5fGJQjqMOK
sFKUXklMB29iw0rXOrULxT2kD2rs3YSRKpYvaVO3xUzxzfLL8hxhl8xd9fgqljjd
TjO4GFZXh3hAhQG++5PACTOh6IRstxDO6tI99uxRJlnHR6q9gPMJV0QJKHs4YszK
UytpuG51LGGndjJtNWY7kFW66JBM2rJDguefS5a8IiJpxAluhc+ESNSerloOqX/z
xLHQhEWx9NbAkWF8Ef2OV74Hh6Eqpo3wETxQkKKf0komzdm1H09KTlbHmDxXK5pp
H3p54LOJZ6VQ5Op59fDUoHIeTrIYS5AC/q5A84kp8256sFusKLBIdmB4QEzT7iSv
T6o3PzFU6M9ZrBAvVZypIJY5KS19SaLdEUteX9MHldVZQ77pn83nUOsN2fr0VI6J
eg58o9CuoJu1sME2q/TPEoT1+5RKaigjgO/JKm8a/YclaVgU03U5zbUKni0Vn2NG
pJlUhXxOH/vfdGVQ4b62cFIMafLKV2gtR9ZT8Lc0bDt+Cwcu0/vTJ+uyqHsOMj5Y
/lbxAHElPk2nUC6fMfmW70Zok01H7kDSW8CY9uxMoCnUmlaN00ZoNsUKImC0mL0r
kTfGFGTsct3J9tgjdnzTZNTIXq/MICB3RgERwmgb1FlH+11wbIEsyAhPmnD3KWh5
UaLx6SrY6q3FjD5MmkGJG+7VmtEWeIb0Q4rrzMPLsmfAyIq8EMtE9CGssU3EGhZr
79N6PMAbJVItKkIeLy7V430wxqJ5u5k+EII1iT7H2JnBl9leOq8fTul6X0sXr21c
D9RV1j32cxIc2IJh5LiCfrs2raL73blI9uBVjbfhlqsOa8uab8RHiIBjmgiPZs27
LScUbOrby0c9XIa6R7mMbdrI7V//y4LmIuu5P736kwFrJIN+R6vYSqsKrsCcQvjL
Q/h1arnnh8utVrcs0JkeOekJ6/5u3wyYF/Pc6j3Vw6qnEOz3YSzDlaXqHbI4gu2+
qK0xjdU0nqA8hjU1zJMcZcJlO8IYa6DFBAKeNnFdaQjFY71mwmS/Y6XPKDoY4lXH
1RTfON46aD8peyvo/emRGp2FWcoG0V6f/p4ZuZBA3sIKnGYNXJIaa447zs0mUyHW
BO4GcQpgeCkr9HJBtIw7qk3KZTJ6kIlC3w0BZyCHXCvlOWCODfQL5VdfwRZzLVlO
kTXWfOhX3HGiomwi+ShaY1UvDwNM8SW+FMKTsBIFXhYVvM5eKKqt85byA17EDQCA
Xp2NEua4igO9zBG4Uibvn0CQ13CHz/kY9StOtXqmp7SSmH6fcWgR2/N1zd24HJAJ
q1Scy+oxA1a8B1iKsXK3jcmU4R7zNKm5bqgRbaIRNNdDN7vn73JjCJl0AuqyZiwf
4Xl0KFtffCp4qjO0pa396lMixgmLhYALsmRHD7qIr/6v8GC5kAtOx/OLbkSqxXoN
T1YjsF9Hm/EuobHqCJglKHDo6ZFCPYLvMi8RQLST+NFK8fmHAwwCufqrqI1NT6fP
N663xnPvIJY6NJDtxqR+XgcHiEShoGjVpHhQKkH0fIIo2HkE3F6UiQNP/tv0qvA0
VwP1gaYnW1KK8yw3bDIVtaSDDhZldWgr8TTOh8gWM4KpGMfnhQxu1Mga0tH5UFbo
R+/wQn6r2jjRph//8aOPaTyn7FxKvwnOjK5LJpIv91roTErq1Fj+P+u1hX1okHm2
vbPi3nfMG+bVH23yqLcMRe11g6wLuiZNGF461KdIi9pwt6Z+h69rxVgWEOalE6SJ
YKEmob8wtslkWWbgk/xSjDCanKwKIrY1yVDLR5WXviQM9I1+QSYLRU+9y9MVpNoS
XciabjyP4AlP88aLbLGL8Afv8zvxXReaRymC6dlqqh2+aM/rdsxKciOeIAfpz4mE
/FEt4moQVu2nnacZ7G1VWs/8tVEBgA4jHI4NI9XLDneep1aj+Y3NOaE3e2wKggzY
xJeGTXFlCjs4UjSgxsygTe/HwFQ6gsvum2D6yc5HqzQXED0jkoalfOXNhc/EeXwO
mGZGYgOT8peldOFNLsjou/zcoUPWdjZMbnFghdRIEwHDRBa3Ei9+pzjL+zCZ4jLm
lJb251dqjhwE8BzUKK8jsBaAwhTWh6lzNU0TrkohtmwwsRmEaempkMD6Xibz6Nqh
DRqJdl9unokqs/H79e7SjKdLFpqUVU1fFZNF4+YcTHP59Nwp8PIQAkxAyrzMYNDm
CsT1muKmpfFhFJTpwppnWITuvoYofKqRXgPnIz6FI3FqODd8cbiG1TZoGP1iyJJt
YLvpLYOf2kP1uAOrqeXSbmUTFEfGlW+s9hJ1rLPlljse5A4pLgFJeLLXk659YS7x
ryERKyIlvttMB4q/fdxW5CUMOvfv1BsG8LqMo8r7gdhvU1N8s1eimX0WxzAOnKxi
MEyGVJL+/EFvxGvrbmwXZSkAm/mc20pH4mgHQPELKsASqeAfVctPJgdhjvVbtt/a
1ir2evCF25Wqsq3W4ZiGWQDiHQDe4cUh14RGtTaEgZdYyCwprgPu5frCb2xJvnYu
nj7kTXne/DKX63dv88Q/Yd43bUHdfB3CUvba73OD+UGimzzmUTV5q+0ErCKZE/uM
n2JZzhSE5PjNIo8a8VETZIbro3fYvirzHvqAXW+E9fG2aDeER6l0tYuJHOsppCz0
anRiMo1uHGL4JkNR6jl5uPm+9baL6JG+N8csf0DzJr8JmxQDbLBOzspcZ04ib5zY
Odf3WrbYjc7mgkfsFv9YWRq/dYz/m6OeJg91/fR6DhFejk4ZyYKF2o5r+bpC0D2F
xPL9OCQNChC77R7kh+8lPmCxj916+RpoI5nZrsBMY7rkdB+dDZCPoL3Wl4mK5JaP
mx8Utx+aXDX7oWGh8KV780/zfOmo7CjLzcoA9Zuij3v4+vWucvvXv3ODRXoJxWh9
3ck33VQdq3HoHGicOHypnjfo7zqDvJvVeS8cBfUB6KWAsvSDfuTsVaWtD9zcI7Ep
wXxKDrSvDJxeiFLOidWrKOGAQJ2BLNi1Y1fHzsNEazKG1TiuF2qFsd4DkALvQr2h
Y0sUK6uqDcq5Pcp+TWQLSyR2NQ0nvu2pmQ3Y3h1YJKxbkLEhDTjZeBLcLqgDcZfH
wOBxUc8FGN+peAneOiadGxZZddya6iAmhcaZzYOqMGfMXytjAUtpcLHdjG+w/b97
J9MiUwNL0mKxmdaPRH5Lfb2doX5NOrFiOJs9oxjBTSewB6jD2fBMArPkqgCT50Jr
gpd8Oy5kxyj6CjwQZq2vfzOJMnfIY3V8MsghWeOgA+rYcG3Mka2tMK3ke+IGLMOw
6Mbz1QrptEfuZknyumyJNzhu/TUdDNu8+GC4sb+o7XBa/G6EHi8he+mAMDeVZeug
x2j0KQTK0Zca1hVMQwMYX81vCun4dh+TDcwFKqSs/o/hLJkAg9S/VX0R6sPmLYez
n7ZOc73cksgsygSJJ06I/NztUn0xYRndFdSq3VFU+3A+nFnXQFDKJHCYhSZH0XZa
9ADriFDMu2ZftvGAFZZU/TdAS0yjz8CRxHsEhysvUkrgBfFQqWpGe2xtS4yAg3hQ
1Z7E4zRFhOnka/MKk/AofWLxSr9emg4VSxFt/SxzMKUsuGUJUHcg2MD5FS/bU6nO
nigEy7OUo0x9qEydSKIZ1WBduFQl8ZJynJsBBzt5uGYGgmo2cM5jSKWNoCZv6DIW
mvIVwfk0LOTwzxNpVtQyHQrYpfZlMWx2VaVRelKzJ+tSDrY+eT4bHdDxM6iEYouL
dKj2LdefoD+p7LrSGA7yevQCJ+kEO3s3CLZg/u57FU/5L6L8Vp2xPmDtviBZu/hX
lsjWzZRGAWK7GUr5HYst1VnyWwrZ8Ua33b1AfCgbONU671r3iofd3HYIb8yQ+SzZ
73MT2AmWexcXC9WGK9008nasjHMW/Nh3Zy0i9zAMdL4GRKEMnLetAvKsaOsfT2zF
A8kjqfR4hPyx39v+3uQ/1N35E0Rdw/SJyvKFcWfhyOTeuTjdqh+AiAhQt2AqOIIe
VxWeGEfxTDxzEBMc+qxFvD4gBvEEcqn5Pu9bhD3ngRNNMhqiFaYT9qWjFjSOFI4c
+wsHHrtO0Uq5u/LT9bBtTWucxzaHUALix1c0tv1HjyUlBoEKk9Drf+8vnPp1cdmk
pquDdgKS262lJ5APa3ygARzr7KnQPgYIIkeRkKSXNVQAnat7ohMbUWcPXIpM7OJE
jPjJEaI7bUd4ju2VWbuQbC2Qy/jNdhZcWgkCKPpZ90FNtJZ3akZsmN1s5NuVfUjk
livk3K5kXVXppMkfyLVKQ9wK36lGHZ5czY4IQB4QIwsjMQZLFZ6IV3whNWoLIkeO
QIuXIiQ+DDwVsqcPgeN/5FvcFPLXiLsl4jnxDm+0F/JIUp3Vs1iN99fRs1/5LzQm
Z7Vkd9tahbQtajBubdQx0nAfdf8KRHbNg0ta6CP3oQmEVapfgHpOc/m+27zutaIn
v0yvniyUVwMzcSzg7Y4Z1R0tOy+ifDz3qM5Cmluag3QEH9tuNhmAsx8UL9ilKtmT
oehUc3sA/LLQ3u6jTrtTYgqG+OzkXdDcE4nnT54KtUrJBqxHvZIBA0z2AULE3OFB
HBm0t7QmoFjKlFY1Dvgqe2IRVdR392ESeac0tin+VsF//UYIDcUMa31cBGnirfsU
UKV5sQeiPOlkz0oD6SCQmJjFQWlOB87dDbZkMGirmSym83iMjYG4gUkIAxO4+0HC
T8XC8z/5YvWgTUXPaEHsr332RWg/CmoIPkKKL4t2Xo97fKNqyMgXafIDn1PovApd
ZkX8V5GegrdMxXY9WPo0/0Ybw7zymwMe6cu/DHGtKjd7eAqyBjye2D9NDgN79qXo
qq71MsdmuVW35QRDoassLVJdQaNqJo2Ub0eTD5BrIXIDobZEsHYikInQ4Stqy01r
k8w2uOJRcsqNzRH9qWaUsBytGyfUBiFR7pnEdGTJzzy5kR+3RQRGX5Fet/9yJJEy
P+PWQnWUYnNr4SlE56D5biYlLRgvgqSoWceJKAnZ5vdsU4WQOhWZBvVYI4dllYD8
MgppZaLfp+Zf6YKoo73NaEJbMs6ECjHTtQqUGsKUAwB1nfQO1SOt9D42YhWz+WJU
w6bXsJ6FtWcsa3GwhPj7DVi/ACDfS1llwJmFm37gKoalkTWoQJdd0j7myv7u7WD9
RIl2T/zAcLL1wWt/+87O7N2Y7di4mtFoq+y4dWf3gUynh0cOe4n+yvOVHb3nKN3h
ismBDxQxVbyi1rC00aMi3Y+ac9ogkm3ggq4LCPzfndV+hdu+Sz0D4FuMbTk1At93
cFQ18cf6tknuWTR+uPYKn92/cBSi7lYOwjwI5hzCicdduKnrsv013KJfm3xEisxX
BvjzRok/kKgbLG1drK27w80e96YPIJN/xKdb06LDfSzEybH9BZt3nagquViFkGNT
bCJjDI/y/1e5Wr9CUI5ej09dPGOjh3A5amCi84CW1XE/z3dQ38y/nFODn2jpgYtY
4bCwnKM+8uViFpeaQJsUNH7lVPZ2GgVkzjve8vwlrZgstz1yh1shAbXUMBqGQwcb
q8O8MXTsxR+MXoJ5ta6rDVnQs5TwrtiQj1vjJHwvyMp6AgJHaIXJDegnVwBw6pno
pm1JtGA4r4BeLp9VRfbnaoM+ilxp31XdF1/BguKjkEr3z1C0RyJ8+xtaiV4AHtib
uy/BHXURKhAboLhAR98P4ztt9ua+BlVp2EOuRqWj4awAvSTf3uqgZi6huh9ZEUXl
1881ep6RocXGvaye3pkYRseqlrCO0YWuwvTwy+WP7d4QrvcXCGuXOcv974iv6uQV
TYZSAokTkujDK2nAkTTZuOoeV5BaxCayZDrXeXzgY4TqN/FXihBJYR5a4a6IJ4HN
X73IhDVev6TbR4FLUPxL0dNep9dYP8eADmwgjQN+5QpSNrjbxlNeyAoX40s6N0qr
uGo12EwOXNdGRGc9G1Q/N/Cwt3cKNR3tOFAt3WGvSkGkLND7y8eMqAaLaQQO4KyC
AwBm4WfAWwZ+dLgO2NpvEEXq9J4wDi5AnPZUbeIM0M01J0aFsEKtoimxvdB5ZKia
m9bCz+jt0+fikMu2eWbrKL2iSbTIJsgT31c8z0yZa6EnrpLkViv0EVv2xxD+fy+T
5JiO5XdUD0ihyIq2Jzvx+yDkERT8uLA7AdVxflD2glglF7rU5u++/aOk3U4XlYao
naXbPLqItb9ZHAdlytwnkLhX4v0YXX+hFJeqeEw1Gd5wd4NMAy6tYytAhBFNDgiE
SZcjsR6sQBgHQKhdJzHvs77zgeMnl+NHdJ6Co3qxF3mUg1O4105oYSMknu0ErKNl
IO4Gx+FynyFIHWIhKnlWPGl2RLmwkW7yZcPI1HagkiQ1u5EpUlXCIrYGo0dpJDCP
hLFxgzvMj+nMMpl7RcPgSufA5rY01nGBJ2Ynw2kK5SybLesvcqe3+yA1xorgg8Mv
u0wrR2jXA24vaYKIOl/QxDQZ9zzr3CePtYeaz08GMFepf1rk0aDrt+JBFeBCD3Za
OqVjpY1CS/ZHfIyMQ1f3XKUBPieuTn90P0zsUttzk66JbSsDXc1/GBORWXuTU2ub
nMUS4cvbrTiGV3Pg5thFZdQVA2dyvHut3DePuiLwIQdlUDiNwdvr/CthjqwY4SIe
WrXXhcG3CJhjQtG0HY4HaOc4nV5031JWSfX+8CUTMUZCKsfd3rGgNH5epm+O3eLw
/76WAJycVQI1op1JvmjO+SNUnYK7SmKCJW62fDHfPn+t7y7osJlpgGmNlyLTzL3u
hEcsZH/HVAZMyiglBVd3qu14PQhQdEDVtCdm2zvdy59UmiJBnoKOGDkgUY8We3fE
N8rAMuLeCgEFVMdSY/PZ2U9kusN5fB68IDVCiJJOoRL7umjwT2em9lu6wSzkt4GQ
m7iBRB7od6NSpXth84Sc3awZFE4Rq3k4CXDCKXKvifACYddV+MljZcQKKH39hrFx
3IEaTBEFW2QezcAyxCdYTzFvSSkb15t8+hQI1o+5VPBtn/H5n9U7zdBnbEZh9Bs+
NyDAE0rd6WdyA2APlEz3km8b6wgxD+BaFPGrnRepe2hHVrNoHaLfO/O6TjdjOqRD
IRCUFTNaIFMc3b1Khq7M0Yr1I/N+VRsBFssItrsmGuOsh6zd8b7k/UNVsblCawXV
kfHu8BXYW8biGQHRVpxV/9tS5H5aVQHBq70rMYHaeZz9iEG3IHUIpUA/x+I8Jl11
u4Tk9kiBdGVy8/okOkIKc3oAOVgSGKZaq+lhizL32mnhVeYOb7SeUbVKVpTKw0nd
LLh1/wuskj7byZUXVwcEWf8r9K5fluLwzUiDdtFqW9m3bybcSQzC/Eff9j+X5vkW
U3Fqs0QB9vr+l3vX69TmBuYqvz80xoq6d2+tm+N9PAcWRnR/yKkive4APHiueZdq
Vqv/N9J7qdStcNRpi+np1Z/yOE2itECX5Q+XY+DsKBBPfviYxAQdhmt2YEsOZfjA
Tz9Np1Y8a16eXpabK509F/n3n4QV4EkYmQZpOuAs/SLk5yotZQ1mw/99yzvX/yaH
TDsDR9IfuhYotNb91STbgkX/7DNvYcwrXApKJpPwrHsATFdIKB+4ysjxgvNBMSJt
+buQzupuxPmCSA2+z3WvIyoq5am1eDbfwER4oN7/lOgHvM/0vf206jAFEgcTVixT
5XdtIg6hdrZF+3FQa6a3QXqbjgfudyA4LDgKe3Lr1lh//YxLpHx4MBf5DJR2ve6A
ZonY2NGW4CNv0g8rJVkhwGyQGP4DpjE4tspt2+ckGIns669M/zGEeg64R5eyUmoK
JfgtwgzR10NhUJ4ucEv/0vXpFcvLCF/xpWPdrjUQC2HBp3eFaBGCb97JHHHQgC5f
8C4gPQ58/LT0F4ahsm7dJ44QuBD2EzSDAtRMLQQznHkszX0YncLJOT+Och3ADKut
JRd4Rayjt9vIhWr2a3GfTEPdAtIyLRRDo2iXnbN5L7wemHspyDL9RBEnXIkXkS5+
PrLsEJ3T6F0vDkSkICOjRQF3UT6QKwMhFimhg/PBw2z3h8y4AisY7Itk7Rd/6VFS
optlbxNd7bpGGA46QDIQJE89rVXuHIf7RIPi/VI8cjcTq4VzFPAFdDVY8X9t/h2z
mfv6txQ/PFjH4GsdhZGLcYPufFo07LUYIZgpU18YcNLWkvQlKx0rRW0HopBpNFaU
GXTT4zcIa8drmJ/yH9Ogw4TFclbBt1/o8rfl28GN4C60gjAlWRBDeyfi5fMw+xj5
e/jo5OsefmjxtFqpyaIjc+LHRLD2oimWjEy3rIgVo/SgstFMWapvPKpfE3JLiCzj
W7q7q+HC76Qh1KQrybFs7rQCMGeqGlWZDYFaOstTdlBYuwsHYwueD/3soh8SGtBc
sYvReXX9hkaLilQ/YMtHZ/eHw/V1opB1et5lA9MlpDLYQPVQjm3OkCG4hvfPtth/
v+Wieljvsf3JZ3V9VZGcqg2sxR8hPiiRIEqMj4MwqcWZrhreW36+KaraVzA78el9
buTxyMBUVnMO+/mPEYt53dbtz+iaqj7dL39kHIxwgnyGjWtT6t6uvH7wlo+H/DF2
FbcLTBrzJ00Rgcb/Rfd5GKGgfFIrSlkWuu8Yej63Otxi0XE5vYpTCkE0syLjTost
A4SFHpoRdGNkY1oo/KeXM8WwTgv8yYp1+EmkegsYOViEhoxL2A0BIbzh2scuwIAT
Y5jRKPfnb0V0UKUpa8r+USln4K2iITg8ZBlcqJQJ7f0i9p7WkoendFMr1olSksPD
WXSEb96jJLLxMwYqvJIKC88FnDPd/t/t254yw1PmwugIg+d4Egibgq4oOLtarlA7
NxShsZ7qbmVwNHYBhOfKyyg2i3QmYSZeFxnECZGKvBTUbdBOP4BdlE+PPDrY6fHX
hZcqLOUB9NIrhjM33saZFP7JWss5ew9bGFMme9wcuXLX2fWJL2cd/BMvBmswYkf0
bvoKSnbXdvGr3ZzX4JqGeMjRvFXapKYyfFle8ggawG4+RR2rokoQRy63g6u0/pBM
0UhhsQnd2sfNJRDw55iMQJJs9yecaTiFmt6TVt0fEkRlmGqmYQNIQ4ZmTwkJ11Fx
fbz/rtV//ETRpsK7bcmANfUT8uebJ+xjvNENb5xh80Em09qLA8US3ZVLqjYDw02h
QswYZCdS4ZOQDpi4sgqE2Ac6mwCZoygkpTIYhX8np5oZDu4Fsg5ppuoTdVOv4E+Y
P60Q2njWNJnBMydUopAPUN/qLC2v5oDSaYWx+bIym8kT/aZRTAMerBJ8wEhxRRTJ
j/X1VTApn/yKj746KEAzjJcSmfaF5tIfiJ0F+J6qEESLBYBV1Xf3e8b6IfX/GQSr
5PZBVIkOagYf93WQL/gBDEz1QASmEUgKs/peTQU+Z1j2gafelQNyWqnyv4pWl1Fr
5R8XHznt6lRmYbwiW7R6kfsXxXav2oB62XZILxsmE0Y+15+bRfcb0CAshj7bjuMI
LJROBKe/Ydyo+aCQ3NpHtMUZ0egErN9sWZ64bjKbfOIVk0yCnX/Ncdjjf47PoEpN
K23hASESYg8jqXQdN4b/mbUYk1tQvDPLpSMUUIvIee+hpm09ND4jkgV6UqLAXdew
ROCbDHXYfFSRn+GgijzhcrwGXu2vaHzHYqk2hJ1zdRVq6i3QBPejLsfwFZJDgObP
9/7LxqdSYVN4UV9JV6gv6sV1bospNlwhRJrI1X6CgGOb8+buOYHfM57ZgJc4VJE+
h/keuGkphd3fqOPnJGQ3pEKY5Un0o5s/0Hf35/xBtyYY6MJMcwBWj6G2OgBKT56S
r7/eKTTekbvOkPXjNm4zEdFtQ2HQLiUgu+4nZq7I3eVTcX0cEcU2zUIWx/3L0JIH
IrbW9tqJbVnuDoFGUuXLBTfJiy7H+RL8tzhS2vnuUhDzCIYanvrnpOj3LA695+Vl
IYh9Cx78MOZtsBGUkhUXffl5afBUGfmzNxOp//qd2Jd6tQ5nLHSmbfgR7kyfzLjH
bcjJbFjzsXrJqoUw38cm0BstlSE5VRb1mmKAq5hqQrC367PC/YyFKcjEs5CtXTOV
8B+cPuf33d3USnjWHYvKkwy68vqUnK4ypZ6R9JCAMRBFH+gQSbwbaKfr2luYBvIK
s7P+vn1raty3kx/FEf6SrnOt0bpD5x7KSZrynlVohwXiSjCiJcLxQYbQ/15WMhdv
oBT/5eKQJGP3HpGY6RyZZkMpr5Vgu6brR/vfQs1WbnwyuGY+jhD08MnepiJ8oX3M
shdxWenEHCCbgvO4Ltlz+KmwMgt8hzt3H1CyQUkX+EAnSDb8/lInuDeTbNvVPwEQ
Vn6xXrqjMpS+SSoZ7nrCm5C2vkp1zSUColEma5R488Kv9MZYYJ8vvOFsNmfzcZT+
fKvVVm9NPF4N1k5MHl7NxpsPdfiiwBQEYHoIMtC6rZPogyjNYMFSTXcygVK3KGZx
cPFFnVFkhsRP5XnUqzcU52dm26CDY2am5ceitjo7e8Ngw3k+4XI97To8CXkOjO9P
nJ8mn9sHX+D3xVfuKYgLpkflB0qBSab9jwG1EWyu/uAhTG9Yey179oM+F1Cn8iEh
/AbIYK4KSl3ztpijvQToRI5Zryb1WdD3QJKjCHxh98vz7jygNRQYp+UTt376ml/m
ptFaa4SLe1U5T5NuviYAuML9lIwh2iq5uivZYVDXPys4AtXSzT8O1NkzJUBePyjI
OGjqF8LSSSZIfaIzwWsNgGlhXhWVgA8plU36PYKXIyRXRidiSpggybzYjCeaU2vN
lAdsGakuzZdd4UNDW+rDYcIMWJ0oSTdgrBv56Y7knrR6puPDw168NEMDOwr5/bRL
YpnFos46hWJYtLuwODRjYT2vvyMIzYXkaf/aTCSWrjYCWMj6CMwPUFt2S/ScpbP7
vH9y5IkHzXJ/QnIKKDqmsNps8g2/5czUAej0cVor30CZu6Lr2u4yq18hlCyzq+mJ
42+4C67Je3/RW006RSfaP3tdV1I8mcKSYx1pu4EA1wVrI9xosHuLNFqg6vIdDzJL
qSSAE9KRc7ALDYQx5WUQZ4PRFQBAsgJbQixKT9cXdCIYsWlnRl884rc09BuOAfIo
D/4PqJ2HBRUGHc8f1qqmcvrao0IOanbBZxoEde3xrCmlCuQtwe6VrbHVwWSS8ujr
9GrYNTHjqciDb44PKNOL4AjjdHNH8MPV40GV45bUeXVXBxIXqj/Hrvej74WezMBA
WDOTowok892yN1iYjb4dENu5Ui5AatlI/I8Wehqhkf01T/SfqNOhf6oX4E9m0bLy
4kurzVHQFZt/DS6W1cKtwEff3PXKr9d0RTCngUzKwj0bViPtHtkudq8pd4fukK31
BDr1QpRRvNSnOfWqkauIqauKq2m4qyVVCd8qWvMYyvtjKh5fzMck17G0KLZzUNEu
LRx5ZYqT9NPC1AfPnuPIBDZdyxII6QqR97p6kw7WBJXWS1ANChG/60ndl20oyxt1
z082hCwxZUZ1KO9dfo9aVVHELlgJHIM61hbM+wjKEr8r+9XHEUAbUE+jXic8w15g
fhUSIyu2uWoke/WmJ4oG2s2Ok/7870TLNhfHJTPXoTKhyPZxhYhleNk4DdXMj+Rr
K8XRoB7XhwO8B5VCuYoRL2CG2/dHHWIeUJdAfdKLbw366sIeN2W95/yx1M/Z8DUZ
VqAyaOUnq4qWVsRVDyUr88Ls5H6noL4pqJ+L8i1Euv/LXx694DMYcy/cTT9COyOt
IoEi22XmLFMF072buWHcUHHUoDc8zTSnhNW21RuzZs996T5HoV5XqZONz7G44CTr
O0hBaq4NdC7hnVhAD8qsoABAcMXFdfECltlIIDdUfVC3y67gFHRWY9t1pnhXVri3
2imoQelePe0NIwe/J4Ct7aVQu6Es8iFPp2+p1Yb4zV8rgbUIlbofBSkF59HDLLkM
QlfVMLPP5Ex5ZMRYJo91mk1aNV8Ht7tlPEbTqPDGVpPcYw48AwRPpooVM3aiXaO+
Za6wBEWPWBj6HPRrThLGGJneQCDly+oEeoPaXz7ySJES3fN4tS9yDf2+wFvHLOWZ
WaOs94JEF8TWXWZ3iIaRsNYOd2UIEo6CUAJhC4eLsSX8Egl5USKkInRXbsS8TRmT
Z2DzEAwM8zEV10wYGFS9wEHMP6+cnlNhYiySlWgdGyazAVZgBVpsUBCDjVmH+W80
p83BgFmw2SvWxLrfOOzq35Bua8daIpG5a8PjwUTj1cIYNtR01WeiLl9hHNwoFXw6
+qw08w5bz0AVkAM/uSMJr41dyCqpQWId0bLu2OawxfXWcvXYYcKPK56qlCXye5Jm
ryFu+Q/3bO5m4OJcYC9yvCyE8aMd2v3AoHldSCIri6PFX6PC2qlTqdo3jyM/6nMv
jcYLTnonmLWU7tDvC9S0xY/nVhA3TjQdXFMkEPqQEAQs4ViKhYBHwk4uIX7UGshg
B1fhoRorXmxNY1saqzD+F8BMO/RTbpkKog5xAYL2tO2I9u/VeVo/g5QfB9FtGCrF
xS5+e4TQVVlCThutGE9qrVsGjW1QKjJUSnmmb6lyATwXl+RGRc1L5+o8dLtSxs27
lzNFcaGOaaC+B4Udc+es2AL9ncZjXVa4YDN9p7EwqNX30nyyQr6cru3mqniqRTRY
ID+PjtMlFR8hbCAh75JDgCTtbCIvG4V3liAhCE25hxSUE6beAKuF0Se9EP+djUs0
fD2Pyup8K5ekgslTavTH9mCgNLedxxjFaj0vdmQxqI0uIGq+/+AP6uwDsg+727SR
6y6xsQddkHgnl0RttBj8tBY1wk2YrkqLYymv1gdvyDYF7/f9BPTu3dhDck7R08w1
58XOnp9RdHQgAQPnHmCZnTolHl/5GCones4FXNyENLxTg8OZ+LoanPVpXBp9TFwT
NvBH9xexv0KD7HnPMmX4fF9/YQZyq12xWNCHODYxqV1cgj2ujO7mBHH7llQQYuzp
S0rwTzBjAH0BwTYOK16AXrdM9gp1IE8cZKG0Qp87oPrJX5eq+M289AGof/6d7wo/
W0oWKGIaPi7xDoRdw7VAAiC8i+TMe0izhrym224ryCTCRtfQkC1yBDI6yeuFGGko
lR9sUeszBkvZZ1XTP8MqpMpZgGXsKTjrJGC9/IbZeFs4HLdgaPYQQhd0aX8uhQHe
pAQkvRDnKo7+NmdhJEmhhLjAj47zfC9riTINIpGCtMQUqWsvT7HjRkC8lhRt2Oxw
cKUJJDjZ1Eit0lU9gEkGW09ao15F0kl9oGvImA1eq1T6D+mQnKUACqqfK6hyRnEc
yaNjPHzkpAgiGadPtAPoV27Q4HnHabr99U16DKFzXJmdm6/7ndn0tSzwtB4VSsa3
38cEVehl8mEWC0ag3DvEVVv3m/0XzFyAywboF4Z+2v1tIvxaynNFMp4HJ6lNaoRZ
DL1dsqi4RAON/b29U2oGgW+8/voEl8z3ldc8del5z7JwkoinGsawxqZykfKlIu4P
M5kXX03Cr9beEwQu6IMBCk9Aqx6uKqw1YAUzLFtGDoMhsBwq6NuR7UlYx+jvpsfP
j73TiT88izP/G1H625QUjZqdx19QkdDkZf7ReRE7Bv9cfYVg/kzW/jPWaq7yHMoc
klKzrJ+isWHUY8q1ccWgeyqwi2ltGEON/UGMLYFbDkFB39rsb6mxAWQ95rBB3m+Y
t7N3bxty1MRhA+7pc+/WjQ4aZlNdmpiSYcPh2NPaNGaWqecNHObUU93HhWeBEMFE
aQ6rd+RdEdteblY8xU2gThWmi8YuD+f/yx5ozlRCh3xOl3cY6uV9kyJeKWf0pkc9
SDx2GhDHiSJuJXEyWbWzVYFQmPpDdI7dI9AgB1HlQT9xxJyKWNcBDOUjNX6onb+N
uyMgeToPo5OLTCk6Gjur5Y4FlJH/lO49fYaSWfJ2eZM3G4vPPd3tG/J2qBaUeNTj
4gSn/2p6+DN9+CguFECY0ARgnzh5EpU3jGkl2dVbkxM9hJxrVU1rkWoVPpI+KiNl
V1YPydyVXao/X/HcrzugljEGCbMc7W+x9pCFepCh5ypDGRrfbEsqXqIxELwSYjCS
vqSOl4yqRC+4qhM9VQ+KWm4WFVr+/bYLii0CQ23kDAMHs9n5hRxRfhSR1Pdfi0Gj
H5JyNkaR9i2hBxYNWofLJgONT3c5WgE/+hVNLJ0YiXLqIyJpcQiENmPvS5GFHdf3
0sjnbI1pqiQjRr+Bok8LWqDGTc6dNKEUOgcC9hK6ynAsN/B5KrMpIrkx8zttlW0C
HNsh7c3ua7wLFndTn1ZhVnLoGsfx4bng4waX7pKJ9cEtOXY1zXFu1u8aIuLYy1t7
WOJvuxUCmdRogyhnfrjDa9Xx+jK8I4LwOT476j266zzyQ6NOtoTSvjvSr1Z6894u
5rpduJGjgo7qXwuaXLM+rlC8n9KjMdP4U3vRcInotF2r4scYlJK1rn2bk7aAuIHm
oApodAC+h/x3z2KHtYBx2aPvZlq9leQaflUalpW3H/mXzgDaGDT6qoavVckRocEg
xWWgLoU5gzOPFHxCZ4MKreOokMdjjdQw7MyzHRoO7lnOfh1znlizbx4goIDKrZhx
gjqXihr8ofnsI2g1hI3ca4csElpBUUJs/aaF915U6sU4f0GuPyolNOljYLPFqd97
5iIB8/T4Mt47hWL45hqAWdLYN4Mu9IGYDNJjcgoJhGY1adx8+L2O9OuXCztkr4HI
t2IFvVHaoUzvdtr7DH5yOxjjquTi7SGrglGDs5uYT9Hkkv68wL81mMP2fXwbgQ7E
Tczu4mmtCTGqiJ/tBs5TTtx8HOQdqYRd4cocXmTTBd4G9vhkHGrw1UWqwJvy4rYL
QDW1a4DK0B1aVhpjE4payzkxaoJ2iJ79ytUEjsdWDdvG5fLQ8odJdkVUaZiSnMa5
zuQSY0C3Uo14oJ1L/MKow+7xk+b0uwFRqX3MDOkIYPE6RK7/Qb0fAllWLPP1gYh9
Vadq1tr0xYqAsqHTzoRnFjtqIfJu/AOWnK643WlR7LRHlqCBKiCyDU55WmW+c7mT
ZtIEG3x4rexlZ4rFID4lzKdS7uSAhMOGu2b16TMZFm209YZWjDlvlHvbbAiDIzU3
+0Y/Z8AnETSYo9ff/rZstc6ECj31cuqc04yNTM0ZjFpttwc+Kl5zg3fQuIFywTVT
O2IyYp3IMbYUPM2N8aoWFuWLcm5tEAHXB+cXNUUyAFaGeeDdxMFZjgzd5YyzoiUj
f3caEXVnxMT3+BOuAg8R9KSM4jLLIxv5no7Zl9GtiuFUS/8DdZr+JVlZSet+BtPV
hYP8cg9r3W8mVMHwJu6ttWGmgdqfKIKV2eAYqU2XpYpCVVE3JSTfL+py54kl8hOe
e3xruaC4No16BIFDZEciopuX6sZvmgw2JZkw3VGHGqbkORpL3LeEtv5iqcnkVYgr
UF3aY/yQhDMFLPwXUlqmO67EgOpnFuDxmoR68W4nMK5150ETFPvcvX7uxmIJR09U
+yg2FVBq7GsBvJJIMzmri4+C0xB0qNKevJ7F5hDjdze7Tqzju/qs0yQ6jdkIf1aq
OTMlCR89Jk8OMCrdQjHV7yWu+smLnHQA7fnpMzkFXVOp9xjUUrUFamp51CMUR+z7
hdrBlppaIN3zAns5PnKJeGOmMNXfTBLttDQ5RuAJs/chedooQ2xBuRT3OTDhAe6L
/qnNHIEqIZXLZ6M2giPaP0IgoNALjEZiDCaK13fYyuBZaLz5KnDyVvuXdsDagVYW
7XmOut0dtu6ttIzrAJ8X9Y6IjJOV698rgM7qquHJItAIHUqRYgmG0CSQHApvjvsM
XR1jk72IML2IuDUZG/0WOLOOhI3xLrCg7qVmP+t7joyxBRMA89Qgj3eJzgQTt9Mf
h4duejFE7vuhPIP/Di14C/3SgGE+Tb+UaBWRXdU9HJMw9a5o7YuRNVPeyJZ0yr3H
KQXPq6eUfiiTNNYsc9vwDtZs8ZOBUThXgc3Ih3+Lrg8TvXqyMYLAQ42sWX34eM3V
W9ugaU/zXnaParVlysrx6QTPTKjhsZb95nMw/PmG8GTx/mTOKWI5gjCv5sW7wTzK
ae9e2LFKq0pxS/TVhaRaY03W1uArx8WkwY1nOkq8qQDss8UwEzGsgSCMBrh5rO7y
ZXNbobbWqa1lQUu3djSBvpVx34yP0qmEiTQJbEoTT9cbzDouzvVOK5Dr5JtGmLJX
8qwQ6jj7TXw0jKFmTMvL270GUiFv/CvKP9mQS/Gl+Me+mzMqMkkwE++FPK16DOOL
Ia55RG+ph1XMu4nsRd8cE1uZk8KdYHW892iRZMFPNwo0h6N7Xcy5uNHVYWtRRlxr
k30LEDSwfqkp6fFwfxjugKx8HER2DQtOmaTsR+tP4EaROzrOW0vR5jgiqttzEPru
StSGA/M4plIo4Xpmj9nvPV7Ff9v2IqVSjyBYzUeyjl7csm4sWGxuu9OZxJFc3sAz
hZUPj+pezWrBEmaWe9snWHCvT2nONcMgvQWD9+PIBfgsBK0hg0RHLfRghSCO3eMh
KjC9zXc9ft71Gj5bG467Al3H6jX3HqIyZiCmPc8pCzpGnQE7KzKDhCJDLKQn9bE9
znOuc0Xw+rNKWxYNHorDWXtjZ59qGlR3tR3J3YAf0qosF9nsFBouAKtYaIHERdn4
YmonCVk7VuSgKqHVT09V69JrmrzYhBKoXs2AL6JsEU8hMXK9NN2NX/GlnQUQuKzM
i2FplApUUbSf+rYC56qav6PqCYg9hTJbKtkK7o8Vh1r4UK4KpwG/dFIoP7usj5a8
NYDN4a4GxeiBoWkEf1AJWqBhBc0DCDDL3qyQWthw4b64I0hwZVFuwTGZnAjm4sta
p27w8zbxmSM7E/qwoxxtpN5nVw7Wn8l4R6NgSZ1ZjbzXxxsoTMR57vzZKLTx7s3q
CTC7PbKmtyEqkV0raMLW/PABQJ07YEk1G5fZ32YCIps62KqyRe8RHe3kwZo3aC+f
WVGNDZI9d2dVmaOQiRHDZYGxu+d3ziHpx5JyDF+SNUDFrNtCNfIxmpuQm3p8j2TI
9D+xGSOKjwt06ie/bGNhdxSQn0xU+d2DQI2SihQQNZmF/LR9W6RaWGWKKu4O9m9A
SRWq49McSBMAkEmY0/6q1rAKplRRi1A4PlmOP2/YlUTAJAp3Z8T9hrwmr8OguV2t
xJc8j8T6hH1+9BminHnL1pLhYwRFiAXCtXpdkPvEDeRpQilIG3Yp/xrfLCh/5xHh
GQ+PN8S8w3Q7Gg3dEqbCTYWFOSHpnlkKm9HCQLTKWPxBrx1Q7ZHuuBFhFzbiIJgF
G/ulfOd4kptrNi+R0eMU72LyEmH/7KfHSLlx5dOi45tPJAhw5/C2c6DpwX5pQBtA
e3wYNBslF6Whutlx08Z0E9UAcJj06OSA8JStGzbf5Mbsw8pAihqJWpAHMPf/U/80
qE7cmBUtiMA7gYLikjErQE1WaNwrK3p2+1pQ5wMpainakE+DEHWdPeK8Gsp3QBLX
+tdCcpe7xhZ9hcX88FUoaeFonTPxMM/w+pU71d5/0ni8KFj2vBKJw62jHBT6/b+/
alEXnl9u/QqnnFPAyveesHoKqlZCDaYFbB4a71sdh6Y9FAYtdaNYGBdkSvr1yvp/
VLXJ7QzvnrNs7mCf+FXahAuwkA8tXLzx0gHoIMDn7DxA16i4MwZF0GiSRotU97bE
j5v0l+Uj0Qz+vczqMfYBki3OpRtDKYXKqYLK3OQZXiBHAAEStek99lgdzDq3Z822
dTTaoD2fNVISPHlecdXTKc9wA6idy30hiHVjhz73sTwXYqpNt5LwmMiqVd9olg2U
v7ucYaeo2rEnzth584ARntT67EF4bWH3aBbi7dbOERmt+0jXPYzhBkDebuPuC1/k
YiS+GJHLarscNpWTnFfcRkAaWZuyaMemEeAU64vHY/wJCOpmY1ZdBWQZB6dAhsf9
U7CYxNm2ET9+wOrORRzRVpOfuq0z1X7YlZ2SYIfciSb1ANY6XuRs/rLZ8d9Yp8S1
49TTd4HvYHlrP5/Q2vK3gdK+5xL6sZK4zDCjTeLv02qFLmo9yo1u3+qzn8UjhkOJ
UePba0nnod0NJV/xG4hHH57Eh+bWkVGcth2gkY1ETYPxq45heKqiWubrnlly7wGi
vfCvnT7rFIzFRYua1cfZ7ao6gmj7rMaDAz4t8ancpCHLhn3BTKddlQIHXVcvcI9z
8cr30tzCSmflbk3++jW8Wvbp98YRXXwfcWkDB1Zrdcsdp7QhB2fDFDPsFJ54f0xS
6bdHzcTqBBDBE+sW10vQZSxvYwg4ARjRQs2iUmwtZb3WNd2irL07NP7UIO7QAaUC
4oWHSNbk/ZQlMJgKH6kBOYFqdGGVcIXMSapD3P2PR2J07aaqI0ZtkrKvLoJRgyee
TtATl8eLXpHF7FNf0Uh5EHc583vFB6tIFaZm8vpBKkrAmr2+6cBb1/HNIVTjxzgL
vATLLXoR0emZv3W4CFJDd7umE1qAk7YtUewnN5IjRy9Lm5tsfzyqw1M+slqFjg0I
6dN6tTs7TLfGZAVpxjNMv6UnIQ1N/+Heqi4ujomP6lkMBXS8IwL7WVOiokdvMGnB
KSTYfF6Jr1AF3VLr+SyEr6cMSSBJe8zjROkQB9Sq8w15uvPg85Qcoo8TA2h/iuoT
/HQUKF3FPy5+c4+VM/ajIEhVdpBLQP8obTaHcm1NNTzl0fqeOezKjCWzjFRMT8o8
o+eUeQL6xCrGKCDN+wRqIqVGeko0ULs9XXfVV0/2J+9GmeXvl5xrsreiaRcFz6iA
2zct7GTUyvS9j4ttFewPgmxjQqKclFRqOBZeUx75ldUb+9mqbEsFe471LBkSeDvu
DdaHCMA5AQsaT7ysILcF3B8c72f7xD8h8aVvZ925wl4qTbt2p3vyaEekXyl5yNQ+
0FCgIHwxIxzevcoRy50uLO/f6snC1sMPZIcPw89yUVjf1YxF1EXVWKs4yJdOfA4K
t8h0iPM9t6orm4ZpGECVag0CIll3JAkfjdzgqs6LBS1Pi6tBWbZfLHrmMuxOHINk
gtT3XuFuZDSULte27XMr/XEcL3qb4TahMqwdKH+YrLTXX5Bp2WEgch9Bs+Ulu2Zf
XsZRKfaF5SzngU+Ov6ZVHNw2YbUTqbs/j/cRZn+XjTIcc/6s826VoU9Jvz6Tec61
JZky6zmbURIUMsMEEH1fGG7tdWDXOKTJZRm+5Pzhy6uXpMr9xhRARN8Nmf5I9WWW
T1saO9Is7A22pDFlUH7osmajslabL8hQvRNrx5qX1ik0Tkt33+U8wy2nD8FU6PJv
NtH2dik5Qq8DhpQxPjq+Lx6asaiu5PYqmMxv/7t1x4RT/2wkDbYdZeruFAplOSQ3
hE7xn7QrsMOJMtKWuft/NUpqAoOCqjjOCYxOFPHlAC4/Zm6AsaonosEUWOZ8Fc16
5GQebZ9A7xQgGJtTaERqtHjw+6Eh5xt/QTyzwovlRkYKgOQbmg2OW2KkkqdZZGKn
569krlUpjhHP4VuYWU1Kuu0jBXbDN0/qHqQC95rt7RUtBxu12Nlbcj1ky5fWQjAC
qSEkkDT4leM/jpP2CHG7OyJnQmeniaupSN3RJhXHqoiNV0oQB9FpM2e4Zj0a0ekv
i4b4Ta0Ww+9/UQ4+A3rXIrhe3MeKCVwRsOq5s9r+JeQlunJYVNQcE/z4dNi+hbEe
83++dmxicHv5XNPxcj6aNxoIGWvrtlrXRJD+wgcF0Shmxnjhj4071lJoDHqzpre+
49LjlXtD+XnZOesYACDG8EIkK0Opx2F45etOcxEgJFMcwuSxKhnPph8rmbM6RIqj
lQIj39ZNpBY2DpNZ42uSoVyV+9u+mZnPHlXTRBNwvLHu6smMLwKclQL5vvVYdAqP
1GlAF5CiVwrm1Zx3Gr5eZurfIPCRi6q+lMsZ1n26Bty3hIsUZmR3rBnQQ8cwdW0I
LdEKtqfyzuW3cFOT8+cg2MSjS6Nfq0PCT65GQIKpibzYixboyMWpl6DWP+lN3MZG
4Sk+R9WrgD5/Ldwb23si2ZZPr8oorbw2KRDr33TIP2q4Um+AqeflNhJ77/nQ8X/q
6uYTJ/VP+gAmJ+Scv7lHEipf7/+42YrUucPmXfNqULqHrZmCgAzWg7cJulxjrHqq
o4AX9NKeHKni6HBdPlg2fcmPkv4JkmwtcyAv2VaOCGs6senwYX9dvWHEZBAsCLZ4
872GDZPnZ4z6Wr49UV9ilDi30IjGIjVQShBvbTA3kmm/cTZGiersnXRmrjy4Feog
cNFY7LUzUiIZA1g0PPza88irquIWlw7Cdy1PkWHg4fAT4dMZq1mAvSsBUcIIyGZK
XyVJT7nLNuywz6OmxJ+ZzatKVpBtQlKSQY9/e2gMD/ASw3xuFmmcu/1+fwmIBigu
Idsyo4n+ABCfDIEhvURBgLVesRVEEqF5Urz81Gq4xzKIKdRJ0m7gYE5PQ8d2AixR
EDJ8su5Qj/c8kKphtCIgScjP3dGSeKQgqmrKoBnzP/kEYTUaySprSWThuJjSP0LV
6/dGt7aQ35KsGTLeKpLNWeH3wUOjBbOAaV/vR7b2gtolphmlq2/93trxaFODfPl4
7INEjAxKo9LkmiGPBx2WXAQ0LT6LZNuC5i45UPYspS1L4eIdlKaZ4NMLAOADUDOT
JIM4x225yUpIcoii/SeP5NfSPVbmOfAdIdkH/4wZ7uSL+JLTE4ffDObT07+czfdu
g+I+i+RN91ExyoLzyLH0+mlC8jfHDaG4zv64RsCgoTTSbql75SAd0CdSKm9YZhra
ZJgRPetOidqdNF1rU5SQyeEHAjGGdAv3ryWpH4aRC3hSoYjeV8flB0OMeQ1YW/me
oqmh19nnJSDVxXbZqUs2423E7OubWLunPgQxIuQpl5C4w9/fKk/tfm/o66bZ4Vcv
PkUZjkUibZ8QbwvnS2JLCrNszxWKOLJbSVgpCQviU5ERoHxy9hxXMctAlT6urdk+
jaUgnTBZ+orLPDrDu415QWnduE4oz+rE7frRIspsLjcTrmVcBlcx1kffGu4c5B7m
iB3JnVR/YPJFXM64DAnaM2Tw+WPQe4RbDPjv8KYdoaoItMyaGe5a1ZRNv0yvX2vm
Hn1iXucDAG2rGzvR5lD6QGvKtlu+hvWhlaTKxVA3fEl55PC5fhraw2WiUCvvI0I3
G+2Az2RwiPNoU/wGa4+CC+corlXWe+IpwdEN1zUcuB13aNGOe5hcrHzew72fbJoP
7kPu+SkYADjzW0tUhXbt2o45NXjUkM8OkhIC4/ZDQ0HNIXHCu4e7pcgwT2vlgn15
OhnBOZVFVdY5rfyHev3+tr8p1q9c4z6QV4xtfeGOrHLyJadz7jsb/DqPYiepEw00
o7JwgQh4NISOaxDfh/OdzMDRFuI6dbr4PKYJ+wcZ78GVG+hHggJPy4fCJjSJdvD5
k37eebD/szuo4jA++GU1NeVr5i5AeY92vK1+xQ4SiHNNhR8FA17pS88f89r3nbM9
dxDuf5IVScECSL2wG83zND2c5FT8ll45KXGLefD7QXLtMjheaj9OJnFHP0W8NfOo
a1ni8VOPAmxqAn8nTNu+7645wQIPsg2yJNnV3GkT8wPZPos+Ur9pEb47DNv4icbr
Vo2u8MON0s1SmloZUnqYuADa1Jj4WdbbOw/meopqEVQWdJ5IRbnp0qMfs4AQjUot
XlgtQ0+rv6gB/zAZVDJ7/vTmgxe/fj3bfnxVwo01UXMfsLnf/LvI9Ze8jWqv6Csg
j8c2NuZQTlgSg5XJahfL5oGERvGbdNkzP6Nj0/E7+ulsWfX63Qw5LsmNkQUn0RXK
rFOR3NDXUEpQKXxHLu9OKKGufhUrNB03SqRVRSGBCS/jm5t0gFeQ4/tZIuH+6k70
Kuy8VthT2FEW5/ouUd6X6ytuFwmVBYYp5ffBpnBDTzsxb6gd0llG+i2WGZ6fWlVw
VetrGHMbZWj1pnwm8+IU1juCbOOTWl87yDpqSM746kVFfpLju3xagtQY5j1mNJSw
Ed6p30jbj+cpH8yUGCqUshX3A8EM2OtKU/xV+VJW0z2Dv+v2XuulMi5V+82lxTAW
EJis9Xhf9DVkKlLZemNyRiAsmjowmoO231WWtD3Ullzv6WjDrQ/GWTIWF59x3HeQ
QOTmxjq95BPJfQuTpWahvM+Scl+wpRuaK+ix8KBVdUWt84DDG4j69UeBclKHJUsy
gAxalT75BLOiyj+zTRPLnchw96M8oynaPD6RgsQWJ09eUT2V8ISrgmOHekyVLuac
aBpvTpoejCBDSRgA5hIlR6bTIF5MQ2AXldxfJ4zecdSqRNKvfnetlTm6eIO2Ctmd
tc3E42RLgIQBpEaDBiPIINhQnGYMzibsRWrxoz2RsERD260qPNWKujjQ8AiVLg27
Z632mH+sj0pSIqaGSSLNRXpjYzTN4DmR4dTAtG+eCefa7b9K7kqg8q9P94uCvEfN
jQ4ZNARH9oPeeJm94bN+UKClQezL9Ra7aap1tKx9Q/5qd9kTQeo6p6rGNsVFEwYt
5yzFdwd/JgvYHVwnwworuy0YkZ2lBKv9FGnlrVJgfr6+VFghBBcof0tLVyVwTl1d
sOUYz3bL2AXQnToAAJxVb5vvIODDxYW/WGUZMpt14+PqfEYUF5T5G32Ksg2PynDd
QpSYUpqxtQqxKhH4cD3H0e9AKX1MmV31jCL7DHk4ZIy6BqnGHAIInZcfzdZt3uTa
18J0PWrYnUlS57yac9fpEpIKsCFmRs/rZjNvkn7JE+oJhDHtuMIXy3rCwul9WHqi
i0hna7ILzjC9sRxLg8v0ODMmsD9WxCE9Ee5PUAVF9Z1XzqeyYNEcwMbx2VbEsH2P
GYbHL6Ki7iPtfPt9CThJQ8CpcIDfqKGf4Tr2I0RjhTt0nZ1hF6frD0EcfRM2IXp5
ZMah2TdqQerFKbTyyHws3dLosgvIxNi4zpc4+JmUnkfWOYMjbd677uLzNYX1XlBm
LFPwKNkanHEekiE0WkgAOqETbElHCfBoIR4SplKyKuSx1Wo+IgQo8dsDYb61qhN6
jH/Dh/ZQ2CUkn65AESvmYGq+sGRU2QhlvP5CjgIl9XwMxgrPPz5NsuQWO7HHhVwP
OiJnWr3/1vOy1PcIDZgBzE2sWUnudj2YTKfFA6j1FNnC1ud9RFAWHjKjNs+BhWyj
ULDPcB3fq4M/5VINY1sQk06mINyOOnZkHTcDI0ogrfGK9X5PZa/i0gQpH6I5Au2k
bfok1ZwLNhKXqPviTHIciJRBbxpcW83Od3HBNS9+Yd+LTfMYUFqE6e3OsuF2bchc
rb0NnK7TFkMH7jIstACdhpa4Io0TTO8nFphrAFU3FGpmGpU6JtB3NHAsbuj/wH11
+A4snLmJ10uIdcAv2gwpODIGjCeFs9xEUpMCZVoANcPCaLCL4eVW54GOH1ps7FaB
FkScxkH/VIff/HTTXCbdlQMFoZ/8q4hDFsDgtwQybRljatZhQSX/bLhgMnnd6qkl
V6FZvbPvXThYHNPS0/iTIPIZOjQtvQcbja7gyLcRDCAMEOlvybHu5GKGROKM/GKx
k3ypVxHvgVoLLakS8Kow6a1eJcR5BVPTOJc1a2AjPoRyrxPJB8ILmCBTqLuDLoAj
uNK2hQJ5DO8MJE/fTQ05k0fgrqifeGNd/TatWF+4ryoE+j6PSmHVGPuDwzr94uS5
hLy8ix757TQUN3wJ46CrMTO/aRxXaRKltMOWblGPwgGNi1xR88B+l7N8cN1lUyNn
8Cu4KNj7wembfJA6qniu0feQjjMLrmdmNoFWqsN5dXo0J/3a5ICybP6teb7ymXJf
npoaKq/dZPItWyG9So7AshYTS8opAF+Gp8uJFdwfkG5q7gkTzDLXbXGXg9+d5OBP
0v09h7ozci+wd7uVXqJ9kLzzpHHyhxqhGPrTyoreGSqi/pHvGqDPAKrQvzConznS
8grShNOrT7BUk5U8KJcEwdVPa4ELWIN6hLk1zv65Ui3i3wqOfIay+is2xcCR3+kk
sik0nfT+Nc3/a/auFL0DIVsHIiDXZoXMbrBzldDGvI3srLC0rzrsjn3qRuvNHho5
LtUAIDWIn+gEHzY7X0QfXpx7AdVkC8zdCobLTXCens4shRYqo1LEpE5E139cJ6sN
uTMOilM3IODDr7R7twCiHUvvYzG0mHWJVLVsdMBUAFjedlS6NjTEGk06J2a2vMu1
mxAljyIN/oe3SCkPAhbhP8JZtircVWvm4uiQPfs4HvsPycDKyr/xetllciImD+rg
DQli5AJQ/a+mfR5JdBr+Fj1O4rMaLyMz+ZOzJ1yFIgfFls2xFiA0QG03OJ1oLfTf
nQTp4U9wEO4+b6q0trLJ2fO2rBHYd+YZEi9c2uqeD/jZHLREdlD7j8W4jLHZWUQ6
x92Necl23nIf3lQ+RGbSC1pg57HqfpZhErVkIz+7yEfv7wtW69lbzsrH+tl4WdxD
HxPaBcblPNBrez2heKzpjgGz60N2ZD/TnB1sOe8goO4uT65Y26UubLpANgVfVhNQ
8SvmFEemfqRa5LAAz2Zd183CnCDXI7rrNu8wy3ypXW2byocubZTX399vAETl/TQk
I50fB0Nexi60OpDKVJIiTUnSccme7rbdsXnk5BqOQNfpb641Ic7K1rwGBlWgWkXo
WQIlxHaork8CqtXajIoV6fR7zvXaCG5gUPB+WpJOEPVKIvuBek6BB8Mj8ykLvh1d
SudfT6KbHZvEN1Z9L0BHx+2HMrW9wZQwMAo+qq2dJNL5wxR4N19TuCroID2SArfS
9BPOdqyXaUietyKf4OT+oH1Yryc0P6YaupnTS84yhpmlVpsoybawBzPW0yYYen/l
2taEp+gOL0BrH/RYhVd4ApvTl9E/qK3Beys3QyMThm5whXed6qqNLOzfFDIWPIh2
uyj8qVuAGB5Cs0UTEdexl2u6ErBz0JT3i/gg6drSpMqiJHXk+TnzEI6+AlLdRYSw
gRK/+f/l5U3mYpjfviMhft/R6chvMyigbeK7E2kREBQtMd9ObnEJUVGtTRike7BW
A8WOGjPuYjJMG8PCQDUtKI6NBRjr2L9ZCWIHiKisuV5hQR7IsPGskuguubHspPr4
muJUzQ4bdJxc+12zCqmFOKlxFnJOP0tvbpCcOSbJMXeK/koA7hduCSc7aoQXqJgr
GuLK37lGwKIBoLuuMBnFPupyMCavQd7BWZtt3yYSL1XxhvDkXkZ3IkExmZ/H6sQ+
cexA7dsoRCTXa6bZOPVUrlH+tSfuP0FJDK/6xB3vMz6H+GEASHUv0ZBUrnj7oAAC
Mtn5LrPoytNacdk/lwx4lx97/xWSWKNEeXovgftDs/OhxWhOP7hrW4siSxZI3RWe
/T2IbPVK5lSVCJpE+r2+hR0cE/LsKI3bA0pJi2XLJMdJQbU8FGObCwgi/81F0SOb
dORdYfc9ikS6YZYAKLnM4WX4pkifE+DgGntUJ7Z55233RS8yemDUT8rrdBtUy2yi
QbYx/lsZuhS5nrZLLHHn6A/rnhi6MYAVI1HIWbuORSl+yDotDGkui6AC1uHNpPEa
qUaQkDhR2R+oylUmQVs1vMRc5rADR5Ah6Mdo/KYsR/rXXtM9hmzL8L+2T1Ki7qjd
kfxNAXVPd+GlYOUMYvIDASDu+BkF8nHAIglEly2AyB84RtriX/vW+prZ8AFCFnzX
4WI3Yi+zCNgEAgbU2+uU4lA5s4L4ECycM0yxPCmVgBx8Mv/j2LNVI96KVui6j8xf
po3fE82RpEBn7bV8OU/LBYN2Uv+TDv1xTDO/colGyxm7YVwZ7Y1vJh8emU7nHjG3
e+eMESAvHBFnc1e3Jp+bTqRM2AddTylyCptep12T547oAde3G7vTLmbawezHk/Op
sBkrYY6BLkMMEuYhmoQ0tTh5FrX+4tJv3KRAShzMMYdBDHTkJqBmKuISiG3xJEoi
MzwKHpOAQWsLyCEnW74m/QnsrMsMfWaQY/+VySxEhE8L+YOGugvzrh9fOUZOSdCY
vHWYjLlu1X5GLzzv1A31Rglxwcjmyv4tQ/TgkgesmvzKoN4JqGRIVTHzNBaeV83I
OX8kvSqKK7qHpqGZgZ51sLT7fa+WWK8Ji5k2hUgObvTx2rlrkKYtAjIn5wZN0el0
H9scvg8fzW/xYThTgKb3Oo5eLEnyWxvIhItEzSNPjOZRq2AiE7UjNsdoqmJMW1+a
cIv5yaXZ65W3gbXUf5+0AblQ3emmVfZbt5IzeMH+YbE7bcdB8D9tfWn2M6JJlZCZ
jkgH2wOmL+X2lz+nfMH6sxGv7MyTafBC9eAldqYxxHI6gCmAIb6UJ05iTJ5x4nPa
+C2wp2gG+HuJD4voaWACbEHNtXPLUyltos4Uwg98STHd7bSj+LajE2JrbaNwxTI+
9svVlkw1AqYss/0SEN4fe+5e6vHCif3qt+0ffsFJi3/hKqOecI/PFOxI23YWR2qH
9XGHVR7vG77lUshhlQInY9YJI93uW19J2D2P1iidG4f/W7nyRUkbE9QS5vZ+d9qr
RgmHJDTWOqFSbM3F/Sbqqt9SLe/o5OWvG/skiKLgYHdd8uNj/8xQJVZQ0ge2fo/D
v1YBR+9rtGjq7MoHpDPtqBT9WQ8FZiCwawGAvowj6RZOaRQPWQNmb9udxTM7redH
l0ca55Ze2V025F/wWoNpz/4z5jVRD+2j8hdcCnVhwH3yDcyE8k/fQhYtqQO3qpd6
DOy+GtmDyDvNdBpU3Ubt274HDlQf+oo/xsi5IIKozicEhR4aOdImNHsW3OeUEiKg
WugzhsD9SQr7i2Pk4tHjYg3kptJ4hV5Q4pZWhwJuUKkL4cQX4IjSCjdnr7Ari2aJ
fF36qvHaoXv9yvJsDaLw8jJ/50jR84fM2HnuDS1vktDgthgn0MKODi/Ct6dHtTWk
hKCzR35xKMsZHCiGVrD7a0qMLOs0ESlFncjnMrxeks22BZIAXPQKkw/Q5r0j7KcG
GsOW9MWEfpa34JMzjN+IdWhuf2tnYfUd9ZhUKeogJ0rVbVaqbiA29kTOlqEPRtVP
FQGkHQy5uuEdUWbrBzrQf802E3TUf51+QE7yvJq0Xl8/kWYvkn701uyZPpX2Po3I
0yamcKXxI93M25WIvz1PFVkXl/fMktcr4/n5uITtUlK4o/kervLImrr9SOMrrygh
lI81NGIIEm5/tqRrNYLR9rNN0iLUcKSvvzlxIMjH+9t75o/nHfs2B5UWUgpg6Ia4
YTdXr19UrwBEiQbw/rGjEwa2L4Uf2ieRN3ygRbm608tEzDDtDESOlSv6oO6Tjhm7
0xlrAbFcotjll9Gai8H1masyLQHJkj9Q/qJGsqioZnlgS67ueRgst5PB6x5z1YJn
RHCps5Eojs2VAkD74qqocjoLXcjzk/m6naSBkr+FIv8e/FW71x2wnPq3ZnACNF/T
E9iqq0bHjzwjisACyNNpO6SCrMmE/LbU6T18BV6rJ+YVVC467keqij7Od8mhGS5K
JSazzKcByF2AlMirlkEaS6Dn4Ghzg1BPCJfb0r7R+IwdVXxRybWNVEQnL6B6Vd1/
g28vd7W/sXyxce3hilsbTwxHx+SWOW1kTtPCgt6pJovL/fhAFYXcoZhw5zr/3CfV
RcQIuWuyMKtii2Zt8blytu0tK7rc7W/noQLTi9eT3i50SN5tWG8dsnmOxuuO4HtR
e1dN5cg/xCgxW+rPz8vHaLXfHmn4tru6gj+BDYcKFwHvGL54CO00APP4ASEOMvig
28OcU8hKmrs6rkwkdIdHPxad7UQhugvPrVzAis888mw1/3Mn5BfRaIMRA6ukVYLm
WInJOO9uyI9SDcsrLSs3Qj/ZJ5VfbPTLGG3DGrD3ZTcYUZXBIB52aHhWaNBHv5lm
oAwr/UMq5a+1wL2WfKR/uDebzonWu8mvWoLWFm1ombvXjfwFQiWe/yVvNC7vkUh+
I0bGlk8i0i4YI1cuvax6OrRh9nVcHqw8m2ndOEOxeVtUlBsxbc3kz10agLwWV2M5
P4ewWQxdznepi6sv50uzTvt57GhM9caT1Ld0tN+lk6hzjQRdVx0L10EF9Q6yFVs1
vMcl/2FpbDUsEIj2q1tm+EhpdaHwi8T5jjrUjugLUIqmURIUznJpUKLkHwvJU6mJ
Bg7jWaiSWgyQ/XelRfsJCZqcWj+BprJg2Hpkur8KZ6ycvygvDhLTr1rCPCvRGHgU
N/1mw1iynPICF43lBhgHX7J25A0lMGGqtBQ0qLsk/4ohVtAxfc4Ml4dnbcCaspSV
gvcv4dXWW+mx5P18j+SUEOvrWbMpUTMFtwa/vPK7ZFF5e5L7QPdhRebjjNMERnXJ
eCjMrJaF+/X/UYANxPHWRAzdimyvOB4NGJgoyBswtx4FgowJw2EF+y04Ffe/sY8H
1Hs4K7QCczAQApexq9L961h6ceGNYaq+U5BrY8Vu3I4agtkZyhhRLSxAMrFurEmI
ujPXf9hSeqtc6SEXVNOdPfHMsSf/AbMq+9304Q/+6s/PApzkhhEffUKSgOrgVphA
1V9IWFYkw9TgiBRLFHuksGdDe/6Ayn5NQ/fqy5/AcESPPwXIXJT+/TGq/0BJjSYV
lc+7TQ82JdBMS7sL3Fooo1+OElujqDiGCU5dQcfsIscQhdUz6Lg6+HQMLXg6NMJA
9SE7czZ42xh4jmaebleLjACPwQiOJeUT5ho0pe2rjTKRrCxCteCQB/DHPOcT3h0b
GPWEb/4GTYOT0zDbG8yF/YQwX1/yoCFMAHvE16GcoYXMJTSZ0KlwGWoY+fdNj7QD
ORXNt7yIxEGWKSADIPqu5VDb1PNLIgl7vzhZuotGe0RIxDaJkBETFxTosaPUMPZg
krmGtzL9VcYatqh9iGl9mz9wPbD1ovbDX6S+ZzkSa4BCTRsL71BR8H3dj8dCW1vI
FSsGccP+v7T1nU2DRoNjKdnyw4LdTxBtwwu9PiLQWx0QFQyNH3rydOdqu5g9k1RH
YR1DX6sxlXXkv4JS5+IBk0jrXVxa3cVHTVBx4WX46Hu0/F7z85o+SX3mvG2q3Z2f
PG9m6R2gy/4M1CJywCOLZLuLaL/9CeKwAcUsah7Hfzft5dDDlSWy1b7pDDfeOPsF
3uG4kWSpqIiRlvx4kI89xIuOqYtpduuvh4T5yIcOybvvi+fVCLVCSptsMS+EtBUY
+XJPBCTAKpLHMIjtCCczP/2nxMBjZrJJ/eo3hLqmsoXnOCA2cAZfKGWP2e530Bg+
dA2oC3cb/3iqgJEdYCKzp81CaYqggs/Ur2teiRvDXsxW/K7KttWdrNEYFDHtXhUo
jbb4Un99uVpNdUGiiwUA4d6E2bgBGjcruh1sUJ83JLASRr9LNeQ2d3nmBTJ+ll0r
+zghMmCuePk7AlWtmHJzkUmrw4IzPgdhsbDrokP9cUoKAuEz1uglxKhdSbV7LbP8
WYeDOtjrMn33OrEYHZNJwIOKyHmsa6MwnOw7nGM/Wy2hhJ8KVllt7Lw+VTEEnkh0
xuy3dHjz4OsfbRCjtuQXp4I/fSRlSTlSFzbCcZNLQD1kHgBA7aiWXtmktf9dGag/
ImOuIOSxr6Q7OZUDGMxG1+Yluf2I2V+cpd/Pi+BnTjlj4TqmGIdlAwoqQkFAbMCK
zbgpbOPtB162RNoWyaxqCml8AhcxuFNypycR68U1NsUSzV/YkYIgd/dbOS7rDky5
yDMvWNTwYZng/QdTcDsSAe5p0aG8rQkXoX9feTSLHHIAkMl+jRv3Mxbw0nY4dyKz
8f3smPdpjqLKLD9w5+t2lR/I2ekwRzOoFiKlRbtFG+v4Wmcz9UtsDazFjr8dhNrB
p6eW4sch7UkGSbsDvQXSjHi/3V3JAQVh7pXXCJDg6QTFzuDiz3/4ewTMQoIkAu77
ZYt592EApkHlL8XKMZNhcZ3xCXRt3RRqBokvMULaGsPdOqg+kTtfFW1kn4NKmibi
pI6PgvglKWGPwAy3OaKDcXqEs8izy4whmo29SjwFhkwSxZh8hGJA18pV7hQb9+qw
rSKJeam2VIBzWStx9URHleqP9XU1ZtUI/IYZMrOeb2oxFGa+4AQJWKBFg49MFlh6
NxT1TJSjbAhhIf+NuwpU4HMpyyA0OZ7/lyLZcPT/I+NVyKlbzcKV9LeE/8QVfJnD
wod0IEKwe5IFOEPkOiyAE8B4673md1olu/GJLLT2xKXMu+XtS+1LFOjUpGUAFdMg
i3NIA791qFYaCXUk7+yJzqituITqkRazsbitBwpjTyhvJtAHvnhqeaxvn3nBXBa7
Uez7PE2iD0CmYbnMfnk3sNJgCbi5CcExqmqytinjirbklflEbV+BgW84XIP7lv/3
iqFJtj/edHRHErpv3ZjuE9+PgjYYt08l3IU7ZjyxET+7zN2ip/rcmURC3jzAQSuB
8aJp4T0MneHCa5W6z2sVOJFj0gQHH60sJlH4ryTKrb5dNyGBFE77xbgHs8Say5Ti
Q6e/J8XOSoJ0p2UsjsRcxxmN/kSnhSlib8mztqLdgpOIQdbLXq2+01dn5pD6aScj
VkcKQ+zzyL86pJRhyckMR0TfhIZYVh5ToRZ3CA8DCz7/+HrUEOy74WHAUe7wMp87
1unYd6228XprbIayvvJq1zKWtqBwpeoqns3KmxCuUprmxDIeTQq2K8bVV15fjmL7
41Ai6OQ1QztfCcVmOvpGYhe4dwpkc9EEQ0HQWw2fNmTREUKmwE2UlCCcvPvJVXew
iYu3GDWKTk/9g4KWAIS9FjOuLiwuSazDtLQtgoCcZKqS4/2HTHLcj+AdxlIEC5Lg
5OdJbW6NOzWxXzH2NNjB2Iq7ur59emLyVdl1gdfwVIpiHCSKPWtqhiUM3SwzWgNH
/pmakB8bcHvw8cdSQE0Egr2ZKaoUbHFb6Pqyx9doX+iGoF1cg/qCqh831IlmD7EX
PJX8vkr2+8GKnDNDh72ORLQR2Put/aXE4nFXKcqJOoK5g0QR4V/L998fxA3fSlsv
oLBs/lI2RCg6gU3ceVujwMdnUM8dIDYn78Yw7t5twXElbMoKYdeyajkU36gT7lhx
FXZI3vTdJ5l/XwS4daSCy1NTELGZL2WeouHKsCEoFfw6jCeDmCa0/MgD2BXw/UXn
LxQ+YacqwfDuoPvSWF8H1NKkpdMneBgd7VWem4h2wJxS/TLBIdYu4obXe8XVpfai
fX7hNXjxhJaIORqiyhKyzp230qYa/vxSKLeSeXWW4lyy5c1S6mNkdsTD8aUN5F+D
gX5F8wO85j0687fMdmTU9/LvhYhVKVI8TE6R1BlRG7XSh3SWv1hASCT6evdaVzj/
sgId/OjbPWbwgJ7RV4ObtV124vWK+vXIBrNvhuiaGhRuvrmp3LOUKrK4pfuER4B5
/RP+oplRtP+oyGs0EvTE4Wdqf0JJBakLoIUoHvWc6tNyMmBK+cRhmygLKx8cO5fy
COlYN2d+zUMH2cMVBgMG+njmX8j6W12JDvFqV0EIDqVqaQS8GpKrzmsX/GRuEvR6
f6S5vVLwmbDDTkg2+K8OFYh5CVMvXZtba7lZITSr3FigFbjS1rhFWpyAtk+JOsml
dWvq2r5UuUY3Q+S6y373dOR7ythSWg3ly+K9BRZEUjWyk8qBIHsp3ckVvsQq+0SW
S/ynCnwrpIx6U0taLon4/cbGP2Y2Swe5IDf9kUF2tvpBumIzRfg5nLH82/qWW1w5
VHhWRLWQrUCd9HMhJ3viPuAB932KmfBp4Q4R27DwRHKY4x0IgJjJzSPmqEdLl2uU
L5fhIb3spS/jlMltiaif7oUM9kxqkTSb/p1sjtMzU6MYmXwhD2Vdmlw5yZtPsta7
WInSWEqYJS+YxFFgA+1PViX5ZOLWFV6pt6s62Ob0HBP8T9hJ7b8fJwR0bmVGd3hx
HFIXHPwrjJly5XFW2fFR9aPIqt6rdNxI4mthmZvwfHyH84XhSYoUtL7Zzwxn75oF
PPdzLTiWszAxczbKlW5NrkWPxLlcxFJ/XjOKad56D7wNojjOCPppHFcchTiA57Ek
5VX0ZreLOg9I4lhO/tXwjh5qWvfYRGzPkJgb/jEzncQoK4zR0if+yE1dA6EzGF0/
Ot3wIsAJmGJklKbSP09TLQA1XV1FPlOPGZW53el24Dt6gqhmgmY/q3q+eRi4hm6n
hHI5fNYCzHxdAmq/veovRD9FZq11vszGTn+V5jUz9yedFxlTEei59oY78zqvYtm0
SxrXYbjiUg0z9jVxTJ+21A4+7JkpTopW7TOyPTuDKP03pko9zK+2+9j9UMrv5SMD
mFs8hxBEH3heTiqHAkGV2iIetoV6TPS8DSrzpG0YZuVW/39xxS1HGTJcME2rUFmR
M6DJAfwKaAMEa+7uiOmJmwu+cpmdjlsSDiWq6zqQ4cnHi6Uc03cFyAFLoGNQIlfE
oA7DMHUfTKBnvEdNJuqrvbVgKvF9/y36lNqTn26mD2K7Hx2252+CnErKRI9NTSwT
2ej42RAfZgCEmxtpagyAnHB1ivzV3K1G8KrdF+H8EUdKHfnV5o4FH//Te1RAna47
0zaeLbdnpPjZGcrJ+hP1fo6zmmGgnzbIaAPVqwybWqYOGJeiMVPQ0OkBzUZ5wh4m
dOBEj4by+nlJ4UABztkGisSAdEVTyF1R4V/FF6HY0Zv65m13eZE4kbNtEXgkUeBu
Txn3ApHwkM7a9qzfw8/NJhCvurVHOc2Mbm0gQB9SM7rxpeDvXaXmilqN+8yz6hg0
xHNE3sg4yIRCIrfwviIYwYrbCxR4kTtvOS1SaY4i09/oOVyM16/vPjSNHednkCmd
HXeCpnUgJUFF1tZtpxNd3ZkGn+0OrM3NeFuSZLFMdW2nnk5RJeXveoX8CQ+0LfSw
Lj8lABEgyCaiOKAUcGu0dLt6D6iZ1peRgnz+xhkq94QGiQ5SVCG5we3fxZ84evcV
F+U4sfS4/qiZJlXwagJ/DqSZBkhXo+Ac2UY6A5VcrD5EuSM2I/BK/jsyaPNWZkB/
7xj7PVOd7NuuQDiRFc4FbMKuDeRW8plJpoYybsTkcBbGsoXcKrjs5x5nfNeOOAk7
0SesCmzCCYSmUUKLGpS7Avn6tjyGYvVIyfZot76+IzbV+WZbLlPesaJl3eXQBQXy
hG2fAF44zNEJAxuLBenIJf7+7zvUshb3U9gU0a7kx5Uc3OTa2l0kD5h8iUtjMFPD
jKHrGxkHIZrORT1A1xpGRVzM7MSdlBxFxbINjscS5bSkKX/YnLAmDn4RcGExnaDx
7HFfBcxOqDOjNElpFqzB+fc+48ut+8EMcachfFFAHyISKsQxlaEgfpqRjnq2CEbU
v8qwI6WlMgJbZfGDugybeMn5dMdcRkgs8C49E1nwklyzGkxhe2lrNbAc3GRaZubD
Gm0B9M3DYnjl32Bi22RVwvJAp7RVO8svHVqZlk/iRyJES4A5qmUxO+Gbu3eCt1ia
IQawwX+fb4kIlmkc2cGGs54D8usecXqBTLHj1OkPUP/gVg8F0aQihiuMqe0agdf1
3lQUuOMcUrgF6Zyw0HdV/0hLRTtWtEH1+LZQCcL+tTUdSJY/bz44/yCfrZpeVCxI
/F9k6Acxxs9SwtLzM+rcaKsD29HrhZqiodKJcCoqerup5jahgXoR1A9Q4ZPu0TJG
uv9OGsuHm4qjY/oz+ylrf2uG/7BQe0aQcD7WwoaiGIrexv7ggmgckGqe3uHvsAmh
swzq/nYobKLAKw0VQ8cZSzsCYZeprPqCdP+PlqBEaa21qGg/xg7brUeGNZruO1JS
v+jmpHy6Wz1239FBDd7QFDxt3cjoG6Nzfce2vs5emxq8Z1LvyRW2x6EHSAZWmIYx
OLmsjZU2JPSZgRHKr2kE3tLEK7bOCtgXHdUPYAoDNt/BXOH3D0ENxh4cTTUqdNeF
SH5h/xGarlpxCP0EpUoW1TIhNyIewTvUBmEWM2o5uGF1yX1HVIuoXHEx6nIrkRqf
S51WBwVUT3toDiUxAu7U6rZrFoO6Z04XsfnPFl9l9nLZbIL9syZ7a5pXRpKx/CJs
KF/7Tzw3j1tb2kPH506St054VnceQE9aY7tMy5ul5RHv3IBxak4AvxUkceMRZ7Ki
6rbsHnI7W9X7cHyiKHG1wyUA+rSF5AbEEz8KQvnqDlJDkO8Xc4exJhytrG7hzAQR
Qcw/b4TvJIwuc3125nlKZ/kFOxjyD6i8dvtpVN4gJPlkColv5nYX154JiQDKvWhT
do+q4XpGAotlBu7EIBtDWicWmdzOVtIu4Txr8I7G700CWJQkvZCuJ4UclNzBX7as
BtvTCHEKZLy2nwkPFKdA/UGapTTFqq+cyZZXs2KyWC9ZLX1KavGMoRMkrvIcJxOq
1N1bEz8Qni6jk0rg82cSqf2+5dJ/ko1NxTxolIxCKE2V+/EcLLdK3DTgzHELAEuH
flJFbnL03Ic1jf47+MZPJWpiW1j0amn735iFUHb4Oum4+wwu5RtGanTdadN9S7m2
vn22T5QK0FSeTnq5ubax9y5/9x9JTgbRyjXcZcr1bUUXxD0P67n2zKzPir0/marN
XZf7v11h0iIVySkhYp7ffjLY4nZ54NNvTDpgkc4ROTDUpswduti+t6pjpkmH+HhO
ejkhgJUCVSUw2uwQ4QnrCJwsLHUqzmcpq5Ac2KWaut+6HBUfjSf1srlln+KnmFvu
ZG88sDFRI5eDVweOxuUWNQ587yR5EhCXxBvH93VN4nLUdIyF/sdQ02jFvxAspMgO
G0GJfIHBqZ//D7qLg/ZRsKYJ6S53YVtbbn9FKD9gU1pklNdafQ4/dz6knxAsxWUq
112FHL092aoXG2zvolGUClhebcVhicQvhLjrkRWAcFcw9AFJGvdOEhqgVqei9aeV
uj+ex9N0LP1C7L65YuXdj2DvaSFefuiKjc4GBrS3X466BCx+9VOyvOUsAaXEAigI
MZhzzgl954PK+rP+gjmlktF3ArKa1FmPg2U8an6B5OECxvs9VQWyKxYfCqkEbeAo
2xgvuJXdArWAYpTrsHzeMKdSllsnepTDXL7XzuTqKYBlulTNIkx6aDSkWML+5Ijj
Q/hKUTyCz65lRffphqsi/K9TGZS5W0q9a7MRVDxdcSdqWBtyvqvbaDACkLiD6lX6
rfdc5yE7+qxfrlUPeLVDTlxKkBV2Q0aZJwIDJQIO3cuw++Z6aMgrhawh2zOKjaCk
65Yklhux/oFWDpIw5HFMKtMPdxf/DkM3YfeTZukxygyMQ+Edoo0Ot8SAMBR4QzHx
GvwhQb2bdznVT2t4dQKr8z45+awSq6XAabAnHQIX8O1AGZ+WJLACnRNSvLd+pTkg
y/UGYNjV7CxSSFce790UjRlncAstYxDEEZUbXr+D+5WwBFfgo7Imnz9MAS/JNs++
NKQ7VqtPNhyM9NEyCeD8NqPdWioG6qO9TDX7Yx8eaOCTwx31+5esvTxVWLz6w9jk
+gcJ0OMLwbJwWHCUdrMNy7Tk4Wb8VMh2LHfdhnM6P8ofAqQJ5/BGatFKl1pVYd6k
ZJ2Jkd/dNs+lZPbFgMgDMdQbZmx5K1gzrj4WNxbmVkgjaFzwKRQTyq0CSXVBR1iW
KkaS7ZyGPDq3n6VdXK2b35LsAM1FPVoe7WG8Io/YmeUgJFTwK9f+cHqBnPXaRD4I
rd+FzqAHbwZkHUozf9MveM3VUYFL+s+8wOjBHfJGhydqq/E35GAyY/el/F1o2GhL
A51VySaAJfLU+4r/blfoBWjqEgHd2OZwCGBlK+Zuxx91ujTS2bez0Zv5jKCXmPXe
OE/tr5fmytsBRNVe9Nblh16CrmkGXI5dsMlEXAzivN+tyP9OY6xnvk3DSn6IUfLA
+OW4KnJvbDlDz/T0sRBmhaNQ+9FUClj6cxSO2FElIE41vEaNl8iZ/Ax6wT7+kSpE
TXCfUA9hHsSulc5Y+VunpkigTgSwTRsZ3kop5PWM+4n2J+6ruoUYMmTQyaDavOab
Q/fLC4YRiMuO6KTlTbCKOiYXLLvbZAATNDQkq996v86OS7GzEUukHNa+1S7Qi9zk
c4nYAa70oz4iK9ZDAlW5d0BH7NVEwXw2S8MEjfsDZvI44W6ZqoRnaNBZn2goaXy/
OhrSvm7TpHqMiAmK6RWqDR8PTMbT7MlT8jjPTNOquHoUXTkJJ/6G305H/hNbstWM
cqqqkbXo8Q/6AH8g1Hi2/GaQOLUM/vpk/ApZgWW+r+BP9I4jNT6t5yCgFAoRVt4G
2A7Vogc9fcKH0SUL0ur9AdKVDQuVk77e4E5yx48oDd1rg8rsOk4Lcqe77sybTJy5
2e5WjEa7EYabWvfM+0CDvR8xu8b1C0sKwZdt/Mzu8qJquisRUtGeBLUgWHL0HcrA
ppEL8zG0ljudDrhGWr1ooKC4pU0z90XVarKAh+Uka7m0eCuPWrH5FFzRyNV+r2zn
wAJIT1atYXEoOrQLGywdQNXlLOxTzG2tb3ADqTfEXlP4YtB6d8gR5Ut3vN/WvAns
BkAbT8g2u3ZXrOcfjdSub7m3l1QDC9lUYxsNDW97s2pHl3DfYjOZjfil4IVsZ38R
si/mv59lyeh4WltUQIsTGA1uEt7PHmXnkeRLLoIvZmXo0xC6qaTQk0YC7e9+168c
ucnrilkFr2/yEZgz4rk2/t5SQolSW/dhxZ581bD/D4QAU7fafMWA6HwdGpYoK8eJ
BpB/uNO06AdddecV1wOHoxVFxBRH8S3PwZlUyRAE7q3WTylJ9yp3tlYn/coD5u9y
oMqjfx4zMmRiyuP2HFTklyVoHskZyi0X7UBlO/nqRzEixhvse0CV9OiaVsDFXICb
kciPok9o5AS/MgcooNDcdxJ3hxB4UA06yMYCkU+LvpoiVG3xM/QV0K1jweK3xJw8
pv3cAgqn7GqOrAs+FtUrc3m7pPyRgEhj0gNPvLQ52H5oGlkMAl/iTnQ7t+z4wvaE
B/Lje8TJWdZRTuNmajVUHnMLZ71fIiBAqKrGQFiN1gV5gf48hPMNqpuT6LVXzT8H
45IslCCMmWVMw5Nv3h0+tfpEQrTJkysueyv+yw22PGeQeg7NQeC913mCklAREq9N
J0jFCQrBM14PAJx/AQqON/VmcF4j66f9LgS7omxwAowWMCo9KRqyNNSqvtb5Wyo3
D/8tA/e4NBfxok25Uv2O0/glTyfTug2sUW5+GkNGj6XehUI7pR8N1q00Mfa6t7Jl
TsjrdFpBwZlvu1XI2uC7F2CMIINQzpo0fvKukvIxAouNym+RtAlDAgGYhGpbd+y0
Tai2DcX6EJONsE9IrChIcM2a1lb5lviZ/YEGC7OfnFS8VRnMJ5UZkeljecixLLfL
bSwAKPh1zRvN3OR32EV/r6AHAmbd50NsRcQO8+50QSuHK5zxzOqO17ljTVZshmca
6horpS+YILK48T3Dmw7yOdYO+39tTuAbJYN6UEM82J68HRIRrhw8TxrhNowmJcbR
O4bkC/NGA73uhrop4UmwNoYxrz/Rbk0R07q+Y+E/vA7Mkwqgm2QvZPUsnI1auspS
I4l9rqMQuZii75po/gnyALYDuwis/PhqWjKFdOcviGe0Tqbr/K4s83XA6TnqIJ4X
Ll7FJqWn4kvSEjJtIuB5BiM091r20rECiJ0sfTfphFLHNnJxmGS5pUQ+N585i9mk
vHz2s5aTbe24n3MdkaDqt4bVHUz5650K+wRYopE/dgrv1yLP8BCRzs9UV0N1oPAB
EoVvWMGH3+LLoaPxvMYJdf1Pj4JCTSr9wW4TBAz9YAFU4Qse1MySNq5s/OeIsgSF
LIExMxEhFYXPe/RZLBWQaR0QN6hc8GFDdBwqsRWx2bVTvSVPTmF2NMT7V/Nlcyuq
CQH6E2W53OGbaWhaqgKMSkOmehxMKnk9N9M3MBFYXuhIW2uhSVfUDWeWOQViL/JZ
3YcKebjkLeAmwerBQ6arqoLK/oUOOzoLkG+NCcHq0blAs0/r1HDF2yO/Jg82r7YI
FHffARu6zNuxFtRM0Y1GXeukW1IhQ/QUNjJskfttk/7GAtekRYeaJdHdzCqA/cO+
vN1P83zdZGpgDgBoDx5Kitkxn5tepAoV7N/g3NOJSyNWxg3uWE4loaA/OGp4hPA/
RiBz3SGq1HZENvOdNcfBPpSGgWgRVCCo4H6NUWZnAUzf3X2nX7qnicdY1bU2pZnf
rYFfYOCwYhLGSk8DQoWeyYUhPfhyp9Z+pPRVm2KD0qSaCufupQPExZu8fMeJeuSY
IQlmbxgTEPtByUxLF32wGlEe95gMWZkJxLQemqZJ3FKVul6kAZgK/aXpNvIeicxy
r9M9XyZCUHUlZVbATYTpuRUupu1F5ammARao6vYkPsTGNw1nShOs1MOwlGUy/aBK
cQ+FN7+sS+ylqh3AS6R5dxE1Dk3Wo6kk3A8YUAfZz8puBpKbDJ+JNBoGKCeHl5/U
6cF5SlMRlX1O2fevQdjvTlzI8FLI3BCrXJAZ637csozDPzKrRsAuwFAc1mGChIng
pp14UTSQFpWVU+MxadoU11uv7LihQRPCce70zwXqdDHbY112rvHnUkXdSppv1e1m
+F85eUD5GJOJHD7/QHDmyZWiu95mtLyfM2d8jiWjVfG9vUj/LJwl+GcmVYvE/ZL+
Z79hlDAUthhQlozqXO3dTG47XrJeUJjsbIGXSN0Jky9LbOMVySwgrHnsw6JY+x+6
Ec7IgsYf7gK6AVcrNKOUKnvM5XMLkFN91C1wNbzp+DLiyy50LOFAuSk7JXSUErwS
t5WdUjo947i7s0ED02lzFBdtiBVB9D3YOZmCGr41RSH1Xwf3xI3LKFzgf6SgoNwI
zAikFoWfGAvOp/MIoHMxVhvRrMM5d/PlwOdyalmC3xYmJhh5nBkfReqDLWPmpd3D
ipsk9OCqEcGUFf4k730uCHaOnxSsYMbD5tIZKOspR3k+iS59DfNoHHkCat5tvexV
PREg7+7No/5MbaI6qgi56qrLcOOLxNYS5ku5EvdEMYzEtKs1i/vSI4Zg4HZNckRM
fhcAyINwBH4ADfjtIH7oN0SGE6yX/0kbm8hPVOFtboUxcXtVxsJ7PbWoxVbHuk/o
tg3xNe9etW6Wx8hwFLtStS0GiudFcSHKUaXZLG5XdTT14zikwxnbT1tvSeMhDT1V
jTIDBrD/mGsl8AhRYRUYT6UX21HHxu6qXaACTdwpbIMbeadDvxOMfM5gOyCY4uvj
FbvoH6GWvlPIVzRW2927U6U6jklOASEC0epVVzyUKjqKAY+b6OS6z6/4Ej874QTT
krWRpgL+y77HHDZsiUvveAkBFWCdDQFuok+eyrTnLqLb0+x/rVbBa1Cyz8kWx1y1
WuA3LjmQjj49jsOb1sBvT1NBabiPLDx+gqXCiqhbZnyXMMwcNkCytkymz1gUMVSE
zlt+kHrQD56teje2fxBVHxOqaQsCdAVe60VH7MgbYaxF2NQ2NVhg6A6u31e0721K
w0a7mmme8C8GNhQ03COxmdynoTDDDXCjm6Go5kpg2qHilw6Ev5sfYZE5N+JTO0Ln
Vs8Pl/6ZPygI4xrUIxPK/0mTui/gd0xBnzz+Lsmqs7FoFYcewIG/WAucwsxZ8tG1
e8pMv3fsTjXTiDtq7Yq5YTD4vOXbz2lZWCXZ+lBr2v+5XzO3Bf2hyjFRPTE1P1TV
OmVmS1G0zMgkucZghOFhgcZEThmXOeSRuoMyLWyEC5CQ9Nd6Y4LTUxC8gGWZJ2J9
YBy6oas9ELOAG+S8D30lNEFBZjYK2dC3wgBr3EpApm++gqkEcZRCXqoACjC0hLhl
z6c5aD+Y7uKe/1thhkqynhw3C9tI5vwf0PaOdNcYHhGeEERpKhs9MFVnLmSr3qlC
ZmNlVQB8mD0il8P6G5aUq4H5eJh1HW1udzHV1Q/Hz+GQHpuNuD3R2/aXft0PQsrI
j1NpOYmJ4W4MBteh8duoEfjRM9bGxEOhrHKgzx5YgfRVqB5DZ8gh3z0EqPB+Rndi
L8dIy3EC2fdJoJrZwPY8pKoKVvmwdU1Y5uuzRSkngPf0vcbLE/IEruxb2oUHbX1l
9EluMrK8rEqy/Ajv1O7+PXPk1Y/RnXgaVjhBck0Dz3H2iGpfaoSP8vyidDSt3uTF
Feowj02kNU+pKUIVFf4+a/1qhClxP0OlRt8aeQeSkxaKB6KOuOYOoGngDygENtG4
Spg2hbcB1vS+AxJL1QWYGegCZ1GHRUpez3MUABg3+rCt1UFTmRE/UaYW89aKLSh3
NhLIoiP4BYgrIg02TxmuWPpASbzLZcKNYbARGsoQBoqnCnVASWI5wS+f4B9WhW+z
x0zeqDn7lJJKsX7SsuqlxCyXVtsSz8TtZXXn5oV+qKpUn1eBbHAPMokQ43FEIlAu
EuGgD+CyRT/4WgiE+UcRwpdxFDPzUhdJsHXjP+s394lsGVQ0g8knbVNI5lmdG15t
8a5zEKKuyViULM+tegXkPSgAhQkNYF0iS9WhMh087HANt7qQQXbK6RiEGdkZ6Y+D
RyqmLB22yIIS2sBSsi6G31By4IgmZgnOSSo4+camH2ExvDA40r6e4kB78uRbZAuR
UAay4wsTEKSRZEvdxbMVvTe1HdNuOUCk6p25cy1eejjCucSnb5pZAija2WXa1nlp
zhKtr2Fk4etGEzTfAHS7S204UcKqXvJA54vbFZC58K19CgpG9DIKjXV+fpIH6YJT
+J/evu95dX+ggq7biBVRyQX0M0YhBEM5ChOvDbRE8DEb48VgFHdTqh+HDJ6PPQPo
l/M8YHz5t2fwnVLt1bfJPWYA2XhlPkF4pSoocscKXGW8QQ6/b/mqTjpc2jrikRwQ
jf4ap389/F7Gdtisde0LiJnJesNqFXjGDzfRODKPoFL6aPD+1JEFOMbyhPv5wvWA
cs6DdJEnEURm51gMXKFw7RmetXqWwqQA7O0gMIPGf/m+Ez4fRUrGr0r/GK9H0sXR
m82wypxXgIu92AshKfYJP9GzeZQ75FTHmMz59GdjCJTqJulIHaUsdY6WgVlTRx5v
xN5FfFj+0KS+bsCQ2F0DKTIFzirJMtRWkWqF3XZEp+7CAWajcHGSbFfRJqkAx39n
m2oiMYB8P7iBPhPp2Yi80/O1r7dwqRkU3Sw7pYBWSNgM9sC56hVSISQkuC4/vMjJ
nK5zkvze7HZXRc6SGG68+VWqOLFnMpxVXQSz/W6QWUk6p3xAPoWPucIlACPKJQL5
sPRzLVL8TtoQqvqZaJ8ZO3bsYZd6wHvIGFkhcPunD4w1aZROw1U+Jw5omTI4IJTd
GTUFCrzJYbc9OY7VgAPszbqNFprJcnGY3FCuT4FSI/lCOKPcD+oa7BkNSvG2pdda
wVGbF/3L1wchNouU25qfelHUcNVmiAKH66+bRLsFPumW6wV3VNKLmc/lZpvB9IcB
CqfmdpR5It/qSSs34M562T6dT9LQRUlvGlcgC4I8AcWjEQ+Od/iNd27ioa13O9v1
9y2KND4lnHzHGRFfENMMTRszURVx+5Wz8FYPeqLsbZ863Lv72oiutkV9DR7G8sr3
Qu/Cv2e9+ZrYg2/C4AQDiYpY4Zkm+uI2GYAf4uU2Lfj1jyKxNoUZFQSdPK8yK/n9
fwOL8CC/yUSQpt00Kxm02jztNf3XuIB/M6yZQ//8RDRKHU3SXVB63kGzJO7H4YEF
kES1QSDQRdRWOJcduuHv0y4E0Mi6vN1dkjBYRAwsegXFa3PmnRJHEuP3Qx6LLhMo
1sfaEKlp2wJU1t2m158rtOnMRVbMjM1fhf/QbrG6dzs2YLOvzwbdxEQh/hvGlvrX
UnDVo97wrPlIjMbVk3S1Zbg/VCaP9QceYzggCnwlHQXAUN1hrJtHOZF8E5/eQRUe
ulTPW10lI3XFRcN2my4ORCfYQXDIb1B76HqCytOeuu9L+9NcgWuVuiY6h+7cDbGo
j2Mp6VQwfupSk7dSQmfzbXvTEdSJixB4jKD5HgMQ4nZAwomXa3SAd4XVWJFatnC/
sFxkRRDkPbzP4qtqATIhZaKmz2ESF4ykD79Vt2ym/nUlA35TGtdG2pspl4Cy+XIe
YstlMEKqoo+ZiltsvVwe5HGS/gDeoZ7VC1fGrPXn/6YjNUN5Lc0i4VPK/4krmsrt
1xS02lZ4CIsnmfJnkowvn1G8gD6QYoncZAlAS50c2gWLx7nw0u9jrNsp52NRR+Va
OpHbvhOf3Uu08GUzGBwqFchUZ2sDIhjuz+JJYe4w1QGxRMMcOUp0QO6MgyVA/U39
IWxYoNPUdewxe9a5/CzSB/TlBCqrApcujxqdmV8k5qfPTRnQbMlT5ehKOT3SF533
OHyswuYjdnVf9nPyEfDT8zS7zTe0mXa9rYOdQ/5OaCort6CIW+X2nJyYRRUCzjEx
YohD/dQYOydvjKUBBa+RdW1VT+G2WBxs6g62VWErWwVUljaCHHUo+a1v7KX+uTNm
6x+5nrkPBEnIe5G039fISelrUGSHyUEIDDVWNJqZ9pjALQ0SifT9hXHRKGLSg/+I
b0lmJfHBav8ORji2GXso35lVOs4xr2pmyo/vLkrVtE7fLoOd3lvnl+W9VC5GWxEH
vbpYP6xxu7wPL1ZLSgWmep5uCzPVph5WF/mDmZ1bpm9PlEUkQCIIZkwVH0AwIB9D
OEdaPg22ENdoXBCMzWejvfkhT8g4e/00jcCtRwAm2zzmKb9EmLCENufqbT4h2IJ+
AZ7//Pe8f4f/GzLhFBw6ZOj5ojiiU9D3bA9+4xlf2TgzflRXECQHX+4t5U8YoC01
rREdGuiJYZ7DUOwKPQE5tNhUQxcewCHFlV/HNA14i9Mq872vbbS/ghdZvV8uOUNS
GtgSIkIVpO4PrVkrIOupYVIPw89cR6vefTKQx/T8YyIxFeChy6aO1ZfQlNTv0rl9
auAOgCA+LMi4UNZv/aDJ8T6ykeZAx17Ikysyu0HajJk7uL7Jl6QWwyw+NuCM7D96
/5foQbB5DEHF8YRdZ+4Z0ggFEMcZ7OW32KCUf5kAOBkgNiQuepua1cCnNqHWnx10
csaGZ/TzAYALTXvxVpfTD/aB2WFrZR+ogeoquFzyhkgoa5jLCgeHiwpuFH1H9guW
6+CycJE4NlMpJEMeVCB4TqMcQwHzR5pPzHtPx+SuWbih7N6XajOm82EG0rr60W43
dZaGpChbQt8yLg36sAnvcMRR4WTWpTsbPHTaBQ9idYIsvxQvuc7qSGxPl0mq8dIu
FQ1dl8LLdM1ndVN+STUY58gAo9XZNz2rAEX6aoyeI+MXtkyk6F9S65JneNSJbnwi
cngWezqVjUS/UUEoeh00M0DN5UyRhxnf++i/8qUZSC+ADDaRwK4xLCn188j6UzD9
GJvEF1mfvQoLFJxBfQ6z3xyc7Q+llo794Ni6y/A8+VcX3Dkfij2crqI7udSBIpLm
qfAJ4LxByPPra+DrW6I7MJY6JjA1Q7Ji9KXgk65q2usSFbPr6QMrWH0YjMNvvin4
Fiym6FGsz9JZsDj1FkbsEmYBR0CkSVKZ1yNfD4I3nlDNhCVCrRWYNSwPCZxiP8WM
Y807oBjwPmojB1Mb+WkuG7xhpiYRwt7lYN7pTlMTYAefieCoc1WW7aeUGO0Pw+Dy
YFLbB/vmX9mdIZMIAjMguRb1p9PkmC3Zzi4fgVh6izDV+re03/LiVMT4gMKKZUqT
M7HTLhYXD6T+lBCWd9MllUvBvFbwiybMp/1l3R1rBOXhmbik177MXKRbKbxliPNo
CLRNkfHpP+efE5NjLKTdGt5KKdWUnmS69k/ap7AF2swgMPlcup5cGmOfO6kHhNcq
nyY9RhnNLv25f8i74Nhtu8Ngv1yKuncgG4+vDm08iqQhq97IqzD8kDWFNYuUvM7j
vt/UdR8pLWkMTVLZziCf7nca/3Jt4mUojJWKNJWeXV1uoAGK8kiiVXd0DX5y+qnE
kvRhEWLVfNGG4IKAsjLxMUaWZFP929K1z1qWsw91+L4JBvPhBGUieMnyz/PD+7xV
jHolTTTLPJkKZNx6fYUM/2W3SioPUw0L4fWqoNBetjE1Om47i0huzbeRq621rvj4
T0lvmqgnK6iM0EH+/hLmGxxD3kurMl8HpJ8hj7yGvfxPVmPt2rRyZIiUd9eGnc+/
t4BWchm3xYo8gWCpL7LkWp/7B6/b8GWJikSLtmlnE5BEljVbZZ4Pz1GzJApXCSvO
Tvof8VNzxtQOtcYZ2gEvQCbw2J+hSmVfFIGnjo57bZstpnEgzjKWJgvd2iQJ3YgD
TOJxIoZ+0ZsBBSoPBe7jfxAlBOotXAsbadIb74e4ioiTQHYz4/fbUArdYxFU6wPz
DLInABaeSf9hvkpg52h24YtrW7IxT1bTIpP5sSZCVkpFknb/qX2WMQZIXyyBTsNi
wyE+MrMSnILZgOSdFYCMo8FFg21rIGlsTICISsqteT1oFdY/SG2PTrgIupZboPg6
GVMLsRaPlt7trtL3C9Y8bu+uy0Ie/bfg90BKu9WB3kPs3WmkNLsOzIFnVrbXJ4Jy
tvsN1Id6JRpb8dvMJ/as3H5BUX6BtwrZhy/FGWrZam46vfH7cYMcyjW8MY1ztsTM
Msg1Sv+Wnj4+bPBo2PAktnd3Dv4FhGLF4YimIY9TI/vOuJFFEG23YexmAA6tXuev
EpveSPHU3YL2TVBKscovT36WbZYGsXhjfhIJjctOxj5X5TF329/crsPqQN8LvYnX
oUvxYOItlltCTOjCxMA49agSU89aU2ZS10U1oxqtFE/ECDG2scdxzESEm/yT8v0m
RaUg2muW+U3WWs22/2dh0oTiUVGk7qvxCBvG12Dlytzt+eX2NblUAszTnwTo368V
SGOSJfGmiNsNOVk+F07Gwx36erI2HrPYanN7osZ5VUKeLjo0ZBsuM30iEyz/dszN
CRaydgNf/hE/ga5afcVaDgcoQgO0yVbljN296GvHyRff3tn0TcWABiBxLHmKvGjF
F5JSFu8ZaBqzBmfQ0o9Llc2rv4Ie99gywx9T+KuWsO8Jet4aHE68xRVsyP1MSjoI
9e8vYooTby5qokaqS909BIKL6c1yXX9aYRs8GG/1xk/cuBVTPTXXlovxWn+hXwMo
qz2ZeEhitHMf+wJbFMItpnDnw56uVU1+1sO0YUY7f+KuDHh1fQ8jch0gn1AmQWvy
/AEjfUAsoKpbNJuswqKzk1CpHoCZ/LeYBjiWtfDTo3HeAtph5sJvVTq1aYjAeP7b
PsJ3IhbKDphrxHGdnpXML2dMLLxV3IyB5ldev2EP1/a9dbozCkl84raawimbA77E
Sg+jQPy7Y3H0xw9+cJ+102PZeNr6LGTmb193XF+I2Sq6TZ5+ajpUy/6RtxZZAKDh
D/8R2oXwOd65SFotGgqrOOXVE1PQHmeUIitzBCLvypakncILrE8bCEFlW43OHSVJ
3RXSQ5mC+xjyJYArGsA72q8Nbx6RkvDCGO+XSVAuaw5aBg0BqWJKofH/Vird6+M9
L9qVkMxyofoI9ui78xKdJGrFXOL02GIiBWWdZHPg0UBfjaold6Em2/i2Oyn7CXws
hs3/nm2+dOeg2ZcfcFbgRoyrr1cTKW4qTr9fYZPr24TzcGG1j5ynFBYexjFu3PLG
LGJ7ezcSr9+SRIzd70ibuGzcfywMFDzKJCM6gNm526nJfB+j3gq0mL3EkDdqOcSD
laNSXHdZTpyKQL5Od/4ZW4r4M0x2s5Xclcsd8VEkWC77mgFwNVwOhAyHkpcvRVn6
uQVwnXz4aJqocFOCgQDTyo5oy7KbvJ0XqVuUZg/IJcANWQhkoz2ghfAVRM0/xiPl
gNcZRlJQrMWPkNQslkfcq8m9igbE/2YYMVa4xMwyPu5SCQl1+mS7lovWgJeHUozz
yO4yRi00tX2y1bKRgnRYgoOQYFf6eW7zTNnLdSzsbTs5nx39WT7aSzS8Tzx5AInB
2oiCOIwnK+G3oIVImSzWZfDsTwaQVMwWkePFS4YljkNVcB4ZSbJ6O2w/ntcY0PVe
lUCe4QpX01uQV/2gMrfAcTec1t3bfuVb/RpXEROioARPxJbsCmq5HEf+A7wci28V
fcncrsrKnChl6zlOmB0hQxmibXigV3UB57X5KJT5ngzsAPpNNx2GvT8BYY7nS3Yy
W8DxXKYm7Bv7XCO4xllDTO37TuC8mTzwfPNsiaY0pIBn3Sj8mUYQZjKm0ReWS7qR
gkwMuwx/epmOhg1zHuK5L0KBClVFZXps2YASc0H7BAajfro40u48wMjvZLGq5C0Q
gP8xtx2UBepoVZ6MzOCv5YUT2HmJnfuVjo1uFc4FqLCeDSHGY/c5K1HodkNsooqm
MgOP77dB2HfTq/xg9Kgrc/vQ/ILJ1GYVIQTxOIjamGHQfuISKVQHYFu4zStodj5k
sCy7U/y7T3+Kr0b8fHzPCsnZ3I3Lv0iN9EsO4ZqzPzrti1kbzD6xZs3xZYWBEfJN
CXj/1nyTACUx747uFwUadeXMslE5vqa9y4DjNnPo+Qrm4OEyknKqK4VCd6kBns9i
A+TptwwKpI2KUh3HMK06r2JUca+e2RxLk8NlWdqCJRsm9ko5iar/0JtijWtr806l
DT+zPoPljb3VSmQeznVuOhMVSFTzJwsdg+/3YESa3s0q8nO1V1I8bAjdP/rGZwqe
XGZXqSSUFDlDFQyx2WdIrdBbvmDUHqmOVLzrV7O59mbnpimaZKl9jQCfwjetX/5g
fdNhsjnT0dS0YS+7cTECpxcIk1yWuJUJ/HzakybP3INwRDAuY5qSsS/Y0UGOxW5H
ZVjRatYuJwgU3BZrJ0x6ESD7v/pjXNwZdAdpgIK+nVaMp2DTYnEJAlePqb2ZbBXZ
I48xfIGbBqzk+Hx4hV2A6VPKQmt1m6cJv/s1n0Niu4Jl5qciXpm8NOyLapc23SnH
W1QRV680VgmrUKHYG7nkr2BJBcmhPJVEKJUGFC05j4H9TkACMp74r134jtabW/a4
TM6DnvIQSgKqD9mr1FixDI3xFikAA2mc7q36iWKcmrIIVneLnJGsjWu/IsJqV7Su
dEnita+YJFp63EtjvxG3XnsEZN+ET1ucvI5xrSDydwVebOP66QNEKMWLRwbXNrO9
Z+oW4oT8bXBb9UiiIP0346eyZKxl9/m0rnor0FGEoh6FfeEwbihAonPtQ/8PLvi+
bhe+apcsjSTYx2PuYWFVCXIZdvE/p1Wbc01IZS2S313GfPavUtgkOGTQEDHzUKRj
J7G6cOChTt0ZJfJvzPjygTEOyL6qOWTGFGaV1ifYqQraWB5KKoUI8RO+sG8qZQix
0+gij2nOLuBUoj1Zp+AEUScTgPWVYz/3fIStfJuEBGE5dfpqP3fYZhxv48z4tBqy
vn/FtB0VMjWFDhWGCAGmaq2cv6YZFeFjXvK56/++tU4Ydoy3sxR2IRHPYSBaSsyO
VKmLp/Zkb8hKhh4BbzctXMHI8NIbEq+Sfm6OGooErolfqama7IEAGzhQlSs33XOg
e7uIPsi2VcqH7zE1cYBheHxul2kMrnDVPyk8x/TNiE+/N3g/x36RNypyhUxJGv+t
DYTuti2Bm+MP/Ealuz5yYL83XgKCtLBfQPQ4qC+MLeMKReKDNPeIR3i69qjyvUjX
H9WJ/mEoqkA2gsnYZYyYPyvw42uAHHHq/5CyXQ2+IPOhp2MMJLE7UCfEgOBWnvNW
Vv6kZl9WCsGAleGkHXtYAdbO26EomtUOTy+elu5iKNp5uRHO5IYO1PREvuLdVLdd
V0qYvrVOW0dqNf4VpaW1CRv2iNGOYbf2scrMgcAnkkvX0AuBEErQhaEAfJcuHU6Y
0I/YiXNGk74qQ8rjLMRjUzZT/dxoofGh9yeSElPHBVLPiUq9tvvw0LZ2JhohghYe
2heNYbqbU3TRZCL5p1S0xHTpA8gcemkEFJ7CsHdB5p6oqld609EARnNPNDrBqmNr
EQhUVoPr589lGTErIpBxeXhtCbg6+fG0Ofp9/0R56Pofb2BNi6lnaJbijMynBAGL
0EWqQRDJaOKpd/RROoQoWMmrAvrwhZU9PHQ0DQDbHpIrMGzuLfcX+bCCy39oiII0
q0ebGFxLn3Ds5wUifjrC77R6G4rWpqZfXtxBam3LMPn32JUFkXmLcHb381GhCOmd
KKbdo2qVmIhcjhTYiCncygYlQVs21832qsYtFBr3zgPm9uBsrZnreVrEKabEw1hI
POWGsVLBrJyEtVi1l+s4VkAS3s1CfS3B3TxxnGniQIn2BwkVj708H+a7amVxET1O
76+WS9neJKkk7Aw3A9SDknoZzxEafASAgw356S5yWJ1ynBrCy1J3FXdksv0ubvsm
qqbG1gBp9ZxsOoivna2u0GLW1EhHZiU3VgJAhfjqdGMgaIFr2VybU4IO4dbYCSFx
okAH+gKGxf1dEyI+CjVLTcvfwhdLrxVOwBn5GadDWwPRyP9XXnxUG2JfV9B6dTvo
wWAfsUAR+/imk63gnzOSzv/6fDnOCTFO99oEmhuU4a789tsK84LAno3yMrr6S0/u
ukL3xumkpgf6R4Yurb4zEyRJwAsh4DUt89XJAUXPzS+ZoeNVuKOlgNsVFm4sWgIs
rO+TPDcbniY5oWQz0LU95adKiAVA5E20pDpjz1Xqyuq07+FtTlSbpC9y3uTRPNY/
i5/Lcln43NfRMj6qPSDP/oZIGgo5GQbOnullC/f94tVhSqd5k7Imz6uzsocMxsPw
v/XQgmieFH8GdSEkA7boh1aGROGHYAvA4/xirO8fduke+btG10dHD/i7t/RO4VPG
iRG7ocG+DmcPsvbZWrumx3JspcyBus9AyCFB0yF04+elDmAykN0PUnk75IY/+UNZ
di8b6gNsL+rbbeUNh0YJymY8+G3u3/2OjdoeulGAkXoS7Ourgzh6UG+6j0pQEicJ
KA7lIbU7i2u4oSmmvRjaBHXdgpiymGPH15E6L5DbioIr25vp8kiv2UqEHmYS8VYS
TTIrwogM+kxDys2lXWdx1Ey9ZN3o7EFUqPbc5ISn66eM3IeGCkAb/ttNdM/5ptYm
Z98u4O0lWY68jfhjm8VSS9c3kp9f7dItLuAH7mxS9MwEyRsnuFaKoKQuInecbtVb
r9bhh9jHqtBuilTjiAeWLVY44OBcscRdj8PdjfL3CUhu0GyErfsh0AHjGDOlIMC3
tCWVd66IBjciL93w8lP2boK5mU5LbclG5Zrk8jYODJpdD5Kjbt/9ojiYhv+l/VNi
p3Yi78LduZ40QeBkjeQZg2OUztLC4j7wqihvLM4zvrfQsz2IPSK5JbQFcuI8vkqF
w+VkEQgz0C0kfgPSbAruprGxV0aNLdLEIvnyWHwGJxbjl71Duxe0GQRaTPkWJEqi
/mMd9a39wQN9kbXK3rhyUi8HKwYgpytEXvZqfQn+NOQG+9q8hXeF/wYsLF+cHFa7
4NYhBuGciZp+kWwg6hjiIFhTZNjuQNj7y1gAHVWlEoPvmzmWpkJUGFu5dtcysw21
7J4UiTk4ISIhNFuzxBFhrY75s+13JOAFaMJCNrdA2In+AkGevZ2+6nje1tks5OZc
kA3SpP+6032XB6XStJScOfDtVpbFeINM7MRG1dJdOBjSKE60MhZcEZL1Ty7BiDo0
d3SGk2S9NpM6MeNolNnmhf7TnT35gNPkznqL+WVPsAnTyB8GOiZmCxp8OQxv2AV3
sMI+MSrs1GyOS5n6da6a8aXqZcT4Nn8SIL0pvutIIrfYrFTGvUCq41AyOAYEcXCU
mXePqF/v0aeGmAVt6pYt+vO+wc+oIn5h3WZAGkRqxzQ5jKEOCS2bMxrehX+fONsR
I6SWrNubnLDDWiuwEKrcjXMnuE21u/DT+t4RziLlKmNWRYq2jAOZ9jMKgiF5NG2e
1X4bHqWSj9zoauZxFR//+2UAs+aV4J3DneI8tQz+UvtYIdlVBi0KjLPXR0Iatv/j
cNcJWuaZ8ki8f7PXzSSj9mk+ji1kIfwf4lFj/d/XQPIAp5JELoSljrPmRji1h+VN
q38HInjBSWORIdhlBopHD2fU7SW93cqjRMEDfwSCRmySNTPkGNwuYsqZLCbDRskx
sOwneYiCmVeAoB4IMB9sgiJTcpIr3NbywgK8fFszA/wbRLwEVRkNobCYeRqekPnl
7LEGhdweFPAKdHxvLhYnk+z4LEDBdkU8XYmPtiSHq//8Qu5i2zW+F17+omFRKmQ1
Kn3W6d5D8IigP8mcM7t37oVm4Tf/vQSMrSwjT018TzKjHHr0TH7S9cHjjuq4XiZW
EWWPcV1JV6/vYLMSDxnkaPMne4S2DW5G16YYnuDgKxEimh0ViPM4u2TsZaArXzkW
WuO6s/26cvxawnCV58L/aZwZOgXGDKOBtlrczdWYI50rYPoDIjdY0ZQCFFyZ/Utb
4pe+mpmkqaZkKbpWZ8c53T0Br5iSsSrUWRW0VAKl7SqeNB0R5yVtGlyk5aeBhJ5B
josrZ0Ur1WVklRfeuhttKlH3EOFKf7p47JhN5fB6LWLGomqx/SmWhvGLCThtLQmI
0DwG6d4HpQngrSIbM02JpPJ8eZfdbmfr+jv9KFswfyT7uz48jo/TKJJR1Fd2M0t2
FEYgvx+kZvzouR2CM8NqfSLVy2f2wcyrflaL3hWYfRqhi2Cm+f2YFx7F4klGHuw5
OM6s9LAe9V4y9Y8MzmTYnUEhhlH2hweSbAWFdFsV+JQeh/aWxPHdhN8T08E5rR9J
bmhHlasWMybs+lYktM0yBUSpECoheZhyyoWnCtnsFUbXdk13T8vnoizKnY4PK+GM
HUB/FPOE5+R/CcbgP4+IAJUSQybba6xATz0nyLdPgVaanD/wKrojk1HzIjbQ29Hl
gYhxEdIK7xQKoAN6oukF5WaUIPH8V/WuVNSvt5WliqPMGCzyGQRb6zYziCxZHUyu
FkLHi92Kj4WOtIvTB508OzVYIRXb3okP4R2miE6THzEhf1oHrpu1vss2ZlulAKdZ
jSovRsv629P0ylbX5UpuR3+Nnz3MrAk2IbqRX1tIdrj4rdP+j0S8oDXlsBYr8U3W
u0yYtvilZjQeiTYxWw9qg2KzXn0cs3D92PSTsmUzeOTUSNr+R1ZVeZLEhaKaUKBp
wXFzARXOO5qq3ebffN55ADPOK+ttIGVS60sKeCaLwZISDtt2Sy4y0ytUN8pslSvF
+NfpV25Wg3WGiOJNFWD6MVDUPrD/IJnwcraY5Q95qD6AnbCG9w2+50wuqXcKdDWp
GIoN01D35JkBEHv4b13LTQA0BXjJF2x8ErVnArbLM1Og6ZyXE5zKudpN9gJe/z5L
aG6qhjmfGmR7hot6NNoMEvje3INIHA0HvPBVzpCeU9CldNusyJxBaeephheIQytG
3STT1V4M6l9vbUGpEcdWb/r/mwc9yyvPtEbM2SDTAFi7F1fdwunsDMF//pEjak9J
EjpwnvuLkAzkHdPvcEsUxmOJYn+GTkVUWRyyl3qFIkrRJapCCCqEqCQaJzYIvGJe
pItZlw5W1WXpU7V6i52zOQgnMiisJKqd+y11vK0OyxocSkXkoohOYCPcByb69gZ2
6sRlOPHewl0pwBVpz6AEfh1Qlropggacve/4IONK64uQpM2TtgHZHcCxXahGX2Dv
6/uAJFdPMy9UkzBFTVUDakBpE6cn8Xo+Dg4qUWxrkWlLTKj3Gb++BuiP3eGmPpr1
KiP1XkPBzFYB5q075d60q6+pY+3KHefMwWwZQ2FCCvHF/gBgvT3hWqm7y2xjsqUb
QIEI6Z92Gl8R7zSEnKOGTXm780Dh/KNXwixBgb4p5h946Abj1xUlPoNR6B4ypFv2
Ao+mmJEWSsZZAm1g5ejawtMDsbXKjAKDb7n+9iHmgFLzf0XAxRGWbQq67sSsyd65
QZILjstg0y1DywI18+HEG4vP8LJcd3j9fjYMDGHOrG3HlKmSzWHb1M2Pz7v/L7de
HYJsvS6NX/lYfX02ZEtltEPnigCw+oI96ivySTcwk5u+TtIbyJvIEX9upqvN+7WT
hVk8+NdbsrICo2va25lGR4zOPQDL3G3/jZLPevhfJFJEBzJCQml4Xr3614acx5aF
bFEfiznET2jZDfdP0N9UgOoEE2C6g8o2usKIy3t78gy0nMBrDo0gv2FPvRIZsjvm
yvBVFuX9txflDjuAD5TjnlshDayOvJTAozPhU0ddREjFPpfuWA1/AuBYRsLFtV39
winuWvflqXd7vgupsgc30iZVAFuUFWvC3AWfa2A42jGxKRyTXEtaTDnspYXLnGOY
OmnzlpOXb16zO3wq1QdW9E3MJBDRlz7uTmk/qL4uKSyBZG4/i/ds8BbBhpS759oX
TXHqAj2vLAcGYTnpJpx2LoD9j6PAvnR5DUsLW33yU1vAwB+BSvLfF9b68KnNaflf
Czu78/HCmRw5taLa/tlYuOmGuXm4DAr9XgC2gJknMeHHyuswCIFeg7deL2DvWajt
zl6Ui0VWyMi06p0wXR/XAJyEy/Q5MY8u8nTegeqCqoQgkCV50S59CjmCC/Gg3kMy
zSDL1JqrRNeqjsld0L5f9SirvMN5SJJKj8C0OYHMLF21NCftuza3YdQzAOOpcMkv
fywxfPX423NxWZewuozmzrtFLPbrYigkjzHWt0GQPx3AkpZ0szFWZJ60aa83Pufj
xQvY3cA4S2JRRW9KoOrBCP8/EwqkA6v9zD+UHT/cyIGS5nBeIEDTrqCvngfGtSU1
SeQz7Smy+asdAIHM1SSH3CiyktRgxSmBcGeT6AZQNk+8hG2Kiynl4DhhEWRb+nEd
Rnbc9y/CZNdV2c6kFXYIitRNDihs01Ujsjnx9blOYU2z6hkON1pUUwPEzd6UZhh6
ocmx6V+fpqYtG0kbb0dbUUpuppISkE5Cn2dpxC/XIRu5p2QBMS3uq7+FJA2nyaRL
49rMBvOfYEKq+q4WUaplfmyPgun8KY/e31svr+H+KJ04rN44KN9fZ8ZLgWggXuV0
50NqChLfRACAlGa2Pp3yUDXk7C0YZqya6z+5fetaPsCCm5aJnLSUDlAH1pHDmYpC
TYiMRd0tSRMduorbWOSi6uqUqDFvtUw7WbTGP41P0QXY92UPgizdyCN7+AoXVIHT
WbvWcSh3NE7L01/vYu3gvOKbYxxw0r/Zk4Erd86g2kZ4Eg39cRoh9DQ+mlyfBiN4
CN1SEd+2S4wV2emDGEdGpBkSShiR8OFVyE4Pot7oaGcLvK1K7cKr7WVsL0H5SmT2
zq57sWzCWW/zoAhUM69dkGrFYa9+TFXZILJVeQIEZcp/dF7Se2MpoNmP87jkspoA
qumWFREX+oUSIuJb52Ub0GaCW6FQ4LGTdCUpaEJcUmzWA/qJPeVyxsP8M0hqrEwq
9M8IRKx3N0YpDJqoj572xlpskXZg/oB2IwqQlBFSgAVp6an94TtoNiwQZWREFz7c
QqZoAjrlwuNV4IWUU77/ZCcody6ukMhbn6RiX3Uv23xdaDC5KaiWE4ct1BDNuq4M
ZrSPvDe1v9CaPYIT0kungKa8X5qc4ltVgLPYbVQnsbM7sQHx6l/t84JxqAOuyEZM
hrQ5GCllPhP8wS+6w7vicYNZtr9XFzjR6ysl3pSU948pCfnu+esAbHfx9b/cDzTm
Kd4L8ztu0hDE/sUxSluu0hBQaVGKTYVJgVb8aTVGDUuPLS0cmtZ9moU/U0GfMQnj
uCgHRhQUNB001Usbr/iwEjfVFCzeuU6bSgR526bdS8cq1sGa8Fwgg8zhLVg1ZvsP
i3s5jWzE8oKqMD43t8LdWmMUB0nd7QER3yq0S49KWWsyggr8zVJdpYGsEKryb6A3
UIDGTkUo2ekaxpvi9S5+y/mV01DcbemIyHNQfvNY9VVoFEc7ZmIgN9DTEYiMZVw6
mfwUcW1ppGiyO9FVD0ul1qHLeubLsyoEdOwMYm8tgDVtXzfkOOK5P42+nURPijkF
SovdBAkm+PPAFNI4eUoBr7ZQnREXCaPHSvLV7mO4EOuHhtCt01LmzoYHgsJRA1gZ
yolD0eHaqHhWJYGGvqnrz6FndDsKzYBRFysklr3ILE55uCK93Q71R420/90gGWnb
Ji1QZlFR2zthFRv+e+Q4Hs/GNCEzNGkqgAQlGSplGvQYnftdrS45HYXsPP+ynyft
6NCwanPfcgbXoGNJonrcImDm5V85QfrtXOV9zoI87FpdWom+oVgOWKCFQhn75v2D
KX37ycXLQObku+AUYIXIsQiZXWiA/3UxeM1wgvhq+sJZp14O4n4ry7OcNYwlhNmF
DABblyG0e5NFS498qB9+Lg9EqiHl/vqR/xOERm78faHnyTlqGjd7CQvkdVWD3RjO
+IzoQsuyma3WAylV+iZtgD0HQ0qC8/vFTi6Gosi4lNwKx3PUTmw7klkL2qVFigVk
KAgKVk77ZYCSF5Ew+BXkx4ScZNQj/TGOky3M02rd985I6Cs14nmpdufTDRzDFXGV
Sb1hcnxhfu5OWmmiH+HOl9RaI24p26JIsPR6zjvIKJ6uVQSNbH9MAZxGtEqkPGuU
iiKRBvrF8CeVLlhSUS4VklKWBt1gE7kobf8QBkFKIHaIPl3MXFHpGjXyx3rXX4oK
IpTzk77o8nn1acg2a9fhWhZ6LSzaKMr8ZfogwQ8j9z3o2XkHR3axjKOO2BAI51IR
1UbRHtIcDTK1Epw1ydT6wCVwlbtBleJKHFXRwPLE5x9jY4nKIdw6o4oLVr7y5oq1
f12Beky2gLebw3O+wJ+Npxs14GDFna5dA5TJiX2F7C3VyidhHVk1ulGHdOVAIT6t
rVVjON+uEW89bsR9ePNjd3FLFnPb9bNZuBsbWUjmqrOnhXtVn/u4txoXN+y4ZC2u
NtNsHdOFKLElmPbisQIwWcMipbRZ9HoYVsKNvBIbx295UPRtw2QQyDipuIBsHzvP
FCfb4sbznx+70r4QNyrDkpRj0AUpJT0wqP/0vB+WiZU7KFV8MKphd8HV7ck11YJ4
ZICWO6BWn2umj0y42BmyM5nVoCAF93papOTJ+r1PH0cV9eW9vN/aNzA82Z/Q5RRO
zPtkEeBgtojLqtdWApjLCZY/5B98ZSoPVz5mVsCNGTEhDXda6pNlhvaSzpBG4aRV
jsrp+vRYISNavjAU31iFWxJ248inzThg2vGEFALIXjC3lzUXGIJVZEpvrIi/UpH5
mHo4SagKGkWWORisPoWpMpgIHcQ/L2Kt+jsUP/EVVy7gh0Zgy0pd3HJS43inyFkk
7+Lv1Z5jOAmEX6wZNqggcvG+smQMjdAGDikVWMEuXR30CvMUr37eISm/IxGX/bCq
+RwlnnVZreqDQETadjuGy42nhNzcVgm+tDREE1w12GbFhKyaCKdQnCMH+XspcFuP
gC1Ia3jdaSqBBVHgwttG2DY91cH1qFmWhHipW/LmDNXtrgJlNgdbXTzySS8plSmx
cfdWQsB9LY6jWaDjKDhRE4kiJOQ2mP+wlQe/GglIIpb5qHELGiBXab19fZCp/00Z
ZN7EyKIkSQ7aQ79KxhY8na3e+XpcJo8poxbzpHuRfGx8NbE+oStqs9kg1Rt0jWCW
E8OScTsxqgZxj2gykWkdrFxbbL3Ww70K3TuJNjaFh4pOmYfGZSUcUxIME+YbtsX7
vb6NgSuPTsLXqCbg2F6MVU+ZhkMyMuCa7OOkhhojRe7KTGHLoBOBC20Lnt5+f3HC
sOM6/WcWAPnwaC9+PsNovPxru77dmpXbrXE9TO6KTmC+D2GepuyEhJfoxzg3BKZZ
ZTu+BwJMpXzTqBc+96wFkV+nQumziT4grkPfc/pMP+Pc0SDYVxw9q5NKWldtYU9e
Y6GHbUcQICaSsqIV+Imxmpgn2YPLQrstFouazO3Ganv6/pkuqDVbhJhmfoHxV1bF
CXbX0V2gcxm/nBIO9NZC+K87WRKlS/JjaTEQC36mCyBWUvVa+32yfMngGEDPYey7
YN0j+OB2sHe1XausJhcOHrfr2oPOo8DAM7lbgktn8UqpjEK2NnVgnl4zjNjVjjnA
+W6lzH/nc+F9oj8ctcYQdvWOrwGZwYaVW5EUB9A36FXjgrzr9UJFtL0jAdPAFrdu
G+soj9l7qVP7JO8szz9KkZ/pRnsMM6cnlZxoBqXSHpzEco72ryqDRNkoqSRLL0US
7iehNgAIFNiPYiKurgZEEdo1xvg7Bm+7QlAN4vsBX+PpEt/g7u3+NA30Cryn5KQ1
Wz8zdiBA8xYSamkhIjELJLGCl9H4B97dfPoLhn4D+dMqXK8rvmwSGp28tZ7cVh8V
q2av/KcKefDmpsuczo86c5mj8CezbOIYwwtMfmWPID62qhW2CJ3f/C3822SvtP8N
VbJAcYBbcu2qiNCFyAId0DuHMlitwXZE6vnaTCCDM44l34lj63hltLU6Ds/9eZfi
GfMuocRJut8tPmHUpnxmJIZMy3VpreSbc4/iNgVQ9Pt6KtptLEKeEhim6159h/LY
FNjXjhT3yDRD9NpXIPV6emI4aoOKoi9ASGu4lUONqiaGw4/jK9YyP7RV4HcqUC0w
p8GFrumpr+gpRuBVB/t/ravelMnnsRWLdWWiNQU0AdJh256X7UkBiCyd/aRdwggE
HIOEceSXqh+jBMc+fi3aYx+WNGie5ukAzHkBa7aXdEbD4nJz0If8RVvRxyRQ/2bO
hcLDdmQMfgKQ+vGo2ogwWbnCnzD/Hs0yOilVb7RNdAJooy6N5cE2hIpsak0Y0d1Z
OU3QjwXNivgsEyo246x3+DN2vekcVRsVt5bHZrdVjbnloeoCnocLDS/D+OghTAub
Hpi64T2OxSMPHhh+HDUxbDDrq3ITnZtPSA+KVo9K0eoAbRIyLCMaEEKvo6/jlkdh
MINuahYML+q74bXsqGVzJ2vKR3FI4SspO8bSQtwsoRQVIqmc+nnRP6Gdvk+SbFuM
I8SAbx+qJ9FEKRTvPSn75dMWax18rSENgC6n4vYY4vy+D6aj2N0n0hJySTFPlKGz
H/wwk8K5GjGcjWIXAIWp1V47fNpqy2z+O0jf5+42BHJwtyrF/RvNj0qTq5ffgcLh
cXKTU++OWv33qZIyOhZe27OhGiv6iMsQ/IUIWD+3NV/RGw9yOIafTzIH/vlO9IrC
eIGb1/FZp6smohUTzwGjFekMOxeFN+X/HqKAR1DE0iTcwS0e4vVCZ/MW7pS33n39
aH8CCBOCS5fDTqRD2fyQVGsNq27WOKcXYGT3QEWgp+2XVpshKFeyUjlDkk9HurwU
PwbVXzO3yiENCM/al6N7+YEYXjxfYcopULhVo/a/wNUaL2BCszzqc6G7bS4ouHJj
EmwTS5qRXWtNRF4N7VrWMlOJCa0SwhHKJiTUu9Pcrcf/HjTGztpR2bt0dj+a436P
fdiy/VKmheye/Ltth8m+UJn4AhOKuEk56N3H97JL/TNAV/PavABZ0x8NGvI/83jI
09BgUCna0Qfq6Ghhb5n85zVpeY8p+6hsq7Mdv/XWPtkw2O0JsbxxtLZlhRefIn+t
NaUI0wP5s8BFBSc/FftoJ9mQDS9olSLTqR0KMvAZrADH3xjPExFpnsJYv4RT9qFT
WPBrQeVBATgOjnBrOV2W929L5XuEUmwAF6ZIUlYhZxlsrj1FEMlTQ/21xdvD2Vr+
5gV+ik9F9UTNGnfLgY/UY1GqbG37el9G0hxtn/fWRI6xP+CDx7K0w7z5jO2DaxCe
6/2sSJNs2A57lA9D2sy6yRdsEt9LiyjklaBbP9QpU7eEPazorHtSuqaqAevA/8JG
aekAxybWuconkEyAuZLRf8AF2rSoqog2bUbBF1MegCFNURQQUDSitfQNWyyvTrsg
hAvBULBCgW2WavdGZaztjBd48rvxUaJJg4m8yCZ6YHQ9bhlmCKP2sTC8zSihwhKK
+w5ceYrde71Ds44kd+UhBCl5jp+j6ie+HOs9Mcql7v913CzEqEHqCfUCnvsi3MZE
XbJ3kY2DpRTgiOQP+qodwiyEVe4QrtNX6tfmmYQV/sbGcFwbprUB/uS0oKNj16Cu
f+ZEDw/gIYwjxS0/SnDPpTL4qGh6zGT+Cc9qrPJNnkUXzIz8LhJekuktaKTesgu8
N9k//rue8ajlOZazknRnQMgL8OOgL1yCiNUUuMalO2x22FWK0t+tYIlKDZcMPH3h
h2y2yc3PSu0Q5uEid8en/+Dojmx7H/fvsW1KnzgPmp6tcK8T218X4Eb/FKvSrY1M
c9X4VdbPweqn4bQNizArfl5CcV9EYTWniVrRh1ZgOtW9LrlPfwWBPlBTDgcbCn4x
iWu+yUg8QySVAFsjAd3DmCFnpWJmoXDtxPJxObpip7pTfVLWfek4iPf5XhESTn5q
4+hmGaZrsaDia+bm4uLT0MJPxTUODWo8O7j09k626nTS6wBibABlzhPOBuKlHOIU
6Qg6a3HZ5uMVlAO9qbOt1AU0HNTP/+CKZlwE+3tXtTF60OpOZ9wVDnHqXPxgBcqD
aicznq322bSEJLr896IDgrbJ73cQcLiY3PBbA0c+Ep+FYGWZQ7Si0NwfNcViLQm3
EEFKGzcQDB+fT1J60Bd8uQY7qK/6HBfh9MfvbP4OpgIIEXcU+wx0pZr7kE2mpBs2
CUi1CmLwzUpuWH2hwn7JgZT8BC8Hwe30/e0/f8bXC8IEl/6ZRRBXYvIN7eKPNN+/
29xsyZvXT0ZbhSMYoK16pXaFx634Nma2cUBkuh4I4XHlUgsPTlNRB5bi0Q+fmdOr
vM9C7vipGJ59LPlNQSIpypVaNBlrDTlsmefCHU77iIkP5+u++536EuhdD50YzLMk
V4jX9WJLG5lF1HmLCTLIcOBc9T9QSdnGD1vYNIV1V/tIItCyAq3mmXEUr8i+T3aH
Fg0i5IdbJrYuh5mHso/j9bdTweCE+uKED/TyqQQCEb/PEOZeyZ5tHRnp217FXPgi
pLtghM1TeXzSy7qJggZgzSI2N/aNbHxpKv/oFDzviVtdunk5dwDiFm3Mf/MQkd0t
BwOv0wWJN3FmrTa1EsAoMjx+Mjsa22xKjbSQpLTEofuAen19m1jIbxgiheeIsmyx
tHIc1L9cOzSnuyoL2TS0C80WwpnXb4GbIz4+qwGNHTl3sK1HdnvAEkWNIU1L2+HO
paBD60AuEF+9dRFYRbb/wBWXp2+srJ1GlxpyjK1X/j6K3ZyZF+6hmiNjp5MnO+kn
J2J9Egs0WJyQSRKkYDbnE/zEJaBohUSOFM9Qq+t52jdsl3J0uxI4zGWfnhK0UY/1
CZi30q5gbg9ypIsFw/21jZiaMu4vtB+3UkGSsiBjJW+2kLdyL2q4D6VqRQz6o9Z5
pm3Vla9YD8xX4Dv/6OD+OzUz1enQJcGATFAm7MjVsfXFmx5Y+gCxwLgIj3KwoZBu
OICm9INn1ZFuBjlx0jWcxFg4KyUQa4mFsyStnkyk9OshPNsV62uveNr1PT+JEVe6
DlxX6Mh9T6QU4V7eKE4cqWwwNsLtEHR/WmouutfNGHQ1koaxUuDVHocPkwRdxBF2
N8+Q05oR2/m6FvShYaTZVc6GiLXGRsYpwDuciERoZjMI21S2cUziFbiyuUNuRdMn
nOVIDkUFFdSdDsngfY1lvw9Pt41gfloNBHXWnbLuv52aC3+j4ZbmOgw4Kd5GUzrj
nrXa/FEH1pOOkrzJaJwBbvIvlm35g+MIdzTcguHiGVih+10hhJ5MGd1kKGpSb1pL
o0kpU0g5C4pziTjuwjrOmDdABxe8bvRrC5nQS7mrywIT7vU8/xWC7DqxAd+Uhau5
PPQTOdIRWSuV8Dbk/qbUW1MBFCGlDcO7IHW4M8uLCKne/G0z8Be4qBQ56PtJbHlF
LVL0gpk5CNYVFaFjj1d6jweVkgXsRxlCGB1O0hjFP+pv7Qh/Zw2212JySFAPBP2X
kTcLrYO4PZv38XEXCuYsLCH1XrNgyVLxEsnBFlsljR5NbkDTLvudrZLNbVcnziz/
6WsnTNIg0jt1oLofBJyHYjQtvlnc7ObR+RxfNCyMUwm9tBDv43C23uY04U7/rN5O
rRc+odDCKOiqZ1LLfckgNBXHJnCG/YWMWGk1qq5p5gV8vZHgehlseJsYzOIMtoj7
Gmx26Jyq1GP2nfZl411YgydizEychpc6i5Yn/Q8vxEJgDxMtj6OPaYSYrD/Zepd6
54z+cekrDZhuMxeUeuE2gQUPZNR5+roE1+pUiV3/BsCGOplbiiDq/wzSUgzlnQv1
kAAssV/EtklcSM7GNeDoovorlLpis3uoLicdhVpC0XZyX9bFq84UTTfy3GPizmhH
fjV2vpGa6MY6z9NRBA9zxBFfSRZSpV/cQcf/7ApzNfxKXmfQoG4di7hfmvyIrgEG
Hrk0SLNHBJfHRBm5VfzHCOVQPUfM50eSvPzCeF8N8+yieJTMIWvbC6Y8cWLahQqb
7LthoZBPfYcTeK3+OJpzg49M+9PLeB0mh6A9RWghJrJKO0q5Db2h/GxuvwQwRJPW
bqFrqToBJlEaZHEmyDlP9bH5QI2AEbtEubqoD/mKN17jXOo2HuqhRIQAshTp2QZ9
ozLm8KrgpOTKB0mBspkU1IhyEGWq6gBPdfo+/EL8pG6vcoQrQ11swEiGrMTec2Xa
SUUJk4eo9aW3WLZ2eK2fL5IO9RSy5iWjcydxPdn5r4KNgcRIosuw2vaUrAaF7v0P
fbX68ZhWdN5BC/u427iLtpz609clguhVXn5l0GtK1LybXNvPvSsVFe+qlyYB8C+V
DeAMIUjOuQfTkVbkE6k8bwlWrqtp2ye1atUlitLkekzUgBOG1mw2a+Kp1mswG86g
0cGF+0QCje75rcw05PVnPlzaugsZ+Shlt5ZWsWTIrRMJ4nsXmeQWfwqfbbkq9znE
KdoWFU3o9QiMqnCL3lA+EYWqtYbcyBRc4pbRd87ZSt+Qi3lMrv5mEcTYw+O0PKFM
+ayNVLhi0WuDZKN4U55qe5C6qOQRqd1fFgWdRbGN4g8/fansNGf78PEuiyAvDh/K
Z3Xt5fgwQfPt7EHhCaMKKD5LED1ur8zRwL10KHJdsWZhvfdTFOJ2DuV2LaXw0KS4
FJD+wTe5HeYrvWbiMcr6zdsiwI6fb91REq+bVVmto9oU7USAByjVcsrea3QdN28+
o+sSKDXNd9L8fKtR+j4qP2yfM9Rpm0BOfMCac+h/m1tVgj3c+bBOq7T3wc6R6/eW
in4ULH4BH3uuYvgkHqTzQh+kZaJg3z8HaZAiqSTJyV12y5ISiwofQ1ZLDVq3fjL5
w2hriZg1yzZNpqg+2XgMO9BnFr8GymBr0eTaWFswxfXaIyp/ORgGhnaVaWfnlj3P
FQQ02HW36rBmF9CYuDCzkckwK3BKRxbK6kLMr2clTAUXn1U+v/mygOQhaKRQh6vU
Vv0b8uIVpAiqd7HN+/wJRMbVHzGswVj90LzSwfdE0SVmS5YG+HHGup5pbGBY6UES
7P43OcoU/yd6JmZG1BH4Blyx1Ei0WKcxQOQqy61wPzHZWsH949FGQqomNgPw0nvn
OoAAypwaoUUDMYu9garbQwrvnzoSb3QSpgrkyoB/zBbSUhMgiko5bSY0519dH2ts
uIba1SsGoG7nwKleblZkZpk1N0dm7r2xSxrweaWJ5JADDff3wig7R1cCQwaMIxd0
9Er0nLqnelzIWCk1X9cEs3FiMUG9zJDSrCGx0fcYwn7Q27m1gtKJ0tAQ2Av7CRaP
kLJTA/JNCkHFu/kIMLsjRQfEtTUi+Rywqelfcr5s3RPCkoqlCKfk6p8bPL388Mhx
BoqVHWxWDTggbEdIQR0aPRwtnn0HfUKwrCzHy96ybEricfamUfgG63kz3cJIBF53
893D511pH5klp0ywZE2VwZq+u+e2BHws8JtsxTQNi1cOjjxjH7vGsuF73upSoPXX
e6OGv1d4I0YztuFlFZBRDn0wC22Co6niZSvIDxMpb1KyNbEaEeYthfF8bxO43/K+
HL9wEyedOIlrhVMJlLcMqj90VIzGxwmqKUyX48yrrDcb9Sg2x0p3OFXgcEJPwjls
N3yKcHEno3aMSOnVTJQ1yxznnCMYIKSotFUot+nBMEJ1jXsdmLCnROZP+vfFJXeO
1IRev9c7X826l+ZfHBDbanXv2ApVmI4tgftiizfXy/vdqS6mDJ8OTwwSZWdxWhW5
yvAS/w+BWuR8pPCqu6lKDUbw8W5DLgWIyjRS3uZIYi7Z3is2Bd+VEVOBmKA8ONbi
8LeesD3ts6nyrvUjcNferJJpImbH+j9CqcZZi9q9ty9ivQrtsgEqrYf/fvawEkQr
EgRfGDQ6jNRmtBkx76U+AjktLkelY1fJ0zAoOojSs/54q9wYRPacKI3oRBvuirbB
5lMgZ3LHB9mlQ5VezUIoGcmZNip2/ykiec8/0+A606E6gRKtoL0eO33ZYkPOR6g1
tHuPsE7Dlna0lPInlmWId6Ub1ciJ+62QKu5kuLcBAtwPza5mW3k1s3asxzTLcSNC
4Jd8OwF1Yi54UEz+Rhajg+T8rbR6nyYibxGCuvPhHnNZ31+7X+Q3gaeRttC0WmIh
kC2U0lzS819U2vItRINlPWLj64K3OOQnURa4BWos3ukLhd4Yroh+xztwTy9vi808
RJyPnrbr4twsOBhi2vI6nemen200QSG2rNs5pr1Nyxz5/bqukHmCRvwHQXcC8moI
Xw6rQ8VWMZG2Ieej5m6zcpfiyEpCrFzRv7ZUuI16EzgE2xib6PWiQmt1o30Zs2b1
0sUPKUQEmasJk8HTAyNd+jUi5RMKTE26gjTbMMHiM/90dPzxJv/58FYAKPxnTs/c
F0ZbdNFJ3DsDh98dW4wzYOhtnl7J4TCjGAxa26WouwBD6nqxFq6h9BSuyKDA7p0D
9yDFDYnwf7AB8d8b0io1tPXi+LUaJ8x23fiQgVMSDOXpkGg4IO0I7q+ycnjxRlw2
XPQr3UiTmzXH8A5NTcIdIEufqMeL1GIgGb/ns2acu1VRza7MR7JOxC6S4CmP/hbz
hg+Tk3j+wCY/PRdruenr/8zFnTGyuULxgFYsMIExj4LNfeDVuqxfRrFRRUrDqUlL
fqVCOPMLAiMwU0mYZO62fuBq4r8kXpyKVZTqdF1Jh6s9n+wlZQBcIezO/O0tngYt
3X5gOCjWuj50qsCpqJdClL0jLioFzrwHFtdg0DnM5iuVfHEukw2jdlo5dTrjtpaa
4CTP8GWLWCs3kxISIc9FG43t27cgTmuTrkG4knDKDVElkssVmIOkiMZv8BxzbRyz
Pvwtw77fa+fVVQmKJ+5rqc6cwzrduzr4e0sxSf6WQnoN4TWoQAx143Utvn0W1Muw
X4EXsAvkSfcYkEfzUoDSY+lnfbcIKZzj2H/wjAhKosPtpfz76EFHiEWItCnBXngi
xYsvePLXeh8N9ZK/CFVYshYBVEYw2AdVXUT6OmGsRLgPcIMuavPyjBaBa8tG3yUX
7UTQIkiUHT2ybj0n0xwpzjuLSSgZ1quCQGbQvK3cjScn93cLiOokxqGLPaF+vSrj
qHh6HODHhUlxBIToWgX+XjHuNOj55dwbRWuxgv4OZNxcshxI8KCoxNOwv4CaaNRi
4/zrMhA7SoovyyLFrT9Ux2W83RxuMaaI5nV7HT7SQPYowYeMyS+zJcez28S4NzYD
rLo+TcXx84vUlAq0OAkaLkA8XXJ6NGgXae1/w0PSwf7u/Se+t6E10ZbDsS6upNcY
6K9l4mzLU0jexBcRB+VoB0CtGf/J+NlZDFMGO/1hq5i32BZ4vj8fGeAzw6BFVCy/
mZW+H3neHzT26IJO3Cr4B4BXklThbSi4Uod6rN1JvjIuzgrb/6trgjP86l3D/o+W
bUV568Y2tOQAMQXrRkLjhM8Kot5NknKpL3sVJ8KVgPbSk/vMYbIpm9OV1F6WEeie
1BYXT+w/EH4oAc4GpYV5yBy6DHeeAlt0j0q/J6bj5ABfS39DTeTSe5ueivLJNOHC
f6D1S5f3Hk2aIM2QPXXvYo4eAecXTCJWJlyNwlWg20ky3POeS473OrLBCl88t3Ez
vM5fCpKKi+eQjw3fhZnf5jjFwCaGnxYSWyOyXo0TuCTJHHrmq56MJ3MVNoA0rgN0
Vbd7/sPsEahwG3/Z8RNWhgQOX3K9ucoxtYEXODr+wKGKzRIhs5RoxKfbUSghd9of
lac8YJKNH1ngn4YMYz/60NlqOXvK3lwt0JD5UyBsa/H4mZEj1yR6NytZmAh16t6p
+a2iVB/wdruPUid8RsYcUQlhmUnAb+LutYfb1t3vWO8j1U1QslP5KdQ4i1iaD1rM
pniRQTNZjNn5lzd+ppb0IT3+8j2PKC6HJ9pQutDCgXrChwQhOc9mohtNy5dHdbH+
/bQPddp6CPK66jPacGUz4Z/zTZ6Yuv9Eir9FSFhgzUajZEts8EClqWiL6rFsV36P
NRzsaoxRYnpVCal03Ic13tyBvCQpPiiOGWlavrEo/wUiTH1gj/mK8FBZWzpo8mae
SKnvRqyZtKGMxjPEp30dnV+mynPPb9jmtwS2ZB+JAW09coP1iRjTBqH7YAZpj7ph
mznLKPXpeOZKtnH3oy3e4z3TDencQLN7w1riPF7w7xXoz0amGh1zE+MPLBbGwU9a
4YLetQANiVnnmP+wK+cld+3yl40py2/VosPZ+D5uNbx2cCF3V0/gwAfhtXEigdzV
/e4r2cojLIAvgwOuVSnerJoMB+BNeD5cnt9mXFZt77ISWxmh1k+U9gWsKUFuvy5G
NHsuMR+bILmkqTezVeCYNSScLdJ9/unf4saAytirNr7wNXPokEK686++f6StJJLH
EFWfmk27we7Ty/NWy4Ddef7wBH5Dsmqs0sUvkAXxokRcwQPuK8P3Mw5w5P3tGQNe
IsKRECsf7j4ihTgFBXhOiqkSAfnHM1jWE8xYLRfaoCChqKm0V2DxGQ3uZwIvKTEt
+FWjxeTtzv6ugunBpdNPfqOTM3kLdSy2PkdxzPoSCCkTbp3M0xDj2QVn/o1Iq79m
9VWgmjC7LTe+q21/f/hqvRxBpOVFHfOvWhIjXEPwOE/r7176L1VEW+6XSwBcs5+x
ZM/qIWjcmcALNfpSWp6k8k7Ip5DEWYZpVJUmood6AF7UxXY5+QOHIfG8wqGfAOfE
lpC0y6KIdJNyuqhFo95knYINMKsaIikt8Do75vHgbSnPgbOYBsPPGta8Iudt8LM0
JyASpyzO4FhfjpjdX5bXu3FgQBt/HoYbDJs/1hNwOXo3PJWuWy8Aa6k6i/7tjs5G
tW4GHhLLo4ru8HqiBluJfIMnyT3bFmbtUhRM2gY/jworaXY2LPg+CA0w9124rpF4
Y9uCNPHEKkARzl5ZngkrxBMHxZUWrBSk/CU6/SdConl+22uw01QdJZBhCfgo1rzy
QpRD3JZSp489sdYqwDVeCcqVV0XIRGUMVdLGYJ9iwRa83hUab8ARecS6H88WhUyO
Fw2Aqfe37lBssZb5Tu1WG8/zJinWxvJ4owebJQE89UeNlzvCO61xjyQVT/ipUwfL
2yAENwjSXXP08rHsObhit2te+uaWGaTZJO0O2U3K9eRyxwrCZnWRpsy41v5Xyp+K
GLpSjfBNLaNvuZbx0LiQPPnFV3DoXqVRPeKV1aTc35fJXvB1ltkUI0ac1wClJl0A
fuuWTUnho+tQmWnMu58TcjyxecYJEXeQuFfFM5Q+qFJnNy95YAgBQozSgVepTzd6
qi3XqKmX5otOxqZpZ+c+Ze4NQ5Rjlf/6Dbg9xzPFjk3l+ponGbdH3bxx4DbnBeKQ
HwmEW2z7ZP6a/4vWMqpmL5ulSWW/qXl6WgC+J0DnAUntu6+BC2hHoNd7X3LB3uNG
xC978vAdNlWNsHHQDaQl1B95kHOH/R42rrMaxLzlbUwtLl5YPzFQAWWUoDzG+RSr
ku9C4bkk/ZlPtv3dNuHTcRWKGa/BaYOEyU9TO1dPHZLJWtdl50FoDta+T7Wl+jps
Uej6xA/8WSHQsmPg/zTzVeDxm986wc6Xonk8ASlm2zsLfAVuFTpl/eDlhMLZKaOq
lzNx8QS3lk4OWDj+f2rnV7Om9XOuyiMO9o4HaFwiJ5SA/5WkS9sP9bK8eH9Xs17w
j85MFMR0QuPKIdfrXtXk/IZGNRKFud+wEAH2TsMGh+rSG8H0JkOublzNAOmXwogp
c2Tcpe8dDiVREVx+d/5XfbYT6QSbc2j0qrv8YdD9hJoL8bTi/EM8DmyO7Yu5uzH/
F8dEp7xjTMkWy+EziRvGK3bQOm2fumnlLjXhJ4rwre7CBLnNENQa+8cZ230mXRpa
FaAH77dEDrmDyv9i0qrs7uglugBcq7FxQcH33fFKlZvFAMWWUyWHxZdLDMcWWtaM
L1w9YVGjPcPW+I6mssHRx5NsGF/45Vv8k6WaMoI6jYX6yDbhkx0wtbbglwAYSHGV
J55Axx0xq4AJwVTSmOKYcgb8G7rUtPeJvbl60+K5C03yaBFyd03B+fs6SgRDXH0j
Bf8w2KMCVQ5WZRuunC9CbFb07AqlyV6/gxkqND9jFMNcIVYfT9f8aoduik26fwu1
TNZSyZd2jJpgkoVQNx+0dTF7tz6bfY7tHo4fcEd8VpA5CiSKEAuBjZn2Jb4Cz0xi
PHodBBnWXZR4QvXYzw1H+Jb/5Na1B2PzU6PMGG8LJqIr+btHkZ8BwQmwlKVl2nXm
snUUmkG3veiUsT+WHbnT5W66x2wLKA7oqSDZIyhSMYIZpELdJi/anXuUUPkmSl6F
xSG//Q2sb4DoPHTN5/snCD1EL6UyK0iFGilYPruM21lP9xktNP5KcTzhpmvwLl60
KsjpgNTi5Fz0x4QJS6e95MynV9POSVjBiIPXw33fNcKpYJqhoxn1dc2A6UOrdiMB
+IkzaigwFlhXguxOqdz/RAieD4IJ3Th36Ca/6o1PROmDVxPRZWHnaJv2cuqtA6PW
aCm/f3s5kf3eyOUi9Fr2X7kznycj+Zt2EGrqwOeJ8NCOmJzJfLe/ZXEWvD1GpOkS
maeFvfeG/TCE9p5c5+gZEhIheWaqtf7I3MXmG/vx1uTwUqWz5BK/ErvRSCt9UMXB
Im/1CwzV2VC6CfqUWvV9nYSO2Ye2qyVIHnGVicuvUE0bhdNe3C/ZvEwClfN9VrUD
AR7wGV32IhEuqKBONaB2DsI0zYdf/xIw4MeVdvAE3JfWvgqdYDYCIrmaPIwct56E
fOm9wr1LX4GDjBDH3btLzhHuCVVSzcXqsK64PsIEHbW+OrB8hv5qW4CSdHpJBmvO
bo4aUp569fcszIxBVjMElsr2YGimPbY3j9Z0QQoZPqrBTigKCO2JiqY0JqEIRgCM
lKgebGvUvisHpyJxacANuP4fb9BBm25Q/x3RPvfkzWDaBMMc5VrbxqeeuFEnHz8i
r4dw6axGQDjMduCTxDWyGckVUjnTz1tQG2vBoh105vLaw+USxIcmAahiHk2TGhx3
m4nJhDZ3WJgETnCvnZ2XJalXhPWYJr9xozt0b2hHl8l8+KF2qRN5eeFLRSAfiFko
E+3qSsIwgleuP13DszvwFRc8m1DtGzYqPZQ4Bg4dCon5uOWQkBtpkh/2ubL/uwvT
c8bs2OtbQMNDAUfDCg+GzBgqy03gR0cXLkbhqpSlhjfBOimbjDMe+ma+bCB8YP4L
GRqL6EnfmOFQyis7w4/dj5D/F/0QQ9qu6n80li6nalSIsZN8V+4o3R2N4uabZR8/
HElGk9kbwSrKs00aBOYmSIJmqWUDmWITBDVgITEM2jbFdTEImUX/S6hpwKK29K7s
b3PH/AqeqpbSN1qMNOheTK6Eihh3HhRXZ8pyAxWAGot6MNrCPCA6vFGfOS3ZKZ2X
gkzyrikTP2aV5Ctdrrc4m1v8x9TtsGJjrKOmFsC+x7o6rEZlHpM6En4xNecKU052
UWzFnLqQBSiwIMpiZHFbzfr6pumaJiejxRF9pZY/zlpmOEYUr4YRafEqCZIalJBN
N02G+3ZfxB8RV9lFw/ZgAhOKlY7396Qec8AXy+886IKF5p+NPe8gF41SXM9Kh2XB
RZ00CzFEfFkNpe8wddUw9sM5kWM+fh7Grm2+CFen2QpeJFfQOFyWPvum/wwkshqJ
mFRHhOkDHApXr8j9ehP310GDuW1iGzMYu1Fvn1p4nyhD1RA2lId2nVVqy5pqEX9S
YQgLy5czDtg7OLJR8r6hdXsGAXu/0dp+nQNiQVQSVd2B13eQcomth8bf5ffg2rcq
egTXM22b4q1pTOW8Wj1jkDu/eG7ltsSnJqq2ojTp7uUTNbvEixLtSJ7jXIu/NO4F
0ZV7CrzJq+xgSKjww3yzqaSZxkzTiiSbD0XI28kMVLD4RUfLwLIozQCpQY2Ltows
iZLhxNzrt3SOTASInTqsqT2ojmdrXvWInk5r9jgHTwKaDUb6/SgxfY45xDi8qL22
WJIGimEvctMM4PavAO9g9VzJXYavAx87xVmKCNGG0rbzveAX3FXQt55VGcZaSH+w
l22U3GfFVut9Wz3d5zmckKl+i7bzXVM279akFOtYHC9csqHqg0TZjidxsuPsKzcU
2MkfpJ8gjZu/rEB8xasO4brYgV3S7yeKBYxKA9jq5jrKoIL/peORkpmV8DnyPEGg
iZ+KDFAXes9tU5bYLhvVQ/REpVrxZscwOaYjwSFs/do6IFm+CQhSIYA+JyY8XPsx
lIHmwJI0saZ9sJqZgbZUOV8sHYCCw8ChnTzEmjh/BIi7pZ6i2je8yBjUop2NotOv
EtDNzi5sZDb+lVq6WhBLir2sVavORQs1uXEt1VX4jwgyQA+zOHIszMS/lT9If0bu
BICKl97r8aOFfaLU5n7x9zUMjHB5PUeI4C2fu4678q59H0KQhmvjMy3sceVBE2cq
B3LHXvwdQj7lbDuxDT/YUoAgc3FlCufIavLAkFWezhlSib7+3V0372GLdVQEPhbk
95kSa6ET/Rug1RrGeE+418SI54x2e/ID2I/rvNNFAf23HbNVwVwkJD4ptj7H1GpP
dDTd8x+vvDDq++HA/9qqDhPBCzikCwjiu/1d6FNgdjJGvXRrPXpWXYa1C4NsOsc6
nKfMkzWu1zDVIHsyX354Z5G2LIYXe4757HuTuIjVSbO1Cb241TrfqCOYAYycDMWQ
mfr+XPuV2F4tJ/jxKl0VgBosgwWH9UbQ4o7SmVHSJM2lbTpzVg0B3LX/XnDlg+Dc
7RYkwwvAwuj7ZX99odTrjgb/nGsvXtkmhz6I8XftUtfz02/GlhYibloXJ8wgeYzR
7TV0tuXGaYOSQY3c9Ypc4gF6seJkAzM0M0moj+tCDIwyR8M1CSeCNL+EnJzMwkaU
Bl4TMET/zsnbxJv5nt4siixaK8G3ddLkxKVXTtSDz599BiYzIrYAGCDWf59Uofl1
5SDcZr+6cqcR5ygJx4OilFXEFhws7aRvolkTCeHnm+pjKzge+KPt/wgDzIH1AvE9
ctOc42ZXY20kS4wrZz+wyRgdSbps+i74aXzJ/BZkQTOIzdcEVhX6vy1dJLbubP0Q
BdWtd3A4V1CChtQL5Fg2Z+wJHi/6kNA+9T/KKnQUIiLRlOt0dEPrhc2UXX5VeiPM
DgBvZl0x92jxMxkgLmRYcK2gZW6hBXcja9BQOr0Zg9AOK4JuE83VjtNTEHM6Vp/U
jpdFZcmr31yXA7k0dE+AgOi8e30THLfjB4Peoqlt2jehIS26kftGF/qgcM2CmZWX
21zTM/lSbI8YtjVbRFHiXWmegf5V6uJwnwFuRhbjapdC7RgMhoqotYwsnBRFNyTa
FDg1AiK3YBbYgZcAxzxURVWQ/3kDDLj2vixvGT/27z+yr9Lk+sP6FRjrCXGuaogE
OUPJHynTcWyYs+UsF60u8sGs01s1A5XuTM3uK4w1HTUcHJAaMfRyi9acH6rF6PRE
KG0FQiowISRZSSh7n3Gg/cOMh835VrbR5QvrH+S+hOJlmCMqAlZnJSva5dp2Q6x2
1sVNufw8zWEADPdpMPVJvIK1AHmZmSyLhnBeV3FgZHsXzhbBGF6swIX76pDn1Huj
OeVC5vkBseol5IDUUvSpib53Na70XMMwIvgUOz1z9Uv+VMLi8pOYHhW/dMx0Dkoe
0VQDQCNfyRcXYCpJdHgliL0EnbvhuCHLxSzW+vAguxtDhWGPajGUJxymlrAgD/7M
HSWzDE0yFvohjScEJk0FDkW3Bu52lwuUaeWmpjjCVeekPz06K61keZhGSV5aTflp
r+cvqzIhmpoN7MKx+O6G//0phMO+qaSBq/Gi7rgfy/Ro5QxnqWQkBHmIYvYIqScR
rnHR7qh3YQZWttsQ448+KwophyjZP7p6APpyypFPRCqbpF+9Cbp9g+3SYNYvPtWY
ZzBZMVETCKduFxJW88zn1wpDJIfTDLN1RBTnR9H9Lwx2X816FG3TFCcNlmMhK2lV
CJFvzco3a01dgSuOrsQWsN3EOsh41vqa6hWtHGBZbXJbOb/lnoVqPWghckSwEk24
p3UQlEgUEeCH7hebp1U3mebdAaDi8Ea7c/Qj1JP/gW+RNHFzKFfUaMYqvFdApChn
jCFLmvbxSpfTH5bV02Zw/NVUX27KGf+wsKjq8GrbGQFGSKaaRorivCSYwcFLGTSm
9eGIFXsKsxIJ4hBwaHuiZmWU1672rJNTCxaMu4anpGh+PjX9696wcVQM5dHLecof
Q6PXGqDnynS4Xr6RuJQeI/uESHN6qhGcrcUiC/AoReKWFHeN+wPh/Z5Sj6pro34F
0ePDN5fsnbqpeNP/HPt8Jm1xCSUUfsFB5jkpWmkPHIAbCMRI68PZg8/32qLropuS
dSLiB8Q8SZV2YA3OpSZti8a2YHUpYt0ZynGY9V9w+hT1LbENpJPRPHyyFzodVNiX
e2zBf+ekMrPJydiICdPSXrqroP5/LUetvfeD745hO0Z+G0HoFalle5lw3VqsL5mR
f91cQBGKpxjg6XrJ1EUZnsCO6sjrdRkJndY9c89yXal5iFk9aLaqs9/3OtTqiawl
FSst69LShpLwAcnuahdrp8hgTo6e3Amdo38YjKqMmFBStSw0HbYoQUETdv4X7Pf0
00elh6LQF4RbswLvWm8tZhvHvImoOTUJEtplX6QXMIxu5/sv8X85Lab1gOnPebfP
P+tGFhHZPjbpgandhOR3fEI+bvZevHXM6i7vWNDAOwM3Hb+CMn/PXb9ZaG0zJ2P6
oc3bniDRx5HHNdk1iAjD9Ma/AnIH4Dg3o2ILNWi/2PL8nMQXMzQwqrHtIFCD/1mg
FKFGVIQIvD5KInxc+FSKFht6zs1U86pt3FfzjLSbTNOweSXJNmj9wGNKSTVrJ0tg
pGFYOYVo2XkycplQBTvNeH72/uI/6FVBd6PVLNUiiGCDIjgXZA5TuWAMNHXCl1LL
/92ottexvC+3pqhNWCPa8erZcWKDbOqydkoa3N52EiLyFTm2kuaZ+WKwzrFqn/yD
YfgyGmht+b+emiWqg6VBaiQ3e+Ke8G0IHofhOuQ1vFw8341T6DBhSW5rQc5p7g3b
wiEyGWL9bZ+CZdpfNBGHVVyHfPIgHgGt3rQcI9YhRF5ftFFVyTD45J1WJaxABuVk
FQd4RbEmQXwW3mtvdimno6ObVnB+DZN4KXf3ugu2UIhktm2CA6kMw1IQPZl/3lbc
ZSMBvTDDQSWoSGXtjVoU920iKsQLne1/dZgjmeheyuRx7O9Qf3Rl4fuW2GVzmVP1
VfketzVsciiLdTwC+PeE2s/sYEgv61raFCGOc3cAd4yeYOCjkpwXj96cL0EkaxwH
iJYcX4bRqZw5gsXPZSaaJ7Vazpki4mCNRPwJ1BskZhSz4S2inCa6WdqLwL+GJytA
dsWqrfybNfFyheOvgQnaD8UsuNRn8vjfIAz8EJDJWzRWE7jqfM2hAhHl7gq6p8WK
hf9uyYL3lex8dZ1KagXYjHdqRQ9epzhOcVfI1ZM/gOf+40EJV8+qbuW8JwHFe4lY
jeOt7AOQ8JrgR6igH/7LT22FNa93ENb8dwLeqkj2HFD57oW9dkHYuBn3YTt7DA5Z
DECbIr/fL6bcap1SI7rRp56mogxsPU07WRxmYfktjjLfNRIi/xfGqrD67+C2Iv5y
hpAF1KitP5ZPBuj5CBfjgWHsMXyPeEUP0nTl2YISlPLYmIue6JYgn2BqNFptnKrC
SEUmU6b9D8DQiI/1YJuhMbFdaYu4LcLos39sS91N+FpKAk4G/oBvmPC81yfCenCh
VsKLAqTrA3mVxlfDH4SDejkMP26ST3ef/P7xa3Nk4vpgSgDddDT7QjdlbEAxkT09
IXZoyDP5CvDBIBQ+M6aHijng60yowkw/L8uIPQIiHZIJJBipIjRByrJC/iXfx4T9
vUHpBi80hSsUj+lUyVCHG3TjHYKckWHiKm4hkwFigQQlbyZrLsLy2zMqVf2N8xUk
J/dFQfsX3X/jr3HCymRlBQahWm5GDrgpVGayrmaTbgFlxVJ9r8aNq3FF3NRWj8af
f6XOjat88McfmRvVsFhg6EhZF1oFukqJlxIWFuoFYz66I6tLNb1Q0pICsiFDwzHc
DUNEZwzj0Uj3/48aDuVcy+C+xSk6+IVX8ltPT5FkpbTcGPJRlKcGsy3FPPs4oEcm
ZbsSEQnBjBk6YmagDkdt3n9MWTPlxd16Xz0h22HxyZSg3B+W0Oyi4HYIoP28C4Ru
0KGrkF5IEpB3Q1Ppn2V+CUF+ErxL266rDl627Jidk04IF4JaF0fq1nqhRF+I8Vq3
lxKnVx4mq2c/p+9EtCzbT7zmsbeqJLs4o6TTjmJYktT828cKsOpWiVNqlr02UhsN
fhPbrJ+8VGq0Sk+SosCW9huJlNW8icxvFW/SEaL5zgaWDRgzebuSYY1qDSMhOGI3
5q3/1UoQD8zxh9IWOXR1JpTeBmSqkP7iuzW3MG1l3+v7DzouoKz0KxYxO+DHoiJE
Q3jZ3J+8/SWI8JOLaV5BPgNOTjJZ7DX5vAXniPN9Z1tx2zqx0ucnJSSm1ORqrThw
JAXOcxIpD+wgQmuGdRqb8RRo6p6CMkSOoo8hh3Hsa11c5hEB33fxDRH8nBHK8pEU
QvgPJQHNKqGZjs35cC5OVliKcuj70S8wjuk5nDomPk9P7RViiCrHYZV98U4LzPKS
LEQ9IUQ3rtLheIQh6+mXpADZWXwRUzCHx+6e6ct67dZA8WOzVQpLFVbi0zKGUsh5
zR1SiMEMz8z6JyL/wLpB5Z6UOZ4JO2PYayccpetiX7LVGX22u149lDKn9mP/y4to
MHtc4XiqcY7Y0XN3cCEXNyCOj31XVQUr1RJg4K4jo3BTyE+akjtmb1z8V1nXLyRu
aUlJC2lR1urDRjbLtgOE9ZgQMAWU//6zEEak+4y2XOGpdl1+NsZbxWhpEsu/Fopt
dGPUiSI8KQxrPGr8v9iZDIdKZfjDEpjivuXsDflY/RbaM/oQDd0JsY/k6sTruGTg
nuvVMFvXPdWp09mwq8r6yrBuUvGzCCGtzl+ot6NDPGHklB5ujlCTraf/w+5HRmK8
EYKkC/83BvYbCDowIC0wkhKi1rbLMHgWYxQeOT9hQg0vcQxQWBBkz9ZjWaWTqkLa
nModUsHmYX0aO3FyyBHVkv5r1a9KYFzI6TG3v0u/I9WLHYrd3abXcnUsw54XBqeh
+ZqNpCLlS4Hab2d6ddsw0LCmLao7LCo00eU8AabpASmbJJDX6rQUs+pUyf8gOPcf
24Tltt+M+lrQRdoxreLrLIBPWyGuIEnRdzSSeCnqvIJSRSmpQ/GJCR9JPuXzjDRv
RYxe5IixbRmjlC06hHfZQj9gogIBeF7FeXZf2zk7ys1zxZWnK3dIb33MnILpdOT8
+QyJ1lshBixkV6sB/JPpViq9jXL3I1TkStI2FdByCu6lqttGn1dsKc0TPW4Tpgs1
ic3be8lqZfF2gHtfeq0YcIwGTO353Bpe8EmD+FfUu5+1ok3gGm2A7bB/kVrbBrba
jowr/NbW3u8fq9c8KVwNWvz1Jx3xRy/WKDnRYofdwoY657kNCMG0NEw7xYLvcFRT
rYGbgZreGUDhAm+J8V2RhXFdc1VkFanPTcnmfQtCJLBVwF/EqUMWWwuKRQ5v4FjX
oeM3kSdyHgHsXVJUhxdBOXsl6clD9Oecb8dfvAtD6+xdXRb5uMHz09EtkQok/Mzf
Jdm6iF+GL9YyHdUMnGEdJGhBygXLo51Ya4ytNswO2RJzW3Q09m5jfWHpfYSMqtT5
GDEND+zBU9gHsHPZnHKjYo+gREMqbbwqTI5czRaGIcYOgP2jFgSW7Hv//HW2Mi3l
VTt+W73rTQiVG3DIkSTGl4VNxaE7fouhjJmm0sMVUmXDg55wh6kH0SeStfSRygJQ
0SEZVcH/BUFAP1TWgbIm0VSbndM/FEloOeNmQUf9chU/c/dFw8JfbiqbDOgr+Ccx
3quARdI2ZkxdwQmAZfyc0IbM5bYGo3Syhx3M4u+2DPda630PcAo+RBxEaI/8Qm0p
+PVxz35BFC3Y83O6QNkXziwk8vTverrCfGG50lbb8/WqIyj8DFDC5tP/WtfYrCSY
CqY0JzWz5a9DCg42jPJZ2DC9jgbRVHkxo7ovX2c6Ldj/HbECdGz4Yb2xLfz8OXHv
eDfR8IxCAmAYlE2pl3hnNkH/vv6/v7DB6zOfPoIgTPH8DH7Frn1BXM/K/N9xE+x7
eyAtGrfTX7hjPew9p4ZUMq5+FWL3/GStfB6QZAwFF0giMEiSHe7Kx1oVpUVzkEGV
ppbhGyEoxj1Dz3PKH8YCAFvjX1SjzaLNdZiYwMAjDNla9iKMMch3OtPZBR6x1EuW
7YgO4U2MUJDFV6/qdoodeGMwN6q08WF++o6FYiaeQ5aQfdo5NBHH8yXziLjjqYP3
uMvQSjN+Jv26i052o15cGfVfDymDDZw2HLLCpWVQCXpEMFVyAmdIviKpVfChllFT
IWNb6l0Sm76BvJRL24ThFf7hkyRAbpY0jEhG/k8PzE3Avtk0JpOXusCaAvowl+ZZ
RzsvTZU/tVjyCBUslHst3eWr2mWvicR9nLBOJOFTklG6OCMr53Vw+2XVkXy5S1XV
JIziKGPF8qnR6/b27YA56PBRTa7qVMut2KPN2m3QKJeyF4CxODFgxjotVQVzDBf6
S7K34vbpk+mmz9rG4NkAQ4t8XhsIM66zWRMUQjGiPi9V2GYVZwoAopeGxjGosWBs
J0a5MttvGNOn8woBAdjk/2Rj1gIXnVT8t9WeX2pp75kIAoWqkVtNRpJhOoS2UpBC
BnTpEj2+5c00zSp2WgFuWwIHYoS/yLt2JguE2QSOiJEm7Igg4cyVqqP03JVUgpRr
Yc+hXSoDTUPz+YyZhChjupbPPL5nm69M5PrH+LlmNp3obq//jF66KL5vUOkqhMBL
hw0PqhcsIA7qyY9dgCFI68Z6P3ziYwNNbxBnjTiOCN/5TCniYNmOKgb+mI4LTyhG
ScseVsie/WKgNPfnFdH3xK9SSNs7TuzxJj+X/Ksay/GXdR+NWC8x1FvTmB75jsa8
6YNO6ImTnwKNSJmLHtomXX2nTUOR+jn1zkprGvmJPUtyEG/4/vdVZfMA98dN6zHY
4n1h2PEt52bl1hYFc56nrwKDbo/g8CPtcU6CD6RwqPbHq5qxNMm+DFgv1pGvEoHo
wwrdjwXYIFqPbEBeewmqx/iLIjKKqmzYTaC6oGW7epGymFYDJ6c7vtvc75GPcx1X
EfN1e3MVlHRJjEiCyMWM6ktX7xOiv/pZG9l6QwBzwRuMtbENDMenA+NWvKmIpoZ4
ob7B90Iz5Sizxexru6ZMMbJiOd8fcYFqdAKJcynfemb/720xqpPDH1PuXlZTo8d5
+wq/iUQlrteNUTT07sKzgbHmimEuC4Es0SyjTPMf3kzahICVsPPbtA5lQeyN3+2F
2bonXYe1AFrN1zikBqG8ullcTx0oW/ssPcmQE+/9P2HzcWYwPfQDdSBp/gAkozMU
0gY9mcoBYJfG8t7cZG+u7dFK8R33sJ1pNQVvpQ4/8ub4hsHrO4VjfYMGoTgdYVsH
ewvicB8nvOG2Xejpfkc06byza4D8IWu9pBPqYP1Q2640O+ZbvXujzKf8vEC9y5yI
6BCzFPtGeBjPjaNsxBa0QmQD2la4X3ZMh4J/+5K8qaOrU6g4M+fPM7sS4Y0QKWjy
Eqmejed6lnX0D3yjEytml8ciknHtxJw9V1M6IuV4mav/rj3HGU1Q/g0IB+T1lbKc
KV4zy57QjHns237tRyyFU9ufcf7Sw2l5Zo2A42O7ePyWknBzUV7ROgY3AZajab9A
R80kRmQW/7erYh6c+YTUf7mPN6d17RQluZrZXzBcp/WNrUdanT5uvnBWHbhJBljV
j8t7IJPdut1aS5xLUBXzTJrCM/VIS79cv6G1C/OfSg+njoEksqukyFr9zngsytuQ
DRbjlZ0CWz9xa8LxhsC9sJdlXkJt2JdOf42wZ/t6Q3nc+JBcdvINGZqV5glvBhY9
lO0QqNSTQDj5EfjL32q3CZh7pshJXz5A3PnJms8T+R8SZEVoKzhPDnk3SGxVes1u
uWvwspxohGWXDdrqK7iGOr285n6yOE6q1C4+TsGJudDup4P7cVCCwT2EUmRriOYq
7VvQClJLBJAMjKD+8LkAXQUOem6ZhNERzjJnPjITWDe83W2511ydbt3cxY3X7D/O
J50rIs8MpXoK0zTwHTWr4dRSKJOdYee3Z5+M2lC3ti+GhX6wedJmIUxYPC0FxQw0
S1jK2R3K+c5oaeu6DDXKIAtTJ4e+L3WH1tEbKusymVyk0/Vf51ZvN5EMRK5aoOO9
FG57SPLxlVOoJOg3/mD6bmimu4jkA76XIBI/JubQ6/9rEQmU5s9CvrN4ewroL9b7
kfhymuznawWMz+KUfnGC+aCYW9Nf7iNbcY0c0L9zJvtX3xYc1Gpg6VZdkNlQQx7j
oI4dX+XduQtZJ0vCMEUckwwFYSj7JjsEW1WKmyfocAK5kx2VIMOQmZj6swUb/ke7
YYfDNzs461OE7HWxuMDZOvheaUrI0D9+URmcHpVGWpouOBUOjGVZWU8vW41hltHu
YvOLfDPeWsaCzYFkhciaetL0stcq6OWX3EvU8scbGp0Gk+a1HTleLBN+ZnMibJVX
CXRpUirci8bMBCfJvy4f9QIUGLaHOa+O6YQUa5hr/5SuUZD6XYw/0jvkwCntf8Bu
aT72tmvsWNSajDoPqn6fFlkw6qkOBKyA3QKyMmnATf+7C9skS45B7Zo9F5+z1z5S
oe4mUI1z40H5H6KMaZgbT5wPJs6MSnCJFPcAbc8DcwXw7d0jHICvaO7ix3JDH2rR
SjUviipb8BULIPYjHrddBdKd1q/s+/IQaV7ShhqvaCKPMNha9tcgpCs19yAKrPhR
834ROI07Lhu3yYq/CnHkANIeGTiqcvxju/ctXyesz5xIT2ZJziBszRXfsfJ9VLTK
EX0hzGpiO5mwaSO0tnBouvxbbu7/V60MbjBqss1Z7pEetJ2zSnp4WVAVpVczNqZx
ScT13NfKnjQOGfpulcvts9Wjw0YbfDQJZfB2Almxzul7SLO6xaEZf99bbOJh95AG
4yzN0c8orBJEM+6x5ThzMUAI0l0l5mCL3zPDtFQEhFmekhHypH2MfMS/pAofTugC
1CP+izGSx/Df+Hms90ppOPkyXaOe8oTKxct4NNqejZCUDwARMPIlrrDyfwXZf1xP
9/PBIpDDnxKqc05vDJOmRQYty/tWM9rTpuejOQMJH/WkT3XQdPCk4qVbD0sIfwXn
Dl4iTX8HNeVDEGWLIWxrTqKMg0e58hIU2veDV1EFXTqD0ipAPgBH5/CaK9LeNCC4
ou4ih8xB8foAt5uUaTR+xPsTZ4OInVjqFhmaNfkGNiSIldWavrzoitzzLDv7B8Oc
aEsU7tNyCaknn1Uw+iMKpi1KZ4YFSxn8EfDROBkACnguM6TcaRk4+/T7ooCiuPwo
3DVa2KJjm7AjNmQupv1siZUkQHo/3qpOE4RMKgOLY81aceN17cNNjOToavpoRzwI
yJRvOaM+wuDB43NYoBqNG8qzvJvgp9nQRvYSHh11MdoueaUXGsD9tc3odF28j7sI
nww5YesE2aZtbp10p6lMximwx3bAcXXC7BCdcrIan2U8VNAVzq80QJJMvOf6jWb5
T0oNuNTXloXEV+VRFiYyKETCBLAuxU2hs8hmcgv8rx88L+wDsOEOePZNYCCY4dAj
Q2KnCBjvkelQfsaCwO4NopUpykbIWuJrpWZ9Delm5YHYHu8lZ/VDBD6siE+NcYkn
1W/SpaIK/ypZwiBRQQPradc1UdebGAfKRPlYy7R/kLKQTooRos5FSj8nWLzsPnV4
qRovHdf/+v8W15yEwsC3b/g1oo1tFtNICGsOoa1vC7dj1p2U0jfIaAUXDPWDcyDB
+MGaVBLp8lAvEOHofNmV2tdtM32X42a7JvyUdhOoYiNsQH6vqa2aWYdGF1/35jcH
81rQZP/46dN4WrEyEEGnOqPd70AntRHm2RyD/gfqAFocGrxOg2hVwMBGf9lUAGmy
cgrKz2vls1wUv+GbPnsscA12bmGp8umDU8iBjRVycT+QK1Ng4J0ks18Zt6YrYMkL
gictIW3xS/8jiRzqjURqu6FeSjHV0rRYmiUQsuTqQYlo0h/xt2SB0UhoOWOSu9eH
5J+nqJCd5/LC9e5dYbmK+Z7Ir0HRDFm8ndM0Oj4cfiEobfO0dsxWOnXcfjQNMxtF
JOnun5Y0lSLsXdoDhL3LwG5FAcDHR1/EluWG+zzD8yOq3PG3YkRgTAOzzZiEc93l
yXS+rno7MwJmpmdTpGVLxL0GUWxLra2h49L8u6jcY0Kjkw+xMh0CK5451TLvWc2p
Hd27Fjsik8tG48QMphcqVp/tsxcM0uUT+deo0pvQWO3nTRhPVop4UKvnjCSNfIBO
yyHG/5opG2OVlh89OCf1IyLCvuy+WThsJbyFhzrz9wMTa/u9jPN8xAUE3CqpF35n
pcCG8lB6R+SHdCQPWNnopS10AMykIualSblZpuTQstcrGfdww06bgBdz2g1sCdQv
laS5DEMmTc8/wBwMSFgoah9QdedoUJDjNxB3LpMviSU1jSYVBWLogugcTJk2CDze
s42yfFc/X/ovVBy8zZ/ScuL2XesHJcG+hBZZVB8YjoZcG77Esqg8yxI6X7Q90bC+
DTTXc+zwC20uM2NkjSRE2oRNh2WRlSOMYfGQe4PsH5EMisI2RnXjhZ9kf46J6+ny
hJG0sRwxJ80/2G9j5+6PCbOflYcjcz5qWW+GzPiDO5uWTEn1pzNV1Gpv8/Nx7DWX
yjRQuDOeozmcfd8SmjfTNEgy2Vj9g9sGiNynoqLC/70HHi5PEZMGVNfZ1FGHxhv3
WlDdtLTE8+3AsHM4+3MJHyRwohFAo8PuPAF18bRD3VD8ouMTG2PyFZnQUsInUWo1
10JUuzlO6bDU8aY11C0vsQIuDxHplaczsREFqSiXkXSaQeTLKiFsKWXJF1y/KTWM
roCAID4WfKaRmpyGY5ICq0PXeuP9GG2oe2ErzlNJCeBcxN1em7SqsM/JPrUtVuMY
qL3vdXtpRP1Wd1FdxHffwEbtaq/XzCMoXxFha8GkvPrOxYiC5juxBVo8Bv0eGtN0
Tn2eyA4wYTlmh693hjECTSUCQtaimAkC6eUX0fT7Hl4tCCHm79hSSUYyBpUUFeqW
DTp91i/HgdnVunGoKmx921TA3qhFBgvUN6+wuOZf4YwkzAPYmAdJFCobHuzOV21r
hKHNzxNj5M8cbpEUz20hlX24xa4Sz4iMCcsJ6/Yt+Bdn8rV5lxDXDEZ5sIOnafJ4
s4B1SEF7qHdlNXityfAWf89CKh0YzsFIimgg3DNnU9J2x6lbRj9wz/xHSPXqEkQm
clhcbQIW8xPMNngNzeAIQDtn8wmK8gF9NoC5s0VoHluzPmv+lmehTqJfs4KJL5Tv
ynyvt2dbXUdwD1JMT8nW4UcsXLc+Y03Ire4d+9IlLa+ql6itJNgM7cRCdL6YrwhO
Z5Vveok8/mUGVC6fRB2sTUQbPLckQTdF+TYR38zft+6zRQW9EiVbd2M8YDCzF6R0
erhNW9cuM2vLcN605oLqrKYzuh1yI6kCs1Bf/y9YsKqez5SoyAbFu/ftW6bJMBk0
cisX/BoZZuBwPzY+1sf1JXhEZ5I7EwSFhGjSh3xo0Nu7+CeUF2/zH8Ew0Kl24Zw0
4yAqO16dzrWXnidsP6gDecdLAJWvh10llSBFHFnreOXNcevmHhQYneB1/1vdoMI2
Hr2LeSWdLTRy+O0OmeD6cniilYNnVJ+otPdvFSvU/9q1xMR8Xdlg7SOvr7s+qsyB
5bKhU6/ZGDW9MQwk/TuKn+yN4TUzL6T1zmQdFjtRF1FwljHKNOd8tffGl+EVHT9l
QEx+kaohBGNVO2WKf6BPE6TnySNpxbpZz1QVmdhjgAPTT4ykB5eArTGB5aUFYERZ
+513FRkhxkoO3NKzmLfiWr/SwrPJp0ZsDXPYAq6lk7YWDGVM3JvVQG3gmeDjMZG9
VCd6XWOyyOuLDqiORGrqSeGFTWMv2bGBcILAsaLKrCfxuRjl+p2EwxU2w3K4/ms6
WFZ4evP4NvnDDfX2n9chdtbZfnGTOqXQQ+ZoWq+skCMFDpcdzdf7WIRz5WeY3upC
dzS7qPflr/TM/xGe5UK6GYn9Ftzgqrh94RgT61l9vno6iDeUWXkXvsyVcZ8vzIE9
BhMUB/F75FCS0gQJjyNTLsNMYNcUN3LjhGcG57dQ2NJoen2tf18OZvMDsM5996J0
TkYeSjXE8AUEiCsOyr5p0sNIj1dphjm35TYEdKx7Vr9oOcdteaLiuU2pRBQDHyrE
j6afCCD9sWizFqsbcvd+pU6adq1qubosjBOnOpDhuAtzqn90Auym7BUJib31R25/
O5aNVOvKRURJxslkQMrEQj42gaSU7IIirC8WiltWYkGQzbeICFTiqVOvJfgQn1OL
FyJW7sDMbP5KXeh8fDoI9i9P+YfQbhgQE0P2y0QLvKPpAGqfvvLp+1G0lVtHHlOE
DGu9DzpFKppUTqdCuEElgX/n7CpMH96xjivTkoDMWE379qETPmJMHGs93axZzagt
bRV3KdTpK/EjWJBLJmNzTQ8zZB1Ne+x5R8cONoLl2/omn3vM6m8ayWwLMxoMwZFP
USwZ5PCuWtiRrwWQNYraJD+r3LjphnW1j/ieYPDyp98fLYMottL+SlKm1arGnMVK
uxXrhikBXX6joHjTTLyISsErS1+UmLHFD8DmKrvy7aTHoe20Djx8vQkrfoJNlZYp
5Dd34FsRBZS8psoVnbi5x/oKRG7CG2oj9S+glphjq8B74zh7s1jgIn41oE1VmxuN
moBj9JVvA5FvqUM9WtI7sSOFi07B/OxZO8qdoZHdKkyUcGtb4w1B5Gd6CJSQbHyG
jM635d3NA+N51nkLyj4Mz5/tFJd+urujGnLIAAMiwQYJKFrujJLW6pF04y8dIACE
C39QokoN/tmS39WfPJS8ofsDkGCwgzn3aNjuEIG/+RDlsJF6O+dUqpnLTlZA8XlM
+d6v2NL80Ol9F925gtLauYLeGDpnoeUU6Ou3/bWYd7fV9ChbX/WHutVvKl+9BQkL
IdStpQo+7NDEyrrAwZ2y6+6iNbDxLxcSfjbMAiT0bo9mk8eewv2Z03La/ZYMsUY3
vGBB9yA4gf3UFbn8XRmzxWE+nzvz4gJXCDApslz8s76LItrGrZR1hELw4bRI3zYP
eqxG3Ml515LdoTYA86LAj0iBeLGVdYq2Rw1CUHFVB3wQOJkQZNu5e5Jy++xxrIJn
HyNpmEGoiDCCvff36RdEJoWbjKHWOeaNNXV8psGzFQPUNycEVf8WZuU//E3Lh2tK
F7ubXEjA1QQzRiGjFY2zFQyE96XI64pS4gQaU5dg7/mGcPh80x1wgbep8p7jnGzg
OURvCNn1Azd2fIxcbx5GycwpY6iBmD8ccBKcwUqAtbL0OHxhUcMxft2qqp7olhZ+
WTAcMHjzJIpTEb00geoDOp5ORisag+q5K0H4PgDOPPbyBIvlu5E5Af06om4qIJjP
c8hbCfur5eDMMOrqkad62dpi5sXgffqALmr90WRZO4EBLghYhDXNgeNuB2F+XsRJ
AKVhqOVdNuFdzRYHzcF57oL+LfazCBcqMsMn9eGY7lOR+bly31twk0aWT7MlEMN5
WzEtGYNq/Cq+NB0mBEhbAOAG8P6tTOo0+Wq7ov1kakike02DWNmCObbVFxISsWCq
vbwO+Ci601N5wlDKPhfwTgT21SINl4b5jF0pvz0Vav814I1UWCvhD0PK1x6gPNi3
HQE5uHD494ey7y6CbfQL/T2ozocmqqKft/Ugcyo0uBgJrxMulevpWVUSg5joHEfp
iudt/uQrDNP9TOJ/K/snDBUI7hiflozD+1OTZbu/JlIo0T4ezCZ9uohI3FqydBnG
cXzY66ob8Wfl9IBrEFj2bFJEFmXgE/Vwdf4ZPA9zIWAGMW3HpPuzGriXVez7L9Nf
xVjeQ79aacLj5oGtxqrKtjhn8yM0/fSmov0qD7tDcWhib80HV0WjpMaz9r5wYlKU
/el1tXC5KfQ7zTw1jLe7Zz/lzq8BX1Mh+onwwv8aUODmESdZBIRcc5dtXrUcsBHK
fYga61gR/1ix7GGG19PVJic74K7Uwil7NzobH8mo/IeRW0dfM3XcrlKNhBGbGqjD
iC8KKiRVlXiLU1gXoNxq6tcLoODZhQz2MmJdvSuzdxaVzD8tER8aumQ5LcFZnOvr
/wf636OzbO0oGKHxRH4UiDKBO2h4X7/YcyNQSw5+edlKq5pm/czxJclErCH0Tx/y
vsW4EVGuGag2w5TFzleTxdKAOa0tvyEtEY7/mU9y+NP+u3EeDXS3mhH/C+T+eVTO
4h9XIPc01unVbUlZlvT0FIugMoedgQOuhwSu6XNHbJfnxN7Z9esagmzVzaoLxQtG
FSetwocACG7Y7GLqFVkURaCy+VFTqul4bp75dLFc9SOoPrEc15UZrOsYh+vWRTAQ
Ukky/Wim0cEFClnDckf6i/jf7bL9G5IwINJw0IM02bu4UETJZ6mTmHkNbauNYDJf
Vv7Cpiirtg9ZHHXlVViOrdBJl3NZEfTpGPhgLTTF/vYQUNkbmuKCg52W6fEBovKG
mCaH5LcLlm5GqRJQdPRG1erVGMhDucPWS+rSvufY+A2jXSlU+UlR2GpC70ilyVd9
r9Am+hL6y5hMA/rugMhrNJYdgs3sTBKOTrbZPHJv2K423z6+4mBz/oJQrMCYbZAz
rBEndDKMZ4VaFpfaBKsDxovaVI1QE7AunteMIbF+OjRaL2mseSiTS+GkbmXg82dC
GJlacKJohWXmYXUn+NpvEKrR09Dzytr8RaCYfGntGrlf5TBtYAUN61xu0GktDaWy
HKrjNfMfaPscU5NyfthUlc+81AAGcc/9SmkJFwJH+dSipQq6Q7vAGUYcPXYlfyRW
L9JhcWvtZsRI35iagY1YVgXrnUZ/5FRbSnIjhzM1qD0kE8lJwe9YkILGzbvGC6CC
PYKO6jXkHO9wDeXDEINdy7n95AiR693Kn/2cZ+KsujV3dyVb66/cfQNkQDBRUxl9
shixRr/O66pvCBw9dVo0ZkF9tDKm42i2BNTMt+0QbzF4wA0p2RiDqRnLVRkR65G5
dEmEUmmdQaHn4iCQroMB0SVNirlMa/hUUaCVagTQqipFd0pSkA3azjs5xLt92awP
kTByM3vfwhu9JqmTds/IhGXWsXIn9Gz7A4W5a+hmHNF0VzUBP/y2aIVYmTTx/vxG
DUm5G3Exq33efjE2xh6v8pgPH3sxjj0xYEbgjujDnsYZRk81yfMaCtTZ4Km8NUON
GigcC1PjDIwPFTfb4VBr9i4mBAv7lEQRKpQx8A+KHc+br6GPEgALwyy9yiinExW/
CqIBdmZsAvgJiOcesp0sPaJbroyLFLjwtHP3B0ekPop2PNXkUuuOzwEaB8i+W6GW
laHAHwfmoe2ep++S+9t7jZW5o/VlWeEjSZ4H3P4jU+L30ZjBguoPyi8+/zTS93TM
Lpw6fdMTnhBNeAl582D7qgDy/Nnlk/UVBf69lD/l6L2RZhNO7yGLv8Ht7Kdd521X
8Pz0+lxlIXG1rwOwc4n5atF35BQSJgbNaV/+NRdYXkMRAZVZuxs03pH+yqh+2Y8f
LQ/NTMls+49shOMd2TXk9yTCFKmh8TeSxISN1EUbq0Ky1SLPKNTDlMSLvrb7LUl5
DYoWMX4UHCZkHyF2lDi0ZHNZ4R1ELvVPo/OjZjTi2cLxYHRokv7kdztRomUDnMp3
hhjDQxPdbv1fJIzS5ZImtpdfB2zXHMArVXkjlADIG9dJl188/wd0W+/taHNpyEU8
9+ozF0QN+Ykw8w5cd4hHLnRR6iu4Efs56mSIrC8uaru2zQtGAIUrlwbXo0S58vLq
vmP3dgGa6Knjuf5OsqhI4YG5KaVN/BC3ZTxIs2wIz/rv1NEhKPTspqcoETnpm0EZ
dXc4i8q0jMNaQlkYpbKCBIviKWaHdj7gV/HAeeD3RWDSxxmZoUfOu/k23peK4m2r
81sHMaiOObizpkKw9GFDgU4L9jSjvaKRmXIYvktQc+GaKSqrPbOL6cdLUZX5zmKx
/IWfqUcwkWKBHLWW3vB1lOFa9GhON3VnHaiM80iDcMD3z2ilaWKyyi1lefUideL1
VL/Vd9ngVmXwDZYZe1dEOMJaLVknyXCoEKlpxoz3TwnT1cU3rmF3DYcXxHJQrWd1
hacdwpYCKaH7UV+ahV+a1RCAELL8Vy74U3EzhfrlC3dH1OMRhSzmZkOZOdwfhEK5
3K2dj/sWfKKNG9prp7lgPE6DYDcvhNY4Nu8yqLVOYgv+/UKOoN+GSVLICjW8IA/9
M1aCkc+jaZfniHXuAiyiXqNd0k8slpRtTn5mISBevAxJbDeoJc0xT5Uvmn+ePh2h
3+mCeqKpm+Gq7fJSZUuiXSt7sxZfSV6HZ63vethlocihBcI2x21B4+QzPyRqzWo/
LcKYHy4L6BNuBSpRx54DEjxCEP3JDlUq8NBkyy2OaQvHQ9xlKJJtk/9NUzObdERz
b2X7EAbhSBBxwWqQfasBLOSsMKwsobxXB+quqdTq1OyT+3Dgy1vHw5jUfj7+Wuf0
pfLtl+s7+i/pfX6R2d2bOTP1yDk8GfSGZ5h/5cEZRN+cxIr90DOu2xQm6oqrA6rU
3l6qEyRtsmuWqzxoYQk4mtencBFI11PBEcjkK/fKoukk4XprpVkdeHGwVfqm0YFQ
/hIloUlfasmcS/7AXqjNOJh80fIT/VCLWHatZbsPbOljG+XmRv/jM30g3H+3RxR1
JyaKfQjhAxBWM+hQIZx6jlNzyU4lm4hqq5DWhuXhMWuMPyR0oK4wDtK0dGzKWAjw
r8Bm0BuQYvvwVjhoqRtWjHW/KBFBDAInmfUQv9MjugulAUCCvFKK4w0AOqgwm5La
zKNARAOTWJPtv/cxbFRz/cmb19e4IJb5vhXcS+wzNfGrnytxFPpvlASbdCgC9ItF
rV0B+Lv+zP2rxM202f+BYHjIMhg9YbQ/WmnQXs86hVqO33iNhqhyYhaeUfxBQHWm
K2+qCJNFySMwCsWyOCG9xZenotPvBZlHqBFMfZPZE9Lp0wWGSzEcsRV9YY6pkv2R
tD9r17sQue/v+sxFBAWP13fZY0N33Xdjdpx0fqu28IROekWXyFL8svqZ1zxiYh+7
QC2iEd0A7oluSSTeZ/Js6NXErX+t+LIoO3553LtF+mWD2vt8Z1ZpcbrVAKLaUqCd
GEFPBe9N3JYPG8GRCysZSB9xY1zqdMZ+ZilYTu6EfqN31YAABaNF99UiZnOWNlCu
nPXoOvpe/Wpsz1jbhE2RzwULUHv8Za370NkRkeGtB5KKJabAeoNsoDptN4ukNiuH
hpDUm9Irgse7F94z/6GdnIp9GaBQW+J4NYaGbaj5XCy8GZcHrU1ppH8p2k9cnpAk
LPxCi7nE5eyq5HU/Y/6GXsVdV+QPaBcA3b/3KlmW3Vjq3wyc7D9iJblqF+tGpIvt
VL87JgZ5SMA926BlAAn0Y4K0vpSTgDk4wbG7e8esS4lN5XaNnoUJIEH/lP8bjoCn
mSZxWRk//hW3pNVrH3FEenpeRaDBNRMNBKPKEj8RN1VHaLXD59fBB+Cb98VvnT9f
WDagr92+xTv2ekD5lobbGDUMLgLOvCmxMnNrOCwgYoQk3ZafRSEpaaLpa9E5EXQ7
QOJzEvmIwMn/hWxlL68S1eBbs36+dLWED5ZCsrAWcf5d4U7ysCdZ+CHlJicAmLA8
toWyHQ4qkm2s2Cis9Je6tlKCcs2UAf4pMGcIWxQlEEZYlfWUtiNJcztFSPgFhZaN
BCT4X+w3Ik31hBJmgCPLix5k8bN2P+XCa5Jb9BCbm0y60/StSKo6IUGeAo57/Lb9
zG8IaNryhAQzWwNB6SrjA+loa15nBuNUe1rz+efrvAt0z8ntp17wrN+vA1VLNGsV
cRDspTu3/QFDPvGEP/pKCLcbLO+99FhR2xEo4BmJk1NA3sGn93UGikuTRgXcsiHy
lPaEOm6HzyLP11+DAIBAU0PhgJwZzcT8oyHGi8wYxq41GHX8LWZIpq40CwcRHL3V
EMDQYc4qmjOv+Qh6FbUeXAVDJyoaQT8m7xHSUJuzwbKqvFzkXhpweyQgSEB8lMj1
AIwHnFTwrX12uPkugBoTztHwzz+KsJ9egAwHGcELjMCXN5bn7yS7cr25PnF2ghc1
low32d1AWjnGhRDoztCXX3BSpwJNpAfg6gHyaqnm5WdwvcwWADxxJkPelxZknjXL
mCKYtBHFkxc3uesb5rKN1YKyYj+cu17qiP0qmHJBgh60c38jjxesvLp9xuFXLmS5
d6n+gyXCQSTGbxMtSPyN0Wempcco6YB59+IXvVm4RebbSWi8SdsXwr8fCNll+7zH
E3t2uBw9FcjPoDbkwTJmlPrioZBQcjnLTEnQhGnzhJ14vZzM9pQ4pqRyhK6IBQ92
nV75PQLu5CQJRJhxLrPDDfJcLWfIdeieNhHU3KalsTrTt+q9WxBNQQJ1IKawmGC5
xZ2Ynu+3OIxX609B3+I5ZvHqw8jggQZQdZquhOh93+L3qp1sEyFvwMSjbgxb0w41
H6/zPlWHS6c2IzCAgGy+2jXpiHaRVtYJfk+8rrEWZc6dwspO9twDR4LNiSkbV6De
13RfZ/FVBCKsxXAqIGoZh3z7REv4afCaRHNkcm8rj3FDwkEwv/xMHLYoFWEpAQ1G
GkX5KvUdYFb3z3YuKlUBFDiaFp+MBchQIxxZL1YGMcI3M+auLDppweBx/TDwcNKo
XCftnlVlAwL9sk3rrs+wGLpJSL48RVS8WwWl3t1Izw/f2MkMlAnXs5jk9udX28YN
9MJmfZQfo2k5YsQQnzjXkeSg7Q/gRkRYF8Dp72FEMqO67Wuz9/Px8THrR/HkfPZG
9i9cz/B9IWTDusGxPrnVupHljiAb6l0FiWRJoE5XciuhGj+xn30lsYcVPhSgScmO
M4Z9mxzmfqpl8B0BY/fYsIwAGzdhb/NqjhApL4m4/da+DiO1ZGUR7wHnU8e5YEUl
TdLmv/EiOaqOSUpcvN+fQ0nHVJLBPEXgBgioELoJ5p+oXNCJpf1ppNwd092NNPk0
NZmX8X80cDxLSmwCUFFnyXvIr0EWBB15olero7iaCYGv6a4rea2YRHY11ZmkpOD5
CloVQZ8shYmEdQ5KsgUxouuNBtoKey2YqIhy8i1meGyFOyFIMEYDXK9M4jX7p2CH
Msu6fZxM3cFrxGxXaPa38ewhdY762YaATOZ9eUO6D5yDLQf52feELraKG6ZOKGm4
7G5WuK6vpfSZGPcl/Q7U5E9XaRaZmiSl4b5HG5UZo0pjOUVxjpq5cclCQLB0bxXo
ReTYj7IH4RbEdXFKnui3L82uhUpT0KhvqajecrzBdcQ4ZpKMivFzKKIBhrztyvLH
9p3A5ZCyeyO+NM+LC89a9vRbzE0wp1YRat2w2Rz4zrlnMc18h4paKGoRI7A7BqFE
0UH5OodTV5H/T0JoJrFwPlT2L8rMSQl/aM92xZbfP2zmiAm9ze/eJneCPmyg4zsQ
X7jd4OrVEEox7OmpURl3KdBjNNDHleyH7t0Lwi69+8FzokIbUVeDotfWd//bADBT
z8Q/kT3YwYvW4IC04+4jgy5+6v+DECxwYZ41Q46260jttfxZVmY01po5N9LJ3qc3
Ev9yICXpWtuMmoH8AxoDCqzT1J4x4j7pKRAr8iioOaeClSzbmdRoqQPfflRjr5lx
jZPe8nt+YaJZatyNDa6MbIiEtn3KOttOAcv0L6FECarTsPxNNrY62k2tKY6oa8qY
qN00sCaEILVZVXlW0p+AN/L5OogAeBfGiOUYqix0J2t4jIQhtfK4KNRbdio9ejKM
G4ashvim078PEvziovVSkLcDbX9SjEedSyt0kqVESYYkZdkCpL8cZO7o4BkdEcas
Twh5f4tZkikAYURTb7EJj5HZWCvgvlS32nfI+rLThAdVT4m98cxBcARcv30tSo7C
6BK7oyYoywlWonaHTE4IYU03iBCDAbv2GUrLSm9wuFdqkQ6edjSHYRQ5AOPfOUGI
nz7PXnX6fXjsY7FdzJqUUQhBy6dxPwSkxD462rE4zHCpKBXQEyp3uUjhmqty6ar1
ipFe80oVg6HEL3l4pjYMOJboqCe2bhETzzaZtg4xxQ9sj91WelWn4ZglU60cygeq
a6pVQhZjK5Aah6qVmL9elNp64Fq6KnoyIsRwytRT6Fgx1yDFqchgfzEG+pVFYbBD
IuFYVn31OvZHfKyT3m7BJjo1MTBRLWlj1DY1EEzFzzjKQkODkcxsqdOo02Lpnmu6
9KUGQ+AJpwp5ElZARlta5OTf8oYfUvk9vEJs/FDEuFYvfPWmV1Koyx1YWP6+rTUG
o2swP2yf8nIk1OAqTewJqzfxh/oxt6dg2mgAnsvKJyYYmUZGoIA/ZANM5hXPW7oi
wnVu42rzy7iMseGvA8uCOmCtf5Q6X31lwfp1kPznrloTNKrMwC3bykO02Hjk00d+
WF6fMC0YJQAjrruzakt7i9z/BkygYp3HTjRG0ab8sxVsURFEjFzOK1Rc0PWiZp0S
o0Qb5yLmt33UIRb9xPTTmS95vr/U/QRpgAs0kuhUB5ARDsHxXSFMTHN3UCoClcZg
WQVDPvxnXrA7BkqNaQDVEJrJ0Ewb6A8ECWqXxBWbiftLOkvUw8TUBSNs6sazrQcv
qiQZq2L+BzehXEJNYGERLUkvi8K3vQklQCesqbFQwLaJTSEwvLIa3XvxnX8h41gt
gMiol0g9gAj4Q/Di6mDxkMGaJb2VGtbqSbQwCCjs6e35J9jWKLL9qoGGEn0auUlX
j5nOMhVfIuAcFGAeZ2GAdDssX995MDhw01EaKAqnUCtWtWYBUbK4+ynYmauwYcRh
LpSEeNe6aCuqe5Fr1BWyKyCVZ1YK9i+pFG66VjVIJESLbBRrhV5PZ32DIZkYqiVv
ZPoOnY++t6dHvu1wRPFk6ZINw0r2vplptA4wRqsFFaeqzfrQLIuCHFIcH3H9YEp6
eBen/ce1lgdIjTadusYYPb2PwSnECFstydG+GowqDHOiVpg8zzoYTpiBEfyNeGCh
nxM9E/dB9ouhcLBDnK2nV3hbaq05mIDBwpcBMLKnO4WLVSbI87RGg3Hi8oPmPRg2
sufZQfCkd/oEmy6IqZmKFOP/jnQpcbg8+vZFh6CB8+Tg+XXU9Sptxpkuy5SBgJEB
uZ5/ehYATEOliBxPzn+g3PztFrTfXIjcDl1mnfJ1VgQLsFjHRG4TIUNPpjnwOpNm
Jseyc9JIhuC2jrNlLrQXMUtYS5va5zuao+yU+ytUhBAsoM97oxZ9+sNdM6QfBzQj
9sZ9E+ZAei8xO2pEWt0X22LY3fRCGOiP1b1U90DsGO5R/uU9tO+RLLJj2QD8fvMN
lM5dcqkq09VdSs/50MRKIjlTnEAWN6MG/MCNA5AiMhWMwfoeInL3K01iT0P7yski
ScAb45cmaSQ8ZPo0k2IaYgnic9dhpkY6EA8Vjglpn68D3ujYjZR7OKd/mNKt22MC
OHxp2l8AXccCs5hyEQTD4vdnhRsVTMpt8jce7jhKsPRhWeT51fCiiCK0uThQXvVn
koH6WJbEYmph+vxohrrOBLH4sBYu2e9LSw34fPHtAYd9etNxF2X9v8BLHJASRMj7
7nG67j5j99zwvm05NoENY9jgTUUaOjpOOLsalVOMyMA8DQv7ozN7ZpPVKUqSoX3l
Ksr0B06pW/o7MN4TNvlcZMlI3zIwXiwsRAQPVvwKe4bz9ggzZtnBAVEazfCM1n5n
6T7k5qtIG+wYsVdAmZZluvA4ixPHnStQfmXblakh2yjUadmH8g5xupXWlNyzSVA3
WtX7DB9JzvFwoK5KZqmJi3+LyyuPLxRRdQWDCWYhBx8BIzOC3wjnaE1CwS4a6o7k
Hkq5AqsK3Q488Z9WO6I4k9liJ+w9nL2zWYtvCw0M9bFfWohyM9PJI9dw9gE+Nn1Z
H56/phBtOLefxIOm1ukg7yG1hyse6XXRylfcVJx/Ib/fnqgdQ0qVrSt2QGLSnP3U
7RyyJVshV0Z9JtVFOzQspVzraLgQDfQqsIVjN76wGZ64KojDQCEhSwN6sJFYjJoE
W69WeuOhK+oQ8Zq5LKlAHYS2F9jeWjtjhcF49KuQ1dZ2mzucUWIK3AV/eIIKiBAt
VC+0aIdow/8b9oXIgDd0JL3CF0eD9YFvfpxujPccyi25IG5N9/8o8OaeidcXQgKb
mKKJcUdcC+sKCsRUtZ9A6NhJSjDRuug+63V9uvpHJXO4eaPaLKJk+iO5Qtix/Cwf
Zz8UW/qWRxV69FfwvpDRKIy17Y6EpLfsAeLN06h+ikBshfUQjcmRSpJ+cCrUCnZD
1CQnQy4D/SPR+7i7/jAJGM2Z5jLIPG2dqpYGiFggSqOWldfUGCS3GWmv2dPMT5/2
mwgAakoTiljzVUW89qOPQXbCFIEcsbwYy2sqguOy81oemctPUnPYRKI1XeJOmhcS
C/Apx3gRM0+Gpn1Tfh4yddGr24JPSUPT9gXGDXD7hHqSbKCqVNhdUDAThggifBkn
VezuEsoS0E5fqxTpCm7xPJucxScaC0Wzfy5hj8axyrL9Wf243rPNT0m9AdaJqcjG
35k9Waia+/hwKqF005oWQI1tr3W4GN+Pl5k8v3a4Z+F4nJSfAfmMQZkxAvKpB/J1
U4ob9qq4kVvdGivfl3T3jL0I7ejEhwCgjHhZZkKDwCyDq5o9WgPUG6PCxt/RNdOx
xSCgo9z3/X3Y9iLz7yOP/L9XJ9f3ScI9BtzvFHAjqIxv+SDyYeFTBN1aNcCuINQe
zsP2qmWXJX+QUWo/zFgYsdEbRc+ZxKAn7VIxKeFKXh1qbcez09eHTCrxVWAkySbI
B/ptj3TUxDR/TI7UIcQ7rcerlNS5PC/cT2225Ktc8rjUYXK7sSjEp4fMK+M1j9le
RwiYNDPc5Rj3q1BtQBf8hCr2cm/V4cSbqP9dqJcMAwnmuzW2YRr2lR2XS8tGdJB6
MYm3E8BSK7yCITYgufpqedozexhfTIaEM3hPxFwW+gajvQeJcUNkTAbeDiRyBTXK
oNZ1bsg860uBhQmONbOJHVY5+KD2jtjv8+dG09PvsFO/w/wsaKoB71PeK115/Tqk
ZwrldL88gKejGrPE1HLi3SN97iXOvJF4/TKz9cNibFtHrwwve4Nmb52ratUwHw92
UJKplrldDfPS4+fN51uVc7uigJYaYuKctNr7XwVqDHDTRSU1Cb7SkaQBuJRvcaG+
tioy30QJjHh6pc4/T31ufZ3yNJDiWct0UCxH4OUeG0SmQtaz1MdC1nX3rrP2GaWr
vkftMaVGIhXHOdKUFvbnlO/I7OW6u6jmrREK6B1QejYZyfxXC05yHAwDnh59gPL3
cRB//xv8uTOfc6QgT3jTR3xSKrKrttE2usnzn4KWUTZ9/7InCT+wdpT0Eoqw9z5d
Hi22b6YE0G80QA0Tv8/02eE+9lmFofXxw5IGVapkzLxr92CJyy+ORXBfjJQKluRL
LzMH1dALilo//pW8HUItTcfIIYwpMyNV325cecorVScU7OXTBB1+zb7npAbZ1rx0
XYVrvCgRy5w30/Fvb3CGbUxVHa1vqVkuWF4e8+CZz1riUYkHtoCBH+GWXtnKHK/c
hFNlbai9GU9tD+CWv5Dyu/gv4NUrS6zksNmioS4AKcObzsrMHF1PsKlt3s2FedOa
mWWrg6rnI4fceuPdLEyHjHr1q6SyXcQcR9CAO/he4cvQC0MozcfvU3CVFjjT7lJK
tW4W2272D8Q9OfBlt/AgSjo5X1LcewdKRm+d6ulL5YxjdVegTM7aHvMO4rhzJ1bx
jgChU1xe/InVTRCq6DAHuJB1EVl5ykzTLiggehvUUvddZKiyjGHczv1PMFdNeA+g
icZZ1Bqx4wXNK7M7MCGSgw6kMHhG625YdnEdS0+5GZ8r31+5/PtEY/xMj2T6DJlC
rrbxBLTTKTpX0UR3lCa+NwHbNDWwL7qvhL+F6R7YPGV8YzF8FsUnMjKUFlGS38LR
91aG/8SgaH9uVcjFv2Abch5fZHld3byB6n5ze07gMuvFG3aap5BRCwuB+fsTRPLE
kzt3in4D+5C5P4gECS7A0sCNDGZeEf5tzG6bWifkuC5JJD/028ZVU834lf4muy0N
ZOita+qETtEwx1G9NsOqC5BXU/H1qRYQfHCHYLN7EkOlVFHctL37mRFs42mJ3lS1
GbNbb3QWeKmZZ5svyAgEDVnSx9k2OXiV5fjPG8aW+7YALwdaphV0Mo1JATs6cvet
Nl8g+4U9YbQH/hFOe+s3hc50SzoB26YiBiIkEefyhiC4qpSlePV+YxnNTdlr0vPN
8knvNGfPEIoDHrC7LiaJ0ZcpOv9pqafI71v51G4EzMGk0xnyHroniMur19nDUZXF
zzgjOUDTOei9tTXHGztTPSTFr/ywhO82GAJA/L6bp3b4eT0Lx6QeQoR5ubGJIgDZ
4EEg4rkHQr4t3oVf7PaketguThLFjQQY6Q9nWUlhbm0MgwZ73n+NOJXu0rbAl3mK
Nsqs8b95LNeAWe1bleBsi04pjoVW9pNWEKw4rAllWYoW7EQDKuoAsdXeABWpzvFZ
0jG6vXQAYUG8hdU+B2qHxzVAnDkqaCInXSY101PI3aUz82IOOAN6qTJwcp/D1fns
9jtvntyTMBUqtoDfqi2w2RaZyjvXGM2zDuDael9XvkPErqkw3jjlycGuza/t4cmC
xs1TQ/aSNSzhaSSwthM/l+JFyt5ryMQS/b2ixWotHgsKh1dePzO+rZzSj82a0NKR
ibY7ZyGRqhoZrIE6X83hszXzlKezpNEjyq2D8LSDtMIaowWNhjp2dH3j+VoIt+FT
FL2do0MwFu8Ar9bYiPn0lWHpAnxoQLouuGHQLlJJXrlYoot3rSD8x+OQ7k1+am/Y
vv0GHKjEH+C62jPVyOgvdyB5RRQihipEifjU/MSR4lELXB/UUclmefP++sVWixAy
sEJF9EhuAKvFdgvpiOqfe1yeshlZ2KYZLSKK+BpZXQisGkCO6X2bbwInBAxxcfTx
5deG+bSwBU2rJYefPU9+VpQKkZLaTpNpXgtX0iKM0ky0eEAd//Axj+TXwDcJsyBP
LGEjfgo+93Ylvwfq0XKdLj0K9cnCyZqxYZmtYM6MUw6+veXmAdHYs0gsnQ7M3Bs8
iwouKL4AY7y5jeC6QKabQ0vR/jI89nm5UfEu/1QqC/kr24aOa1uLNWu9NctUarhy
tUlEDYDA9mwqZwdFjIQVgW1XEuiKCYy5cD7e+8wKvGWcAd55C06tyPhGqnhUAnpE
Xx9D6hBYiG+hgsDPCaVD3EWDVW11z5WIQrXdUZqV8xhRu/0SRf9/wI9Socbu9J65
Vr5Qeu8RSDYLRFTrTy/4p+Ts6yHc5QlOglJCTElPGNq/soUWv83C6zOg17rsT4kg
dVczNLTXfitQwtDr2u2jcrqxlQSvDWMpUnIB6Xa7gGHdhPZJ/gUIDGequHMeDkD+
G37FdeV4OEEIiIhiyDjMYcwsNOh0WVQpHhsLRrpPKVu75wGcEyZ7XMj/DFgt9x2p
HX2u6sECkc8GemBrtcDIxWfh3ZdAea8p1tBdxqU3iz/bDIu9Pg4kZkETYNsrOWNA
duHdEnN3/56UeC1dn0RMgcSkGX+ykssrkSh1Paus8jw8suFuqOVCUKtYMFonzcjy
8OzrmTIzzzjecYwaWx0gRqr1d94Ml4A46g2JKq4rvDLMis8KiGq1s+soLZ/w1MXO
nmqZIZc8v9Wys6vUJN84V7+f7QO0RJvozN723eol7CokPsYq8kTgHKXPlaZtPYcR
zu0/k1+eJAcpb9xN9ClDLZegKwmw1OJnj8yF40sxUhwaz9fAD4HUuJFEtWuPeMSh
QDd4S+eY4vqJWcTMdiWN2AIpOU75ml/thB/loMx2CmWd8sn51GnwdfPE6zpaNQ6x
sYcSLs/oTIHDM2g3Wo/VGJDCv2crn3sibDTNoZE6fy6bTzip42rzKY9+asja1ZKE
d5duvlAntisoQpoq/CsWV8/p5JCg2hxhOB6rMG7ke4nxoTAm00am731Z5sEvXZax
neAXgzbmzeIFvX9MSEq52tMzsH/MWPQGi+FHsC6js6UZ4lqiUjNZSpmiSyQaHMyS
v7H+s1se3nO7lkjsFr+et8PAUAgxEBY9Fvt6Vhm+8AwjvlSzPCg+piboxHNnXO2h
z1odS3wIVuBaSfM48Z3JqxuKt/92aSUHNXG92is5tq2Ap9LkcVhJdJ1V5+qlroJP
rusG8Z84YbW0zPrvXnVQwFTuaQcgn+pvvyVRnUNnwr8/4ZWzq2rS6WVRFrKUx2sv
ko/EipQKVECUImwm7o6iMrCeG7WV7xOWxSSpGF9yYO+wHbfpM0mlrLsUYHIaJhP3
chLQxsqVQDiCZOXsCxgQL/TcM0MgJm9SWoSZH+bXHEM9Bhdl8b/VXfbrSeq8zqXG
mJIoBUMLAFmBUrn5s0jqRSbMxi9rl+RYPegWX42wUFvKxtsez7ZBTkpGpQVu9E92
pKldnZFYM7wKtyRKAxNOGE5rDBEVTKlSu5PrMh5f1vBI694hm3iqTsOXQ32bnx7/
dNiTvxw4NMGY5AYRml6k/N7nurMB5tVeT40IecLDxQz9bHQWtiRygIkmZKIaAwBk
37qEw3FBWQtGQtfVXF6XWlPNbe3Tg5koQA59lyUg5CNAYmJBdfI8T83g7Hg1BBiu
bh3qsq8kgT043ABKBZ9hSq5mWM/RuAp3vamr3H5OCYHcJ4F6IZq23cBsTqNb6xGD
QPk3LEy1zY5Ns5/0egWHpy8pMAtsHDdd3DTieLKEu+j0tj32j8oDbQG7YeLZLb5c
pN/7Zvato8fJeM9dQ0V+EDEo5+ry7y+SmR/NQTSNI8FCLVhe3xbNlo514VOGObXG
ZTha9YSGUoaBmEYLH6eogfpfSyzNegoj+PaPUwWD3FZTUsqQsdDmaHk9GTkk+Ouj
nRHDcn2TfWLmuv4Q5TYw7hmxzkGQcESJFyTuoZFfUHI7ogTry8P8kZV8wNxXuJZA
vKpWW+nhSfKLzcQYrRoyVMVNllfKpEb2ZcMP657P3J8mjtxOBTJOu4fpEdolKV+J
O/leLSg4RHIgRm2G5i8/QJXcULIg6HwiYxbPJHCLbsJ9MqhOrS0cNE+pCFPOnY82
eAWm6i4eojLjZuu5QWvZvoqrZD1WmKDxrWeuOW+arNuw2okrhPppnPMt/9J4fj+6
34dmmotL4kFWLiDRi+VzYorey20Cjea62JBMIlqj0fVXGyO64z6kx5V64ml5l0+L
IFJ/FEhtjR13xyP4tKjS64fOvyfrZAz24/AyGx6YUgirvV+VScPdnwm6av5yLweX
2SLq7aYz3E05zP7WgGcvgY1Zt88ACHUIgga3LnmWTx9SugxM5FZW/mGaggtSC2GE
crPAre2c5b3f0KHhaKZDq0/ltJx3H3BJ8BFi4IlH4doyPDex2VlWsWF5DfIFtdRT
BP9rH1ZpxQyY4thtAqvcAzp1ARqI1qCkb/fuOS7ZDlRl3eOc9CKpZ28I5BdOJYsf
xYi+i6LndvlXanRfWYoYCjgRBj2GS08+z4nVcWgjyycv20MrFxgdEtyLh4r4PnFi
AeLkJU5s+XVcMBSeOLdCmmee3luGu/n5iYQ1TDpbvHVmkDopnJMpJ+Z7LoCHQFCN
fD5PvoNAfdwwDyGsW0AyB7NR9+yS28zuis/KBDd5yoDqnJTL10ZesREWpbucupiB
PUDTC7mrcuVs56RYg9PJpPgh/g8tFaU3T5KVnorIrenxQWXxm5czYISx1LmVOF4l
qQqYEAQL2T4QfY/iP5ShX2wDs6sk4OvQVRT3GSZpLhyiPsPWV8xKICcEJzpuSVoD
5AckRqGW7o+31ikfROTz9aDWf4Tm9FgvEGhPhBEmUKfVDSQsw5qs0U07UbATinjc
UFdhmMJl08wMDg+RdwUJ+tCEmFRkeu41uIP1XosxsxVmosQDVYGUbxd+31yEd43D
QVFNtRFJFC2VnQlNJbXUVs6NNAJhW3mj7rkUjLG0CWTjXIsX7Q6BLCdZcJQxmt43
RnE/MSKeFackZRqHIjA9HZg+3V5xQMkRhHGdoAP7828tmhvJhAzXMEOth8Qko2Pc
M49husI1486EXVHgv5rjZXv2BmE9NNb+oLO4Hyv8ZO/gJ0f0KCwgK1z8uf93ot3s
XoUAolqex2bdXBfx/sZrnBsEghR4/txJyAPZL1C1hTUykjtG+legs/qiCNmidEp/
wwlf/smY/Uy0m+eMn5SR7FZYKxUU+AiRH/5y6jqYcB26d+8PlHiWFiSlPfJFiyuy
H+lmQ1+5WJJnXGwmDudRMAF95dFbuMs1dXbTS2OeEucEe+inr1olsUaQ/ubHFkhJ
jjv0P/snTm2JstnB4v42OJodBJ4JbHu/RRwE12eN8b0tHHwEsZRPX4Apo/uYXs+6
bh22oyy0gou+jb5HVyLgTa5IS+tR6RlRYei+mXyZfd7Hcdp9q/6j1Ckdc+QSMdWw
CynwBr7LsvGTbwTqeZ1J4vGVOnPURTrI9w3iR53MARwbcW7cx0pBxvdOKl4Ou5xh
pwOEa5ZVdjCM5ka2Kw4gY2B6BogLJXcfuxQEkUf7tB/Yf5TKyEfkgZEJ10t77oTc
4sS0nOchiPSZETjj+YCYOB4rgVxWJfH+Dv2Oi+nYRp5CAUNTYCDfF2OD5Xfeylaj
U6feTNgkBKccJRnGZ04FR0sY+fetoAY2bWmnFq6wNRMDxxo81DVoRop43iao885R
BpvT6FgehLzg7rPcIFlO6AGdN4KZiph8djKlcwTVtqdLFSJgva/Z8VJZMe0eVEAz
oOhlbkQ12DQxmuh0MEAvZc4El4SNiL/KiPcInNyhq2Des2PZNlKVyCAnsGvtxiY3
6n444CB13D01QNvRPU0fOCJ8bPKqozpPDOPPi8j0B7hfSvBDSPKcovWtVjQVbYm4
8z2svIJlQ8XYPD2md8lMftsNEiOWhrunttIKnBvgEWLbYVR/miiGNh9KROvN5EZd
qRLeTlIko74zAvc5zj8MqwUzda1yqB4mgWkPVaQu2D8KTaSNjhOSXINkJV+giHd9
ubUdY7wZzL8uxXg8rFBiIYyvU/ueSSjdz+mE0uDPKZENeMN5RlhjpX+1f3PRwqcL
wIa8JCK9WBegbWv+xOjD0qwaW3Vose60Gropip2hvyfIYySDlCzkgBHTy8Tm9BOY
8dKZF1HYrggS0hSAGjZL0LXILf9xs4AggpmP5wHk0Dk/z661s3G2gj9LCrch50HO
w4hyaqxbpDWTN1gkoGTTtUo/niu2PPDIuIzlQWpmF9yV7w6ykZfxCpmeNtsB4LAe
E3qvONKvESqmZCLGE9oQ20zVhNZgehhsHWbXWfaWckXzM64Mbm5HronA4vULM+qB
SFaWXwuCRhHMfgb3UkIBpMoMTxyzMWIvZpNIHzOtF4fn2htSPxGfsjTO2ksrKWL3
DsER6PVESC+oHCukwAGGeKd3Cf+N6eh92KV4n7LFfqrvMC0RENKfnI7ydNDNcJte
5tblduHBOop6lbYCeRBqXSgEcJw0k+nHMDv8MZZAfnYG0O3wej2rBNW0B95VbrdY
VSuLBmqu9uDpfGyUyRQhimxGpD0mxxv3aIHJOtx+Z4YrAsUGvpMSaKCHydyDNRo5
Q0dfmYNSEiPI7OOH//e5J11Oa6WAJAVmUlLSbYlCtwqRCxIH7yk7VbfKNAxQBOee
AqQK8CeRU76hTWVbd+QX5j4u6dC2T5lv4/bJXy6nXByR3/7ycGB2OcHOhVtNW27b
YdtsyCe6n5briYXlm09ugbZb1iyHJB7nDeT8+1n5mFW04rZzOnL4fmynb/BIGcM3
IXyQaozQwHGBelqewHqQLroMS+Us3QF3sZTUUosak12B9Of6vDhfUs9QRZ55S/Y3
a8fZIoYT+zTfDYXTgZi29DRAhWgPmszFv3rWy6fStKoJbCENsSoR75QtvDTHQBVY
ToBw5L7KPcZ/ufnLn1EyNBdc2iEO/JqUihXgxf23cBSA4MNYJD+b7abezRgVVAxA
FHUEacbhfBnkmmeBE1+cKNlooWsT4QUS8AMzkv6RvWjqyxRSJOA4/doLNClTwvtA
X06TGzk15Vgbhchz1qecldIQ/km/pS8RkxEUK6tEaKFS4g/yL01QOcuysT3/sqTv
wgRDozrShTheMmD7j4afmPaM311jAu5GBZuzoOHMHfPJIQP8+IBIk9rRgpfaiOFa
bJk0d6JBUqU4C/47hMFkA+IlmifUrzuCjaRW9gALERJ65Qy+ye48ZzhYyHFi4OAB
qftoyH+TXFSBdkdNxzcX+sGYZfUas5gBOJ4KSn3K7FCGKFb5TgEUTimLbl2SABvj
xiHDHp0M7//ucEgNXLLPUZ3pwclpFtTy48u8tkQtr7LAVlgxRxdv4GbLoE0GhYyV
F6DPZlMwtFPKWC91g/pM7WTVUxPavEtn3tMWQ28MaxaPqjsxLERqFvSkKe3dzZPe
7aBDbYA+OuWZxd1ULZXq8kI7elcXkTTXvanZQpkJpSdDqLO8busdPlhPTybFxh69
/jvqje0nh1WI7DHJlC9FP1B6gFRgxh2Bdv6dqrhCCfXGdgox/1m/C+kPeEpgnX8h
i2DZY3u5kxNyMxg/59a0jpG3uta12saYsgJBmGhFdCz6oO6z3rT3vx4masdS9ZV+
lJH0grc8+AFB+V3hbf+5T8wAkFX+wNZLob44Cz2i0e7EVFUdZa7Mulnj8DUnpW8Y
mmCWTXyEVHB1aQlhFmHtKoQqTY0LxBYBWqQzM0qdWBOEh6wJ4kMF8inOJGjD6PaK
jvQXnkMAeALmrPmZ/JqJhmCPTMo4t0RuqRzFZSuVSiAuykaT2BTLeiP/AVKrqt8U
BuygZ7o0mpRKKrqDSNU3PXxlp8894iuRxdBHhpv0k/SkJ2LJncN0kGXtWoyS85cA
nxihYZVBtChA5hpu0Wq08twmgMlOL4eIKkPRAoMB2jORNr5WZrNl2YmSXdFGz7xy
rFbuvSNHhrf0GQmnQKbYios7Ca25Ee/MpCRbCFUEsdUpiCtVZ8ugJ662j52TjTOt
yYlFuGDeBj2dz4oT8WnnpJyZZup8mCY0W778Hb8weB/MSp8Kj+qTQrnJ0KcTKjx8
Sp0z81tARCvNgzAoCo/TuR/9fZ8BFMnhUDOPKfqywvb2vVCS0QRHXVT/SBX4OAnb
tsFuceeA/Wtpgh2pop1/yIEWnZX3SuI7P+bZNri6ukHWkBLKYdVgQAjhyyN8u/43
aH2eevDgB2HR0oPRgVdYOI/yiRBKIpZLvuxJku81Kc2Q1v5vfzaVYyDKh4KK1pnD
YQeq2DKrl9mGTcQ32hHlyAN0Y4GYRmBiwjxYWwbCJ36NOgoXz26Eu7cQRCyfvsrY
nRlzgv2MfiMtqF3ifxjHPJW1Y1CO0Sa8xpItGkGYoGNDDr6ETGiZtLQcmDYt/v9q
7ZL+VmWANJdYEE2VdJAfmtQgmjKi8eC7BhSahqTW2jY9iBpZUWEVGqyfpddj7djK
4J3SEWJItQ4ZTqI86aATFFm9yW+NVc54e+2TgzM7UC8itJeWp7bWdpXmLotcq5lx
hwQCnAIBLIRQM5RPytPmSwr2QANSVtQmSrBfPbvUUuB7A7L73qJl9QSLDg/uVp+H
+hwPRCxLSe6IejM1Vdyk/4pIluQo4DJJ+tGid72NP2fghvZrDGl+oA0kXEl67GIe
J4CwCNuerTuDXjpqVvNCNw/5NC4eKEt3dSz1TzqudgIo8+qn4ixAmkx8TEPFGp+/
oMjIds1girCA6SpWYHH48oql6DFkc9JWdJAI0motJdjxGw157ADZw5pP291sF3gw
VQFhcyxL2vYHZzX8Hvtprl/UD3g9gsV9vnn80/PQzfULv05Ee0itgBAGQYx88Tq1
ssWjictBYBHbRQ1b/5PvuOxesIfAOLRvrNVpg/atG3iiMtkUi9S6dgsMrlwV2iCD
O/fHweGsut3vS/wnTTEZn47paSl3MCFhafqFhu8U1dsS1yiFSdawsHMzQlNhHeTh
S/gEnTpQu8rRK5EAT7hDa5cas2vZWyHUAZskmIYVMdmWQwT/47bXuHSXSNRrkVZp
tbi2szkhaB9TaUHn40aVIiB2g2PL0zeR3+ChWeEcVdH3aWONlYjD8Aoio0vYmiXU
Yhs4tSLMsJP5D2PmEU+ferHr8kR6bq9cmEzlxKnY6pI6C5RKW5rHpeXcO19eIww8
CJeEcAiiVc3DGNPpQz3zzOGSJJdGq/XxJy7xFmnz4lysE56SH4SzJdNEldmhJBjK
hE/A5HZpeYBa/cpE9LIQDLNwTKpLOa8Qv13VWtRNS/W+TXXNPc2n1WueVulH/nx1
cWrWD4gF1CfXRyWzxIirGFEQKE7rm+pooAQX74HYytvA5Bu8irePPY9PQFMt8//a
twD/Ae6vvGKiJRD8pK3RBnsaPPgXNm8jYN7yAkMJaDuiMLvoCBplL+kjCPAv0r6F
EEp0TgSPMP4ZYFvde5fTBZ2Wx4O4RYR0onBAh/fBLCs+RkKbawawN6dob+/Qjytf
6uWEQDLwQAX18z1k9fC6LmIT3JQo3T/7Gj5i8P6QJTFhFCvjqt3RBbhPrjX2dbLd
zKefriFDoueQ0hAoOpRuwtXLQ0Xmr+Vm/a98Os0zVX1iUWzL6/sPwWj5FocoZwT1
uKUJU7yRqIXqpE9uk3+5JYruGHImw6I5O429qe0sUNHBAxFTAG7wqMYpfcsNf9WD
kVRGvZjeeeB05Or37o9dF8FzNVNBpFiZ2JJdgnZhOf8O9v51mm2HK6Zqx/ZIwSlN
ppj6/W8m0lsLkcNAZwjhHDyb6CwVmljjgzYZwsYO2D8vXzSwsHWWZKw4KNUKr/v/
QX5J+0UiTnQ6HhhyFNYajsSwynosWPrxmmJIZcBw0AiqP7H31S2DkwfFwe/Wynbp
veCYU5v1fN35HG9HF/LzGaH5y2PvOyMlWbKUCnpedX0YN3NcSXm+S2wexmVDai6K
UwY9hvv7jGGpRjTmymNsXMQjLqDbYk4sNFT2Dj4JL37Y0qVzERRj4+SFFUfYZrpB
T0l2DC00P0r6rrCV4OjzIc/VeBOXmV8wdNBGNh59HNbWNNOqeCboknDaFX4O5Bxn
4eGOnFv7zxgbahmVIBhUjjMt148RxYZ1Wv6H6RmHgzpxGtXVbQP8yHs4ixqp6Kkq
WTyTs3eagbjv6SoMn4jhTCNfQlB3ZPgmoTcAUNChpD7emiFDp29HpSTrikKigCS6
n3bMePflGkVis1WwEJMlszg51O03T8SBp2ZoPEvL3qS0BvlMO8gKOkCBuW93pwHt
76XEyq07o6xwk4GqqnvZz2Es4uZFc5bS5uSDdGLHVOYZnce+9+BAqB8DUfHMCaZF
SDgR8Y3BQBBm24u/gXRcslf8kLH58cACBawTHFZfW1hZYSLe/sDprGPVt/22wUrZ
oI3+Eux5qRrPu9hVtZUGwbqSJyMm/YaMRlTtXLARg6Daj2crb9YhqxE+FqMTUrtQ
q5Rd8xUgULNgO9XYJlBdUb6yTLcSOLWVt53OO2UVsWQP/Jotfy9V2+ngpQ+jkqHO
O5TZBljOkTOL8B9pBof7LbmacaQIj/i+Sp++9SVaFzaUXjajshrilgqj7TdMYT1I
wgz4rSRO22Ds5O7vU6i2Ffvn098ECTKFZdIbmO1yGKNA0o82QLEr8QaTPIoMOqd8
9FhgAu02U3NCyKlbQWiejeQjXoCaBWtuyH3/qFSRQbVSOpPm9vqOmamPk/MjIKOK
0W4RasQ4wF3hWub9XWuAVmQgUkJjZN5BsUxv5chpkleDZ89bejSkZCQ3fD+Kmi63
sdFKK9BDkM9eEac4xPaFECV8Hw7Nx21CynNOGa7Fvl/79WilkksWXWx//m5UJxl8
7FeVlWM8WHidiczKDggqeVp9+D/o1s/YQynr9C3UqKOZPg3mKMKZG7umwR2Vg/fK
UlbeiLrqLkfIv0OpMxutnvDelxuRcyJCjEg94Sr8VRfeMEqt+CS6JAHkR9fdJ9o4
d+6/kMbGjCTLAWzeoq/uDLw5+db7ESm4Kr+zhu6gMqKMhd5KDlXQwM+E7rdp3AcT
cHjMI5pIDyKA0JEsyLGCnv9HGLHuhjKtpv/OMxjtXaQUdCsSFnh96aYEC2Zl9j5D
yGCGhiw6xtlhkVcYQelTHXzE3sSwy1DzfuYyj1VaCUphTj50zP8fjKmrkD4Wexr0
KGhiSQlR/NvDQEOJDB/H/VkLbn+twy6u4JzlE8jcvR8JItf2q0x8vu1+PiANcMrp
3v7X1tAijS3yKzFposJumkBzoq1WSEYy2e2sTmxCah/6mkgHLaT5mHk+hMtmNZ3S
w0hRP4xW3N78yXIl8ftM0wRhAf/IZ8RH5MKGtUz3XQy/6wfCd0bzVGfLIM6DtSK+
iqNJbK6SW67hln5Jua2FLRkEyAc4Lio6G3ddnckymGEc6PCp72nfvVsje53p6b1A
8/k6vvCbD5h826RvsJRFHMGyWbnAJNMoLAlKK8zBOPaQvmDKU449WJfC95OhqXJd
wTbC1qndzwwSxIJLFuyuU5YF+fwtRUpzbMrQtPhlbXu4QMDRz41lzTy5wzCkhGdf
UO6NAtaKb7oF5TREmvlEZldS2pf4bo1vld0f4FzKtdXYnD5jIFfq9YqJvDkWyFtj
fugIQvixUtI8YI8ZJmmsWk2ewncWzKttGcUQHDek/4Ys297DTsRIYVX1zZi4NvuJ
+dVM75UxAlqegVceZcN5Kr4zBPRRmEI5O0ttCTXcjpKauGEsTrMh3MwYZSTX0rje
mMSkEKUzXzPLyK0za9ngJX4/EtlAMApRTzNCTwUytSVI6dceqS/qLNg0MqHcaJCu
a+p2K+YQIxOwricmDL2PXR1pw1Do8e4D07481dE3khk2jLZgUTIrbe0xYf1D0o+M
oS/cNHOiFA5/e2CkYVyqmp46U3RiH0gzcuu7DLHjbpYp5SVRQFquj4BuJSyl2K1A
atgbM7sojQsGS2Gh1ODss8QR0yOSnjQSHAvaed6nT8hdE8Fwe7x8khETNXC20h09
b6uAak2vORM17rClJJDH2M6vBiXqhGD542KQJtF9bvrHtIs9fZ0jIA6pMJTSpyqb
QlWX/ExW9UZ23FfNV/bQJ/orIWoC1c0pcBPJZExby7hRa6dB422XE4juwTQkBYds
GBmpbrIoS9ru7pk3d4X69qFLMLKn573+OVvMHgXiaypYXujz6h4nQtVatNidCVr3
xLchQH2UzJGtmghyQcV29ddvVlq+Hp+IvSfQUPSorEzo6JAlqvZQ/yeuef4Hsx6r
RC+LfXibCaEjnmVXmRleOfSo2o2KUBUd8eB7C3CTBZuWXsldnes8Itp4BiUvL6KK
aQvy306tJEVim0ievoBoL672V6fmBpE0JgHivY2QmhoYOt1+baRIWQHUam72oWq8
Qvvd7VeysFUf5mHeRCHgLgC5VA5Uztulw6eaCw7VsywWnojZOHlM28yDdmpdE07m
eNT7my7N5wLYNmkkInxs2JfA+d0G0seWlSrmtfJIaAl4x/w32WpKkt9WiAs+bkV7
jlfV0ERKXCBot35d8SoX7ScT3Zji0a007wg7aCpDK/W4vRcshfyiE0ran8NnzGZo
JuyQDk6fcjcJHn+wHAU5upi3TCqqKYq3rJgFH64ymZK33RrJsa4pG+xmQg+S/0pF
d5ppKP+lyfvPuhO52ST2gty5qDl4hglZsyrafCt/3HwkMe2apHBsCyYIY1JdRlkO
jSNWM3lxMfZUSWQLt9ZRd1FJxsBjqT1YIBlAO+z0ZFlP/8Dndb+YPBkJfbWlWokp
g6Kcq9GPyC2E/JaeXwyaXMPbUzyJ4VmNgV1dZI3kWmaNPta0pI5n4EHcVV8XMQah
aoxKcPFwmgBkI3uLAVpSeGtr1KrEtlfUKZELuSRIP0CcIs65l5NdcsBVDpl/qf0g
zmV5ugZOmgH1GlwQfIaIuTvT7/TTDVKCd/1v5zQIYm2uFnsT7I7caTE69UF2Thap
j5VmNak2esleyWqU2D7N1gYBWMNIvzawZskPV/EVid9jAk45mPCL1BX1vaFRHxb6
55YX2ijBOGpqI4fu0uXIXOTsdRj2Ib6gAqGnjuaetxH5+vL6UuYB5af8tXUUZhmB
OvcBz0hpBwhkU56lfIyPELmzVB0y8owua96mJ64qd7Ia9tyhLSpuKtUtzzR2Fr6P
2hgTFExSMnTzGZ0TO8nASUJ71MFtbaJA90DIbc7BGsnoFrFNwKnbP5FUGuSfekFm
S7cpA4YgPnvCUuQIMolq0dWhsEDLMWbpXJP+9ukygR5rHkFDvWfsd7yeCCAJS2so
AR1f4T72gR2X7RA/BI8QNjxWIZB4V9wzAOL0ny4g25TYt0fhFnE4DlPpQE6cktAV
aYBEA63sMbHQBvx6qBXX3jPTNa5C1F7k72WkY0IVM38ouBrzxtvGTXKosvX00oWv
8dctmpUmPRdXCLDJkGJu5CZhQdH+Tfn7/jd+kEvee7DXCCqOM3TUvd2RBbqHYSwb
ZkETmU7Xfl3eql9W9YRYDmq5YrScCW2fhfrUgN/KdQfC/ruQpOF47YFDx6XJ6wAz
hrzMk99+9TO01Q+CRgdnfuGSWkIXZceGTBh6nH5lQgXp7KiJdsdZnDX4Fqj69vvb
BuKNGBlsU88AZVbwr6KkuCIcvbJWi4d/qQa1hqLvBYoqD/DpQHJmr4rrnrGg8iq5
6stdPlvBOfnTECy84ngVCWJpR2q89INfsrBrd/7kv1cGQ2ejwrV9NBlCIedIuMqQ
cSKeqRugusvYnY9E8BHLcKsakB9/x9BcMIhZbUFsWZvhccGLa151BkF7YXA3pQ3h
CvUWr6VezZs9A5oZYdo+ZeMZIyTgLykKsvKajXfHHUcoQqpgNvZHcgeqAVE8AToZ
RrmrZ86dD8gpq6abSM+gv8ohOXjINQAtQhBCjDQuH+5DIQsk/ikLKZGAabLHYD5Q
Ir37pQNJMl9Watd59lRMc41JUpVqNUrKdrFujR3LchQsmkHwzWoOXnmNyZfc6VEH
Ekv0XgfzQeD/jxuvkvEmqWkFWVrm7R86rlICLfF/Wpz0gwZLKw7sCWWlQero4I10
KP3zn75PrOP5+m+jI4EjzG/aPFuWD2NjHoL2pfZjdomhTKyRqwZQ+dPyWwD15Esu
Rcz9hVUGPSe4TSKhz/Ej3y+WnChhldwOmnXq9fSB/9VCAzQc1S3ZuFeY/jn+IN1Q
vYx+NZbh7L45h9RtNhL0O3Nvgk/6WJomyAy6Oh8zah3dvzVsfkb+VdrR5z0TDRjc
n0Jnnx+WM2+EN7/VYNIW4rUssjp5+xufHL9+5NGOSzNMYuX0B0HozLKKltZqhByN
rI/BtWndmQdQM3cElVd4CGmwjOfpxMh6izDRz0qaDym39C7RnvSO/I2ovUbdIVjJ
G+uGVK1CII+potyUsLZMRLYTHd4RBZczlI1gZIdp7ECNYDEDYc6OxD0nvYFdw/zZ
283D3Ve9JwsL+YpC4AFsthFISO4OqwVis6ND96e5BlT4WrAouI5gGYZWEmjbhoYb
ngaxLBjTqkERsH0JFcjWlzVmZ5AGgzdH/i482AeuzUZqvTiGP4FjlEp7n3NOPGLh
ZIzRcUVuD6XHboUO8/gF8MXH8gTkJAxKfU6HeKU+nC6nyL0G5MBgktRpfI1qsf6y
XarN3UP/MwGMfDPDA4TpeK3g7cM1fKWikNO3ER0n1srtO59nfVppNWCE9TqsoFe0
DinI+c28zhdTPH7ceGqm1qtYiC644I4Rfig2QcFV2TonD/m+H9PiNiQ/QHHFfTSD
bfI5kWQ0gPyzeeoiqdjC8410tDPCGqRTVCAXii01VwLfc0lQ4PedAE1ls4z78FH5
ebbtCQh6ckK7NOqivnH5iZojWYjw+y55S+BOdEwdoojT1xCVAyHl0M2D9zZqoI3i
XnfFrpFgrt6pd5tG/uyoTqiAocbxc/pRHbZ9lsdx7IVqh1oCE46u92sS2X1zT3YD
DUcQMbebbmxIPUgTSE9V6NpPraqUbScKr8bx12BNZkk34kRrBA79QQrbz+0P5ZhM
92DWiFXYjQ7RoDkFvTvkowRAU33qvfLMlf+LGIFeU+R6BfzkzY/0ikWhSfUrtBRE
JrrheAwvtx/WHY3q6jsOmv323RE37JYkBU64HFxCs+aAM0w6WXk8PvVgPPeaGnVw
PSCWC7dzJ24f3njC5h2+Uk2Wua/Ir1snJ35Zg0waUwiWqnxRTVETgrWKSjI+LBhA
yUTEjrhW6Tyqa7Mr5BREmKbL0txay1C3NR4mN6xJicnyuAQ2vUS8xyIqCoAKEf72
ugJ0pc0onJt2JDeh0kEHBpW/EbGGcyyBZl8/R2RphIb2TIc8xtsE708O0e3xo9ww
5VmHEW0cODl/gTgSHUFsXOF7XR+xHAfJhGiUDBwmvI+2yuS3ppiocXE2AD3YeziI
UBEUj0AXYH2M/a5ULM840Eb5pyj3GjiGXXK3XM+FpoNfc7u3NkzS6WHYvadiPXUL
Ka/B/o52MLkMob82iLzwRNUBp9GDkdjuiG1lJo8//Y1NVv5tC03AlQAPO1EAfRuk
aDHAvTv6AoVpdvvlwelH6UuRkDnB5cSWoNo1NE0UcahuhSH/xCMRz4fK3vj5i/ln
yfgeGWtUkvPm84ofhdFytOxGn6lx6jctcLaFOiiJtMIyfmI5Ljaja1q9KHxJEtKJ
ZDYzZ26zMtbA8yECum+i2b+/HhsvGTNLPSCPAAQ0HBS3YRCptSi+ScHz9okTbaip
p6m+Q1Atm/qcWxBuaeSpc0vHfgsVvf5qVdA2tqBgfx3zy7NVvi1sBiGh9GncFu3b
ELXufnzZwSpfXtpE0i+pseC8jZ8x5E9hVP+u7N1BxwmZNOpnpYiDKnlP/8i/4791
UPrLlm5NsOsB2qZ99dP/RFpSGPKoFib7NFxIuPSxonrog1RTFnrjrExx6R/FPXys
rLSMaHxqMzq4jB6ZW6DCE+kAvTyjPa8yZHHs+pr0X6KmMSDJLpPf6ZFuvu1Vgbvw
2JD5gfHpLRL426mfz4B1fNKap0wT2wSRIoHCyQwnfxbUFawiLs8nqkEf4acLIwd3
e2E+UhKFul7BFcn3atb11sCansILd3sSa228Ehd7fcZQo4Mr0YFlL1A9xTQFGp0Z
ZUJkizzRtJC0etbAL+MRZNkpF+SsYE/bEbNg61P09v8fc01E3d+xOuNuKfGVrtAO
O+U3b/44zEXSeuKQ+Glj7YCOR7VK8AQkgIXtB039Xd7hT0BmV67Y2awZB8qMseC6
qx9uz00Q/dq6Zc3ofv/W8CuPQjZZ6y3uESxwQdxTHo2CNzRf/y+jHr0PMhysTLGV
2fBukFKt1VjAJPf033kHeS2Geh/dPz6GUBaHSNcxrR/ZsU4X9d4g86opBhTQpacF
nhNkxB2zGOuyThEwQi1uTjirCaBbHi9EBWIqr7Syd39Ygj/2FEcLAwgroRRERRDy
A5y2nN/1PrrBh1vL7bdeDnfjn/rtj78hMV1wzBSywRjvy9EElzC6cQAqa2nYStDa
Bqxn50qqcCU1GVGG4YcX+3djaOssmy2kCTPFkFBX1CbwXxRe+jRMNDv8qfj/Xvz9
ywJqH1aXpkbi6sYOMDCwsLyBZhx7h3fWEfLhOnIN7d2gDSJCzr8zRbcPHBuFZ8yv
mvNRm/iWu+LRvK84TXRVTz66J+xqXr46nuszQvbaX7MHTeg1PgaNE39p7ukg4Eqj
lLy5ljoAwJxj5D+zrccl3liv/wPrasG8Nrq10zP/oAueuRKudWSz2noFq/fh0NcU
92P5erVHW02a5RBK+X+WZNNSZN92WD2VZtBRAivzW6Mu3Itrt973VMhyC1aeWkJh
cTmEEb09+c3fHsiNp41ZqQSXrKVaU2+gWmkDqOIjLL1sUguD9tsPEoLUKaXPQzqh
xIgefc0QwxTEDwKEx6J/mFbK9j9wxM4lpk1Kb/+KIFurtU0BpWDZX4x2FUFZZ/pT
zScYdnL5GaBDrbMSwQfTYSTH9Ootens0aqUAaAbSLUhSm7OKXl8Kl2OkZNiuNRkU
rclxZjoCOTOpA4PsYP9lTOXqj35HkKBM8KfjgRQqreQFetEMUg9+QtV8eE6zRzZw
njp1HFGLKHVrN6X1wfN4H4BzEsmcuhpLU7j/tRuDyeay5lLdPSCOv4wNaXb3MPye
7P+5JIktpE+he/jgIQ2pJYkKOJOF+gY9rTw1CYuRZZ5Ge/p+hHVN7hnu7eTKN8rF
H/BlZtL+UacqxdShniVRmGv2RYMTGukhTjhPTxb3IlP6oKu0hqx5ISLLciaezvI8
4Nyv2ZivXrV6Pp9OQCsnxhciZsTlS2XDhMfzVBtbWkZ/tsYjZHsUratYtqB7TUOK
68zrKyVONhlGtyhzK22jzeElsMBPQlYd7eiiAwFUo0sbvpGnxphGdgiw7e6jVTfN
BKKSVcChDshvUzM52+w/GRMmMj20sNq9U2glqJ2gtB0jrVnGcEC8Y8YcrzAYlITC
qtT0Y4ObEVjnBY9Hjf2uC3W+wlrGeqmbjEiL+9IepyyU6Z5MY7rdVEqpSTxamqbX
J3I1P7Q6ono/r9MVrkpMfdjm/JSEBEPq+eymZkC2gzr2zxUeAFNCSoojxJCQKeL7
D+ExCEtpc9Qt4hDqKG1nt6PA/TwIi+AXm/PWy9w2fwWLR1P9mmfJyd6wX+wI2qdO
t6DQkK9R52RpKzG+3sZD/dtYc/8na/su3zN/pxOl0AjJM5BkfEwts/7o90HAETIJ
2f6O5fhOk/lVOBN8y4ZZXll85cmokqOa1RC+DiscE1dPsNwk/nUEVOiiOrAoDiJK
f6fvr/Ybbr9zwfpMP9dt6LndCp2AC5rHfk0pXpiw1Eh63SnRGSA19fel/XmPjawk
0YRDCE1VEUhSUsWiqiD/ZBHThZ0QnY/fFYlb/vCumJ2QVrQjMnlzQkh/BPSoLvC3
LVcNmYfRRCBOTEj324rvMKzpAXGPWhL5Ge3Vl35eRk4iQzVlUjrO9YsJaZcqCCou
PGj8bzI5Bsg5yrcBne9O+pGgmIgMYECT6ZEmAielsWwWnOvT2srgug1p2wPvzB7/
2DjE7Rrgc8COwHh3fIeVMKNC6Nj7KeHktPTJ3b6zU8cy/sk4++Dzje+uzCt3lsSD
pii+5lMWYBUx8JvpZjFoN6HjSjto9PMNr6KK5r0VAgOojfC/5iU+fhuOS3OGf5A2
GFlui1vPGZ5l7qirBihx9A0B+W/3JZfvXaEQ6evNMgPs3R8WGei6G/Ns+WUXrFCU
GZNJxpVjnSvU+wxY9wQz3KA/kOZALPkzYETN8WMlqDYUR77jDZqBsen4iLF2Cctl
sFZqJJQD0TaGGjeasdNuB9P1X+IAN8sh5vbzUhX6KA18HcXoK5LSQVvSl3XUb1Tf
Nc5RS0NBdMgTF2h/ppC2H6/c0aOAOTmxZFLPDNP8ZR2rGiuY+jqRz7GKRn3rKxad
x8gQbuctMEFSyqgyGXPG95zTpvXPI/zsdQszdcFvdu67Ntuo1O9I16/yzUGLcdqM
bCoCajUPhJQ6viZbLCQZZ2ufpeuNsv2MfQXgqIothEQJEK+OozkzsnfAsZI5wvY3
IVDbecCGjrpXKwVbK7kVZZiyP0TSy8T1fc59cvrWUVkCOm9jC7zptF9HLaQ1OXUP
ThAP9wICHyv8b+KqJzQQ0YBb5g8QKUastX1PTgYqQBAGw7hEYR/LOYXbEhC6vsk9
0zfNz5ITZwpqe9mq/ZywmC3XSH5fY3SrLeuYaT0o3gCMi6s52f9aVkLRoeBDReDN
yo1JC6EsoCQ0uYwgr7+pyxggjikC15xJVPZLLzzN6MG6UGLdbxl+eOj0gnmgpFCg
lTH/OE9CXv1bs+PUgYtR9yVoMpNIJ7u0sz7cWCJsjtTWqoBErjD4lYDgl6plpsgL
Gc7vKS/vOE29jtWsr+e1V/A7WtDEXQGvXHQXDhpQeb3wd/7PcAHrXGr+CeZQhW6o
2TcKxCYOkop1ZfOKSGGcjJIAFodqzlPyaha3+z/TI5aHnk98KQLkzwgg04daxps1
JI+crY1cMvEjf/OfnADdjcT8InYdIZspsiIo5aE+qsCjWWP0XkjU7VhcgnZejENC
tnUdIKNfOasQnNvhY1HzAOpYdWeGMykPP3S5v3hhZMjqHbotHZjp2i9/d4bAAP5t
iiUVP0RUJN5a2zypObkEwZbKXaA5ytSwUCK825dHMa/bHJKyP2KPeMHxD9wl5xqd
1LxnHwQeRViLK8U8tHBR4gYhah7IOKJ5N5oM3yzW9U3yiqrKRgevTj+tbga2aIC6
xC38bed/ISleg35k3dr9El0+lXeKa5BSpkJvHnYdpN47KSUVjwWfC61O07k0RECu
73YaG6M29qAbgSRS9o3WYVP15C75nm1SO/tQVOBtOPmcYLjecQXSd6+aQ+Jvjdti
6xK5OXln+T1YfpB8pAgQx9eXD5nWR6q96HUbfV6CGverRDG+vuUhZDfMqiCLZxzM
ry1+Ki5VA2kGB7qbCuob2O0Sm1Il3ru/aRWVGtf4kwGXl0qSHGXMZgvQWRtOU7hl
LwD3cRM1ljx0PO+/m7fyRI60PTVmsp4w9+NZuX7R7tdhGIHAATNUYAQJTikbrFnV
pMQ8l1YiDiBYTEx7fgVNFObSYj1bMHPyiCX8YXa5E6cF5tPaf3yN+IImEJHdNWY1
uX9ypiD+adGhIBz00GiBxReZrO9rzxUkiUFyl1yx6foZLfr7AulCpWnRi8PuPn10
xq/3/pOEGwfT7UHsA48QLRTd5ior3k1WDSMoTPV0eCgdV1fp6mQD/5kIRGYhEfrV
K4aJ5Y4r2ctZbFhbAlRt98USYv+jmc/10SQ0iKEWHQUD+h+50WGUkATmBMnzkfoo
OWPEiWQAIXKlMOmVOM6OCp8g6hYjR3LHFo3WHEKIlo2p+Daf5bgnkdUvXnqRpwFM
cfN+czrp8rZg5k52t1eWddsG+UCw8JSNqJSET9K5W56JqHZd2vKNA110KfEiNYoZ
9tCEZpuAXAfgjNy/+DXbFE1JLKY8Fn/HfoCvmEqM5XHdBGz3gYGqP5QrfSHoTMek
pj2XjWpoGJOrxxNLenHjhhJIbrpisDMUDgYREg2km9+saBW0jNOUgU5M1uSz8pEK
ZLyHjooYkBdayJDBMFyEpA2MTBnkMSDf/JKV1zC9/SKYr6I/aIw2fLZPuy35WkHy
yXa8Px+xK7jk9dBL8X6t40e47QkGvfaDJCKEwxZ2thEOn1XQTd5+WU+Ucym2TCQa
Ue7zpy1MrHRW/hHsIG+qghldSvao8HLgZpWQtd1yyqyadw36X6VFM0inEH7W7s1i
eMQOm1b5hw2hqanFTY9lC6cNFeiX6PqPmyLyrOuCbZYlEiuadrfBP72vdNbVFIYO
oyaT2YEjgA5zsFCwqy8AiprGAhhbLQm8sUbtCUg29AdVmLubNZqo8f9XUSl8MJ8Y
F7j0emP0AjzZ+VdwWomSxCX19AHH/jRt6BcZ0bS3SkE8de+9uo3i8qPdQdXXtMi9
tllfoIwqO6rjobYdq+iGdOHhjfPkmu+PMb6nCcI6baSLceaLIpwRWTntx3uHsAS3
0f4JVxHXl5zIDL4WavhqL2OPOLSvWzzYriyDJS8sSYVHZBy80GFl1sChsEmC4prx
tggNHOgNZmuzrI38zYeoPl2htLIM1bNPwb1jdDRiuprLEhCgRXH9Hvy8t/Pv3sPp
mCAMEsKZHBdwLmE/pITrxux/CC8SNCu2jXTiKA6Z8NT7JtVrhkdzKNuFzcyPLGPl
jm3ogYHNX+GZnsbuS14z52RiFZD7vBNXgO2ZCBbV1asrZniaM32dBXPPnRLbF+8N
lPbT2VWKp4DSqZeK+vl6RE9EdboFLJVOhf0ywIYrMLsZHn5GD8OphZuqs0F2k9e+
Ov9kLUPLXh+h4Ct7p5MBRwrrVGJnHb5rKDnooLesPk84Lcc5lU0koNdMqd+n85i9
wG/oJC7KtkNYtSMgD7wOB2U+V1pEFNAoOU5D0P7A2fLdGYN64rQ/H8ihUHc09vNr
s5tfkTSugGKW2LRovjUDvH304rlRwzpmFM5bsXu2saovjqerHdo+DMsPetGpqQV6
hbtvNb+/WkihshMkQvB1v4SBDaWZ4sPRas7fuQhxCxkCNxxLK22fwVryJMxbAYg2
r3kPzT6AAgkqKswroheDQ/00tKoTlvol44Lc1PalkxyISIN0AXULQSPTNxwX3YYU
kwcdveIal+KB5IB5Cg56605V5C5nwtWVJMoxPpYDGq+fAHNrJdP+TdAveh3c06Tf
vP+Gf4SideyWgos7zSD/nGIbfGtoB+dbNcsL+GOch4SdwJFQmvbIPht43KpOhHMc
HXASwVW5nPWKwUXjOsB6IF6q7CKE7C9YDzeuO4XzlO8xkNu8u2C+lTLw4ndlhtwm
TEioKokKDWF2n/1XwHgoXoXE2o/1GKluaVXwAcOsrUH2YTyDbQXQ2nzT902D87Kb
ApxlsBzAZeIDoFX08awvWyG27XkbBvvzRuOmc16hloLDQS/WaqLojk378vY2tg3P
Hj2wcV39T8dTiak1NMQUo5YjfiG8qSDJ/26xqB3h+Pjq+cxkbbJWOoyOVPVJQk4W
iSawnmk1mT5U6ukpv7uIX2QJ0+eVF+0DfBBRDzsM6EVDkFzPvJWEdJZvIn3AdAeM
l1VX4R60TdOGSjRCyl60iKHF9QjuDM4fXgNBaVEp8ZsGH341MEeNMcEIW/UJTk+0
+zyCIDE8r6w9sLDinSgOSDTTb/cUCJjKn3ZNVarTVK1+Cq/9rFlFuZRx5FXPezQ2
LA2YxRfGn9xbldoCpwML3YBx5dzsL8awT9amESaRaNDaLtGvw/P8ovgZjG1SHm/s
bPJIzKvEXeBp3Xksa3fUK2xUflp/5bWC2IFyoGJ081K0ZAkYi5/iol45ZKXOiFdp
65hAymOvvShBTtEqQcQ9rgzN2QTvjkxIKB9tVgq3iFrJRfRoHDANH5wse1lLI+IR
chxVVICDQMbZoxrgQYC3jDlQnNWd9SfoVcA/5leuDOwCrxZdqRObconL70/B531t
eQHAj+3fXHFIt/2ZQQvVnklp9i7eMDwhbcH6FjjO0dYbhEf/AQMM1oC6RCOcGPwc
oDUIENWm35G9Ne/toUpIt7w38dtWTjd3Q9aZ/PRRO2XRwADc+hXvHEop0lBeYSpS
cR1x74OMlQouE0M0A5UgtCHS9HuUfyY/7wx4AHCrvQPP9wPhzzxtPQH29gEidGdG
3wksHKpExXLXvwBAo6+WsaFL0CG52SyL5CP5DreNCo4xcjiPTLk6JJwToJbbpRoA
CJ3Zix8tcJ+mhOQKa1V+EhPqBP74CAyz0kNbBeOIdootUJ5G2eb9nn8gcl6rrws3
TmSmISGCQLBo/aa9/3XnbcOnAOB8HBmwKWQGYQyqShyuHn7YSVInlaaFY5jqScp3
8Z8k/FYiloZdKi3NwBb4vPkGTqk7jkVIROUM5BlafoPFiR60d4O8qVFjBrBwDxLY
892l77cb23g1BDHTbCnmthjzkzgy29tyGH7CbLnTowcADhPF3hjc7a6zMkNwutGY
LHlj1j8NqZiomYBSez4Cg9xenW6lLs2u2XPxmoNbIU9SmQjn7gLiAHQUZ4L0z5QZ
m+ZV7DXhESu/l1HGAdV5/1OEHXi8XxASQhFYoWq/+dhvoL/b8UvmDWGcJ6BNlNnP
9He83AeE4ar1WjppRzgWs1Kqvaays++Vcug3QPNpiUMQtsFbJxI6dya7hczlS3we
AxPfx9h5L8HimbH14QCmZWlNKK1Pmpnrm/hl1JaHd7cjBhOKDFuu4u2VSIvSOjAK
J1fgIQq/OaMD5gy5rMHV6XASChNgrpcxLx8+E1QXt6xv38t4lGvtYEabcO9vm3ey
tBLje8UmV98JqdnBPJgsfGxm80hTJ1AZFSmYHljFOiHqwmV9AWs/+A//syNMpv2E
ah3zHWiqmCfly4cPU7aKUKO8nMlpknl0Dj08r5mor4U0UulTge1BAUNuQn+Bxm0S
XFt6uG7WgdrYGwciZRuXNjuC9TRMA/HgAnc3BMzF2Qglwf6bO3dc08FyPeLiZHRb
aNtMQoi7LAe/LEY0u08pEN9ZgLfe1OObATb0ZObl8M3JAT6lT49zPShm4FofSuj4
NhbUMHwkh/sYLRMr6JkJFqOQYhiwLxiDPXjCPFNB26EAIJ2/y5wLOWJNkfk9PaFK
pkwae+PWIj7/ktEiFpvkh6Cbqg6WG8G/i2PfPZ6p7c7E03xtVWwRGYgva3xZDGOA
wMKOWu2lsCRW4MOE5/o3ehU98EkJj/IQ+4FGd/FAuwtISVSebfCHRCW+YYW0HwFT
2jPrIWT4I/f8sEo5LC9s7ZBY00iDwGlNgLOrkwzkiHJ17KEJzGY27h8i/3BGzG5y
Rc31krS+vDcmoyK44RcLhgg+rDHvL23zBCyiOUymwZa7FbBrQSPlUoxPchbHdCvM
kmVvLkI1uM/GF1G/4up/FvO2ori7JSrvNnCHmJZg+JwRNIovTyyyOy0qqqhji1ry
uI3yRf/MraK5UBU58UdY1QC3ELsuhmM4Grk3bP8fzLXl/okTLBYhUxb465xLHv9Q
wfDQVrJqNueXEDUynr/mvSDi45nem5ZJrYV6Iyc751N3MPAnwrDSR12k1/5a45rB
ysVMkDZi1CTz6WIAItyd/bkT+UaZxVNfaRIiZf5QVtR4llCPPbtgYPCb/lnvAW0c
0S+tc4of8Ie40UDC862zEUoRk14q2dMShcduhlN7D2IyPWjmP9ZmO3dw6yiEBeu2
lVDGQUJXSHT9NFKKSrMfZ3TkvsDn2DGFg38SJVjz/A5B3xPFb+0zgj71icYoE9Mb
f9rjeGZWHI8+7+DGznXF/ZPI/ZFAZ3e0yn1N3P/8bxx44y4RicMY/c5c9E1NwD6p
F7SCzeuDaOP1liuD3dL9KU4B9MMRw0pW19SR8xZxOdLG8kXf+MhtCYlKcU1Umcju
MN1y57txN/NNmle1rAQpfnIWw0rySMdaLjVOWGcGSHI7VgGzqwueG7ONkCaPlowS
wDypmnvKT8+CN9Dk9+aUhaYIXuAoyMZN9xvUVcUWjO2nwxsXYvkXUxMx9MMno7SE
9wOKM2xLjRhPu5e2LztmYIQmIdURFUfVR4n5VeiRx2oTmst/1MIWEITtWnDk6v1/
HTuvI7GF71Qp8ymmMBMbxwIxMRGL3VF96/8Y/Vibslg0ExBXDHu6w5xHMl2T1/ii
wB4lmiYk937exl3SOsUbu+et0uuaV9c7IBtmaYHZIjIq1sj0jmWVKqtTLR1fkuLo
AVDLTUcM2xGjoUrhyLg9UlFN8hL8tTsWf/z3z6uCJX5jm9rmVGaTpkiv96jPt1+y
PLDlcpd2k+Qe+eJ9497Qk+3hvB/CiUgbiqwljssmMY9huaiNt9VPe208BHH2McpC
XNzifvsdB/DcyxCbFL5cdUH3ZRkQahynqelfFHanPpbo2ffP54RBU59YvZ3dWRQu
kstam8HwnkAVTilr4iJ+n8tpj2dkt19Vf9cm6gKWFny6QSz/MzjbYr8N/ZT5qIpO
LWsGvoNxogVnmHK4r1dJnGtNa06bOo5PgnFwI/Nn078HAFgmcgqulCsN27YiIYsi
6ArvZgVyoudqV6m71/ZCQApOqFA2Uz81AfCg0id1RqfjB9AsWflICGo7dMZGbsjI
bVtjGDCekkK9RyihZ1UEpgs+mWjeVaur5Cc2135gGA6p34CksZ9Vptdvl6lfcruL
YbgxxYc3Nvk8L6g29ic5i8gsxBDVQ6yRyfvztnOyU+FjFNl05Dld0EWtI4n+jvDg
ZHJ6M1ujISaVHHqvH3IAPjE9O4551oAZKminv2UT3IRExC8G6ZXEUQjI97ufiYZC
eCby3wCZtskc9BstmbCuExeMJjMg44aMyDKI8NEItO2dsyGyDHrLNIL4mLS4Y+b5
BpQmWeyAlLOOWctnakA54+js5Nl714iROqiumfwwU6awLSaCF8z5LCY6z0IgW33e
+U+AY/Gc0gcqIZOHATRSSHCi4dzEIgRa6oLW56GDctQGJ9ZCYRbijj3QNN7NDDtv
VN/myLRn3E4Ucz2IEodFT2b1vLKaQ4rnFANxJyqEWOgi0awq4MJKt+5nS1Hao8OS
s1/rJHU5lOy6dU+l447sFl/Lf70gsIPLwzMMmK2MYr6nyfcChLUiC9D9pBv/wK9f
xoxituVsiLNqc8qKghkinPzdsONB6h6aUvY/hYdPVwlEUmC8RGgmL6jTEQkxKUYW
uZSZVB8MhtOFZicAKnr47VcPmdjItzH+EHCyIp+54/2oqbVzXKkbLULzgLSHeNCY
vC2aDTdeqCj2oHGofrDLDfWqeWP4y6LAvrTH6jXujiPaKRvkzFXj2MCN2QbDOwiS
UtXd72g5WFHSuHQzhv3uRGlrxgoCjre2dM0aCmzsMgpKpWLyib8ZzOrh8Fy5SVJz
HW1VgEfD7LB2YpomF3bdpv35w8KnEt+QdKDys1gOceSRoVvN4oD+lCmtfINsUs5x
TC3t+urlKzEzIsnqSmB4odiEpbx746SCA3HYE/+ZxISichcR9DNj0m10wbXjc1nz
Nh807OHpxhlbOa4+w8CpGK418G0hkUtFVr7E1Jq3Ra1M4mpKgxWamRprGRiKJnVb
OMWc2OQNnApKrvHW5kSpBeve9aUJUk+1lZCEz3RGSil9LU1l0yTtRMOSNQJWGfnL
e68+Uqpw/sY/+3hF3gN1glpEQi7w28zYWx+0h8IskF793huUlwleGtJMqdUXZo0i
g3tLxCibxCjNI6PdywmU2xAtOhC6YwzqUVNB+wemaFV9Wuehp7mMjWJjmLQBthx+
1zpr10JVqbWjv4Ud0YaG9UcPzyMY+SGzPhK5+fpOzTPO20qgOxYj49G7tp8tgFG8
2Md9HuDs7YikpPXwXmr5SwE+UpK7Rp3g5MbyNfIzYcwgsUnOtbq4fyWhkd3WGalH
PuUJ7Bw0q37tScnQrdKP5TzfjKRqqdbu3U2VKXJt9r05zfdrWAQfv/E1I/0pRfgP
kqVTc7iNAtbMyQTvUns3n7HfPQPH5hSOq7ytWSWFkCVhIhqrUdGzPeP41/UaZtJM
kgJKE1lF1W81UBI7DsC78zq185liop6WFxHaBY4lVNtlxTEDPARthsu2j0CRsXxA
zmeDVx4ZHRm4X2osevGDpjIDl/wbAftiLHV3Hr3fx0Mb5JHyuwpG7w05VIuCt6n9
aMyKc2kISvxSc6syV3cmX+hcq3C+mtntnRaLJi18pqZenZzlVEiaV5SyR1wpuA3/
EfISHQfH5KxGcTdEp1XlcX+kwx0XEfxmF7RbxalGYy8pa2pGGyhuBAfmQGwKjGga
92rqTR+Q+auIU/R+trx33EBlk89H6JxHkmbzKOzsp1C29LCHMM0UzqVmLw6ajMY+
eRKxesmo4Np5zzOEPOuDiGFL4GCm+T8CZ6zNAEgzD4B0YhXwPOHMzXQ5yAr18Blb
osLyfGNC6t4zal/gKiyX/A708IT5duhBDGc+3Anw/fg2glHQSLoPfxYj1leA2E2/
AFGLo4oJnJsZu5DZljYpuWHsNCt5RqpIvw2kWX9fIYiGmTQLYMfArgxWA2lIhhJp
OHLqsBxtKYTZGdnS/YObtbDyIkty1sJeJDcrZsEgt/CTg2kFaa5AWyRtb70R9ema
00yIFS5hzU42p8AoNCYa7mim7DNHtu7ozSxsQ8YzSKfu8l06QDc06QheAJRcObrv
uA5ygm84IlpN24MhGhom2in6sQQQAFs0WZBcsVPWzSOHE+L9Ha8Ohm1F8AL/+EhB
I53sSQkd6PspHm6/fLkbyVMgyHx+W5v7lrz3LDL3jzfAAir8Ofk+I94Jo6a5Y+1j
j0wILVfEHGVCXomDRbX5CKsb3O0PgHgdR52/luXa0wAfgZCGiXxOapqLDAUussnq
4gC6hLmlyCAna+b215+DvUWgLtvuYXWbpY+pdt8jCv0NimTAHY8gZdFmiRwiN+Lf
2aDGbd91GyvokW74+j1lF9dNkFONt7tjYDT7YEVbajgj80IdrP0MOKA72f6r1Jue
9pRqsjSnpjcZtS0o3IpJMbvE53amoYYUaOx0Ytu0qUmtsEWuXk4cB6FGWnZEkHRs
ZidqNxy7H7Kt4HISfCWjwNOAK+kxbL/B6mjOazq2BFI2XclI5ZWKE8oT08h54c52
sU8mrHBLTBMUsxkWS8bggK9kYCdJ6dJ3XoWBZc0Pba0494dzsuOr2SoR0cR2pm8s
1JBIX2kYUcgZYaLNNTCWHUZ9r3SjdAtdqREbnYUO7nfyZ/xbKXbfVbZu4Nh0Z30b
ZXHLV5OhhA5ryPL3gbBksRZ2Dx157YgNFGaEPbzZxMvpGb29z4ujGFoiiteZyogR
FmLjtDr0ic1Pwc8ht7Z00ejlFtFuYo2bPt2+haHehb+jEcpeD+qgZD/ak5MPO6Yq
jPQjDigeUBeS8qqFhuqkDyECctKB6jc+d4iYGnFVjHiONgyCFQl8QcvxwEbOtiae
9Wle7GGr+svx7L0sFrKjp7ORKRGpobLA2OO5hv+zM5J7AEfTwuTi53GbjtLiK9/I
siozpcf1fxRkQQQqCCeBZxqf/K76QSGMuyXzHP70ItFwW85veRyUqK367hmJyko6
dpA1LfZ6hN/JSj0lx2GEJMx8bEUwNpSsYpVU9ndwfxkEGXJlHhlXQbj+ZZAmUwxe
fwvLmmaWwL4EeRTN35wDj6PnCn5xEVmT+KuWYdPxJYgy0eWxc09mPH9ZVd3AxY54
e9/WQeBN6bmH3hYyUmzts/vVRJhuVQ4YNmuQc2nZGztVOmiyHt8Hw3I1bdCThM1P
0S5pVWIdbd5C+v5sH0GXxA6gbLDohn3irzyQ+Uy4e2tQkGCIA1oXkHU8P+6lQL2I
QDqR1zk0sw15qQJH87fvY30YkxAE2Q77QWpNCPh4xpH244SEASsGcw5ptRTVEN2J
fSWg5aRFIxEPbAtmUxiKFzreVujWWYhUWvtjrukSQK82ijrUeE9NENPA1y9lkJDQ
homaZtmx+C9+AQEyeZQ7khiRXRyIBrCSAJBNQKPUUes+NBjjHR9nIaAMOuvYl9tp
wJ5tbynnmoCtQXBGoIH1LUTwGIKLEQ0xZJTHLMc5FTXmoFhxEWCgpecaeMoeHVgm
8FgGlH+0+R0nHy6fsCZIPwXHbubQW8suv4Y1yk87ZM46TFsDZubLNgPx6thto1wW
4kxAvrt6SRmqasCWBCxugO4m5kIvCaInWmXNgBC4n0fkHYRiq09garj7WGrPObGe
66eSdDV6XBfeplT2IHGvqC/K10C01fP7ZbdxLkr27Ugl2jw8tFpPbBdBilZ+9aM7
yQ93mfYUrfBmK5cYvU/EQEkfLP6j6ry8dsrisp5I5AmFcthV0ZMYPo5jzgMQ8nH3
m/7eegWXiLqe19B1mtMYH+34ZYz8J60SuOgOcpFNkuz/3o7YMtNpyKSjGUxGFDPU
iZ7x6LjahInyL+y3/sjw4ez3FYTYPz8xGLzvrR+P147JEvu4erkmeQoLjuP6GQBD
ZDM5oiYllO9D0LFovTLamjztOunYKdu+pwU5N0dZ9C1OdypLUe+5+xWfDtDECk2t
AsAFjkNkb2aj3Vcey0GlOUqex00YCZKWpDGC69zPHubGCTTK9jB6PWYN6ndINWfZ
ilK41uTbGhFIpchW5O+GxmSZeTkkuk/XhtROdk3WNO6gjFklq55QTIAONmONy6PL
HroFPsl6E2qkLtU4i4MMtovma4T//eUr6zw1JYi39X0y/cOsya7MpGKTkdNlFnGt
LvwWIrotdMrRtcuPBR+Q1FQyJ0nSlJxSUuYBZSk4lryiL+SgJBLbwZIm1x6S6qlY
Sy4eBjeBwOnNlpIZHwkz5puMEW19PR2Qh25R/Di4VppP7lgDsLq6XeaipjftgHZa
qjA2SeyoEeJnycucUCFsmqBgc04LuI8eMX+pn92pdpx6ko05d9Yd1a7MALV3+nhW
fnOTZiu+6buoXeUGiq3II3Tj2caVicS55vEFI09wX1j/xdp9lIBfOszPv5ygrCcK
vdarHrcwLzy3VmckbgrSbkVgjhkinKQLsdijrW9c5soOAd8/Up3qywo0B/BeoT6W
kJzUsyH7Wi0DEEte7Ww82JrGsw2ltStTXhAUfFkKtb01dECaNmrymo05bFXiZI8x
8HbeEC+DqpczPlIMhlSPQtbhwTuHh80XHQheBDBl4L0mfhAPIF6IgLQC9w7yTWYK
34bnOBFiKUDxm82X4L60bycykpblhyCtfKVTDUNF8AqRQYsvKcUSpds+/nanfmZn
yttFqBpB06tEhA0Jw53F9RrcarsQa3DQ6qdWATWzq860W3VFCcBKghW4vJSICHtT
Fuj0RQhBnUSfitSm/EsPn6mE08GgK4Uy4AdOs8wb/Fd0UT7haCtNMvcuHVqxp2kO
WYRgw6i6JKCV19sgsmyprCR+EGBzRGjylqmGzYNF/n2fwTTEI689AoghJ1wotEJ1
Vege9EPEzn7+b6B9kwc4h7Bv+Lhf02U4FUdsWaXYQ1zLw+zrX3kqFWq7uGEgBSzP
Cgfje29I9cNoxYzJGhMT/IbumrQ7QnnY7QdYbaTiWNZUVyTFy17/cmPrVjP+k7VY
HKjrA5bhF6Y+uFmMldG0yijpz2DX9WwiW4HvYm2yUlK+bCYy5DpeZKbQoledjG60
mSW8B1ldxdohTwooxOur/nYyQZhhh5rkhc1T/bjcjwkgQ/I32HSyznRuzV6mtrna
Kc27pO+Offwo3oAwm1VeIvYmBf7sbALg41tZ+2zjIl0ztYP7CElLuamjaNFOmpya
fVPpiavgarbK6uIHNNBe1UvcYXkZ13LaA8+xCxuPNgz+WvhrQr0Ojvj+bZU19Wam
NHXUpp7ZuImyrdCgFMUnDjvjH2qeCq2mdEtl63FrHchiOdG3ZmcUUir0Vu6SpN1x
rNHEIIZpidPsM0avdgOpNHY7DFs5tzl30mDxde6RIpLyNKMFDU1PxHQW2YBBL7p3
Fxgi2ODiFBkmuOI5pUsSByCFjpER+B4p8IriTOjbya4u1WpLZA81fUK6sS9ZhLVl
U9Ou42PoDsxkprhDE8mCp9gmER0mhDVmAPRy8bkWQ14ylfskZu6JUBE3gYm73n8T
13yI3KuY9/sxCG52kZ2R+iuw2iwGP4YJQqaoBOA5HeTQBCUAUTVDjGgtxoCHsKio
nTTZghEf8gKh6zCKLcaNDV4qMjHazCVz4UavZFg8EgyKNCwgke6gx/LEwPFceEia
5DQcw8aMu2paOV7d1IwArtJOMAumFjz3qjhz0EIuXKEZS0Wq3eBJUJ6Hk9zUqOFB
uReojrvN7OCeksmJAMamo/uyL0xZ4ElyaEDJ5TsHRUD5b0NHkNqtj9iw9kvM5Zia
3FG97ot/AcRtE8EAdHyrAGQ9UB5gLt7uI7Wl2FH7gBfMgpEDcSMnszvUwLb5wped
pxn0g05pMNfbN74RtJVg4PZD7qv1v7E2tDs++10T5jF8ukN7E83Lpzlp5R8MxyFf
pY0ID2fCeJW8a2xNpqUStOU3/3rcJIug4Fm8GAvpcWrZPK8+XXSY67FN1HG250QA
EYEcki8joUYSZ13zbzgbGy9uJw14KQUXoHA5pwJ7y13BCCTYGZ8RowHLWt3OYB5x
W49opHjNqD2cXlBl/L04tL5PkOC2ud5QwpH6n5d/tnkV62FaPSo+DDp+KLtA+Bqg
i/c/k4QMGwLG9bzOSkSn79KE8hgBBcT5plRzuvzPTBEzetLDccdDnDMg+AYbtMjR
n6wjEtXVO1/gxxzfZNWCU32RDd6qvwMDLzqjMKr8SeXQdzHh8pL4O03rLsLttHGy
lFV/tVHvVeoJFJ0rZzxSXnRF3zmO+2QFCzBX6UDuVDM7kZZm8WA8cn0FHYaLSWzG
m7kKVWjLW8h1NlY7qvClBBT7JHllF+Q/66ESoilAEMwBGPOOCogvQWrTB/UrspN7
jjTv3QcuH0LZ7BQxPNIXCFofIVl4BTxwj2NtlPmyUKNVTZTOaI98ItvLKMxA4cv7
NSt6JQ2E7kFWxu8TW8dE35/TwU/+eghS47zAmpLF5uQIhaaEuEljXih4tULHlobC
Iz7dZNK4Pit0gYh+gUoy2KjEgcxmjOTTPl0HvU9tOwpcHWEAPWkSCfXONc+T1tJK
guJNjVSWYMsXHqFmypsukzmKfFs1r8qfQDcmlpWtLuOG70FpjdsTJZ4/O53bARoi
Z8uzEfACSUY9qPIGQgqdl3baXyY2cJzViFZXR8vCuo3vLrRNUcY5dRNEsYgZ1pCk
gN4IVankWaBMN4Nh5ENDgaIy/erUPMlIncZb6cR0hdsl7lndA5iXVshqXN6FmhMD
PtuOu3MKOaUwosU5sE3PTWeoWKxUlxMvpO0YJkYU8wJ4TJI/y7Ii7J3Xw2rOXhjT
7f8Mn1AbF+ltDL6/u+zsH71XjSPJr0tJSVanR7c6KWUVCMPDdcCt8eTTANJDnE32
ZZy0eCadlRjDXx9bpFsBa4LYxDkH8M9teyPty16rHlkCklTfv4Z4rnw/YpTdR37K
GFPM6Wt3AV9DYGBf4hjlIZFdGvT1xOivR7YvGQqAp+ZeSNYbxmSr6inUKtuf6Lf+
7pQAlXkBbl2zTs1PA5H224lEiY8DCdC0jUPccXS7yO85c3hxyEifceH7wYpGPq1G
bGasLLu9n4E3vCv9a55pJs4BFDzVBMA8ym7aAZibm2YywcOt24m007MvkbE7zhqM
wuGseY3VBnm/RwFroFXaUemsCmsXL/HidLoXyk3obYbK3r1C3SvE4D/dm7a6yMuA
+DuFqsiRWM/J0Erlqa2nzVdOjahzfUjuV8Gl9Zrh1xY8h7XsgUZQ6DJrv+AyOE7N
LKHZJPYux1IsZajg7Nh7AtKZBQqR+5GVFoMaG49YifpSIxP3s2MytVBdYiNFJ9q6
H/qc2CkHwgXj7uq19+YF3j0FACiZ+gg/LH4kffyoNxTTwNUM8bfYqtBxH/4qxD4D
MmioWuNuRXg+iS9pzKPuoq+DVQmJm/PNjiWIt8BFq8o5r16HcrhcLL61vuPWWzwn
UF9/OcRWZwbrlAYUOuisEaiRj4gkQXzLRtMEn7+/rVrhnoae9g3G9FsDc6OrAqTk
9uTBJHCVLo3DJIv0gTWmq266/c+8WQjAhnu2B/qMpOo5aHL3pWElU4A7N6N+DqVH
iT4n9UKmoTZ/cLYkdnnFWlcP+wgNEeQbn2MvABnqukYfMDM3yho1Svn9JOkP0CB4
agaqn2rR8SSnouxXeEtAYgnMSqYjL2H0NbgF5r0hzou2d5IxPwQar4w9C5rgBZQp
v0VJKp0v5nuDTtSN7GPIhV5+pfdgp8Ez3XAR7whaW8C9zgFXn8khld/1RZgQ5bt0
FJZVlJLXuQ8jxKB0E9GcWVH2ZVgpywXUM88I8kaktg5ytbKSZ8x75k7DgdzS5VEH
EcDH7WxBnmFrl2vJYGw+Dhqxc9ngbPP7fCKqPiRhQfYPx7YVOr65ikFveFqMBnxr
9dGE02YKafnUsP5RpZs7qCWjbxPgDUxoK+deeSN7Og0tWKywJZRV0yiRxsip9oe2
DWrSWNUcUO0Jz8T6fW+TeF4amm7xYHN0tMYwDsAQAvCrO9AtzvKRHi99tR7fw3qm
o23ybQDJyRdeiwa2x2VM7PJ0Qikbw78RGVSFlE1kygfiVWTIf0uk7sMlgMHRZB93
JFhmI75VEOMtByhSDtXCgHgx/3Fm23dsyzDrsDoQHKctRfm0iuiFmmDAVtMhEz2i
RUblzsmr94tODK14m6bVz+mPT+707UdU4KP6g61bcMtcq2ypZveaHBYdq0aiEyMl
P05yxoGTw/Rs+jbBiFqjg6E8mA6fqFGZhvPwUUBUytQ+koY430xTqI3KMvSrKhKc
1MYN2Dbk+MRAP5yM29FF+rrKEWcs2Ti1Oz/SIPuTQzQxgywQ2lDgmDRgUnLx9LtL
oYpDuR4Dr9gWiWD/HzGn8VemFu3zPwGauvNs5IKtuags4G7cKNdonwN+fK6ZTH8Y
xfJlA8c8KsJI/F/SWhM25elLDab8JESIuYQh/NFe7DRVg+IHUms1vFeD5ZjQcSaA
FRTXjSllJ4Hdqp8Rmbwln06UgpSLhUdF25kAewX8hSVrblnZ1HXGTZLtWubAo1Md
6u+qE6apNklvcb8sfzDpMothV42VYDO+jV/fs2471Y02CQ/1cNINnhdNuqiYyKQt
gGVuxf4NPuhuFxTKVZ3+uIIObAster4hQPQxJ6yzVkdiqwqPMiUUFtJCLK2oa8k8
bo6nFC1+mXVHv0gqF7iZLkrRjx3t1BxJFaaTYp3KaNEj8pdH7qDI8rpplPO4+Zwu
8uqhmH2xhSdMdHq+2S0ju7qlTcX/3ZM/Az8xPSMo7w/W+dMfRgPd6Ha6NLgkeGAu
czi3hgnu0LjnFScaQy3vaJDwEHP1KCS21B1YkXEhugDR0mYQDt/jLtwtEhWabyxe
EqQnWMZeG6gkW0T+Eqlh8MrYMZq3CDoI1fW0h3v7VM1G2/u118q1sansPR76kV6Y
9DDamt7LoKEVpvkM9cKOm5NPEYp6v/nm+sKT5/jHTRL+6ODYvHskAo6ISEbFVAyv
8/oSMn+2ipUQ7sdtF5r1q68kBKlsXr7oqQy7U1B2SPtYy52kTrXxUFceXBR4s1iR
F9QHsD77gpG9kKi4AN6NzqeAO5/HCFXRP8x5ssqeEpdUtjj0l9XLy7wrz7JeFZaq
a3ORC3M+XqFiJeVwocwHueQU0XgUwK1dTfb4NDK9vUdYIYS9se+Y417nkWusXr3i
PKohGdIsV5Wi0kL0acX5Nv/QZ2MC2ecI50AAZpyaKZFP59pid4AUxqDMlLZ7Tax/
xGCe2iEoSl5tZaMyHdaCxA6RoAQAr0pI5+YhVtOAQyayE55rpoBn9cDE2nYR6d6P
1fHAttoivjAEYrNcstRJRmJt4XF6iB7Q8C1KM5qqTa0cHPbeAlen0SkLynpRW2d9
lhJ55JQwz+uuOoBrUWWF9U64HQRcnmvuURqWFBVbMscWLZYpfBk42Y2XEQQpXevj
t0G8eB4Vx+U6BpfIgQzwhmz+AkLbXtEvt1TQhepLTiXB3smzoTf44CB2gRfD3Pt0
7kaUevOEzT76eV2AgQE8ijnNMO3oCP9mN590XupVXtzjseXb930mhKIszYSfxNOL
LHMFUxFlwcaUel3w9Qv8M69R/mhJr1Fm/iPv/H5ZcQEqksNnwKr2aV1kfdxBjIU+
uLf4X8xtZaIQTzvWn+zAfyGpipvEmLLk+eO4gO76JCURay9JLEmmy7hxokuFaQTy
l71OQX1GOe5Bm+CKbD+IQaaF8YKLC63xsynxEG044/dUNyBC7IKWJuiFaT7PINoD
2kT0HFPlMKrOW+a0IHKmL/PKHZczTlwIzNVOwd3nvPYyS9l0YRvVJKE4O7bxZoYo
fwIIpZ6Bj56vy2KoqbvZQ96SpqW+a/41DePHsAQbsHtkl8jQ86VaBVCtcdqXajnu
5IMg8cZC90zy1/LO989qt89VTjr6xMXc3kC6YOa5Zps5cXBaTTzwwSqlxF15x3yP
boh66VbTKfe1dj2PHO7kXvtb/tt86LerLddkAPncgy4oEtgqbDtd7XKVAiPvJRl0
ypM1sUzukfFLI6oaNSxUxStYSTyrGinazbMcgZr2RNiDj02mxIl01vhpjgs5zbR/
Rqt4c4YlyYrKrwpvVZf3P/kofEKmGs7eEDGUh97lriA9nRGBVNvSALNtYc+zvcQL
TWlq9DIoaRSOyX/OvcNbjRVi1jp1wLH4sy9e930Li5j4BuFOZ8YYnlZox8jBFJnT
BRg9YQTT0TVYaQKIxr2X6oiBeAUTsOY6XshJNF37RQDCCGcKqEUCPtW7PnJ0AHk8
NCbpPCiLhZ/mwMb3iojKKKEZuEfA49vydvgGxjs7NT4wjBMSRcwCDmHOUxhcVn3r
aWopwgvyNZLN5jZDkI1gwlAgUOnDAFOJFv5trChh3mED9alolddA54oHqs1igRaQ
dr8Rt7NhUBebgxv6tYb0MCeLvILHpNHv9NKr420QLHTOwWczImji+oFnXYZ3YUtL
z8nmmNcPkYjdAHeIpiZ098WR0HMFRVaMkPZOV+aX4OBjfG4g7BK66TEUWHtRIgk/
zHqZWNjV9LjM1LcXMBAB3zYBUzm24r48iu1tq/v7QmbQkFbAy22k9WFSuPiLPbzJ
0eBiL8Z0MKw1lSO3BHS++HWJz6XMbvKTYoFO23f8M6Tsea4WfR7o+7xcntOS1WHC
zILOZ+jBFXIBBM8SP7nBxlvPg9T2jebBh5zRIm2jX+9pvlXBwPBy1kNvk5D63CFe
ZTucsHKc8aHNu6M00DVPdgKluWtgRXTEoUBLy0Xmla7/o2VWCmHmW3Q5ACmIC5xd
Lq6jfZI4evp1nrRZ9RF1nuX8uxq5qyculhjW+q982CKAO1EvPP2k9UAgaTpTf9gY
M3lII7LEnQ6XKjBCNxRHKGNReTbeURTgS/yJVr2RNOLm87BdgT0RhMrfFB4lIGXs
YpQfLe4U2vG/Kcz1eEgLioNeuKjPEE5tXhdQX9hixoASdxzbMzK7uPjTq2pCFTqr
RcIGrJm95iB8iLPE6sOS/SCQ96KZhX1Hfex0PPtY3xbM4st2fhXT7fi/utSiOL8R
cpOMUP6EBraUTYYlg76VvWVd3xU94HqRGHHmYifqBAqn1Y98a3eDfXIZHC9bjst2
PzcRqKxu9bS8fKkS0MwwC74wlE4ctou/wnPgGfOBbH5xHVrflfvA+W2bnpZbHBK3
UcvQiEDV85tSM3HpubeeNgqQGqYVhSOzPzpVhjCr+KZNiTHuPcMbDs/AFRm/d7Ft
03+z1axl2CxW+22SA2rBlMEudkmEBiwkBS3MzNnAzDTZgQ7TyFTj8ZHlAs/Gctul
2xdDx25zYxzSE0FMo56tInRi/cfvG321bmlP85aZTtx2GLlbZUoOmxttwycoRc9R
0K2M1ZLFxmOHg8KuD0mpANeYo9a44kQF4bsqSY5bKQ9AxKjQFpQhPpDwQiKPXfN1
Iq7d9lQFEAC8KVYNszQgx5CE7vnQQTW48RRyeyuiJBiX0GW3VaI0th1sDYZinb2w
aaUC7PG/l6vpnFbkt8LRHsE/A/PJppcMrgYgKVF2D8wcdEQQHIVjeasF3cgR5Lj0
NuwLyvBx9N+J/xjIC98kOkKDZD0OhHZOeN89wRR9Wu10p573VURUBh0ITVDBjg1z
qXwgfI9aciR0Y8+FgOqNCpjKoGBikI/HrPbcxfhaxDS6Qc4astmrnD8tqMsti2b/
eT8ZAFEdea495jK4dw8ol2nwxyphoTU5WSA8am7qCdVSNSIEafXCk2qVNaqVta+3
UbaSJAEGfupSmdunQld9DDaJk1vEiQ2t9z6DxXPbjqZn4/VOwjD1bwWdqzXvPgWS
j2wmNSjBa328moJNJnBGKq29RA8XKmPpjIWa8Rw50UpSGwEYEZ1a0sj4i3SpLE6y
icT5z+NdN/OdRq3IEYdYIaSTs+KSMnqYtrWWm6wRANaV2QwIbTlxPrbpiv1rFDnz
yuu2MlNT+5vpZ99tS7ki2HGXMm9X561xtiu3/fSt5PwP1fUI4dgrnfbYQ08fDF5v
EO/u2qZzVSpZnw17jbiDJXsL8CXZB4221E/QHseTNcFPq8btRwpfDNuuwQqOKNXT
TVIyNBxkUC+APHHj+4mHjmrH7IHfoWLl9aqom5B5e76wRJXb/Ra10361WgQad1Cb
fyQuHa9cwwCqJNxjxu52uOFTrAIiVNNdzmcjmKhIuEA18gSR+V6kaaNqVlzPUPnD
G6rMdu35xxg/+HXqhtB1H0LjSvyPtDE7UEq04rlPrhNLG6pODlNfp5YrD36uAK/V
X8YHFMTG5pYo0tQ49BcJd7VaBNm8hO4H9lWrrpxNIzvmJu3hY3tFCAO/4PtLH4Yt
4TMGx2uIHPeRXSaHnfM0UDqhf885+TK+S0HuakQMzaZ0ckycQ3WutrxDMNrpNd8K
PvGO/IHVwfUYRrcgbIZgn8+O9Tl16c9ujJuDaxQyQ6bLc4JPVyNQKWHPtFY59F5s
bWbzYjsUfhlEKca6ixGt9iOws0rDwlO3f7wwha8G1vIlkiugy3Z9lJ0/BqL6Ei8V
1WjY+SaYmPtZi4JXwv731VpdNLfKUID4MfxqVyfcdc/E1Wz4k5ZwQTaVZqkkJJhP
r1+ORdDORprc4Xt8GmJpYGRLUrKxxSifhQVlP4bJpvPYOSZ3VU1nWnaC2jO/yij7
I4N6/h9/I7EUJEYUYaApzuOCT1c1ve+ldbOdpw/Mnp8srDr2tZVFvxVdgK4PcOln
snBgZ50T1K2dnHd4du4QTxq4s5IqQoCx5Lx9mcsZ7lj0/jMVDJT00FVXtcKp9JZL
GraSCUvD2F+MZJv5JT4rvsksKmKBX+cewIqlXT6PWkmHxuVmbyL/PVNkYG8P7B8H
sLNE5AEHkkntFfzstnpTZqaioqTX2kbGWY+b7VSkqcb+zqa6HLrdqjsvLpZ/WJ+x
3akoXgfDFn/lHvNb7NmHAkkyYNyC4o5meOt8AU72t8lSeXW1t9+97AZ4V5OG5p1w
q+8nWIql5+NSFjGodiJhy/ngjSAfxrgqo/v0cW9K6UKueFoV58h6fjvzjqXJLB9i
dNuSbxVHToVVLX4P7JuFT6FdRBv5Yb5XKwIMiVPYFwu3ye6jsJ55uxpvraPqAdQn
g8U47DtEFRRP1tTmjV/Gm5ZZhLq2RuM01LOfZChHpdfl8e2TDNn1/UIi0c+knXf3
GnW6+OP8tBoGBlqTWoLlOXKFIOQZZd64IPpdYfiXxjs/V4IDnM1zD9fqSXX0vXTB
6klJ+7IMnJnsj4nLf0+ZOtF0kKT4Hygzm5najinUSa872xZIG0agLDiXhtclLD9Q
rFlvLZNN7BCqHD63w8vzA9rhaMjNsrluXEmpfhNuqHg9hAaFYKCIQu40nvInp9wP
YXP5x/vNrXfdtO3Rf0JHGRAK8QdSs2z4HDsCQlutXaQMUNjL1kPxFd7GPjUq+lbo
iJc1OySxUHq21aPMkXBDItGjnc9dKUnJzp+ytWQEPyLdLfHm5/hvok4QtzJEHCrE
HZGa0ipfvUoiypMAtp4ZwRPjNqn5r9aYbwTfIEkvGhVZpNNZouYkGJshzvUG5Vb7
YpDMKsx+OW8MBp9YotwXuoNRGLoq+7eZSPR1jipRXIKWgwodB0cN3d5TN9V3Oa7A
L6OBNEQWfODOGXAqz85kybwkUUV0/0dGa+WcaCxnLtnIRyY5+N731buP5GPu9LeB
y6fHUEIzlhUSCzo3FKrk4jkcCVihyO5j8k6a65D68MvtJbBDwYvjgs7yB4XL8lyH
x6D5jJ3xzcgkbkd0dtWJAEYfj4t55kQySSvo2CFHPnBYRzgyK+w/u7mwEgeb2Xtw
9Y6JVTybQYbqSzesow22wnGjfqoUl8Xwl0v+WQZaqJJfVNhxdUnmoqCSzzN3kdxF
X8we2VJKKT0T/YMcG1KlgukpXRp1Bi+VMzC54HcoUHWYQT0pawIjhmfNbr4kI7jX
3LLtI61F6g308SpE7XUOSkKhTdFS8DN0bYds0EETnkKA+o7Sb/zpgvWnnE6ek7OG
V+xG4K5OQZNZuhnP8p9Csj5ML/QhJNoyePL+4xP/foQVTPsR91Z4GWMTy7WYfheJ
Po1ds1O1to1SpDmkwe74+sNdLlu2y4VGQQi2IZRHHk7BTPx5M5hgeQzntDot9LRV
NQXKOMMNiVZFVu6fbFwNfDVS385Z5bWc2vP1uvYJiWoaosO/eAkTiD4oTqcROwVm
Waaz1heGh4iQknj2yC0d5OK5A3zJAITDy4T1pVhtsnZcBTn0yLEcGbBvpJiRuhlY
C9DpYvMDMaxd+pWmHKyNLx1M76ZCgXZ6+14ynTxo1LE+iQhtPUH50i3DXcXdtsOk
Ix5CzoJtsOQjJ0oljHLNapWLGvybwi6eRYQuBNrjJF2glT/cswrBYjI783j/k2TU
53HEI7XWiyOeJHBFuH2mAi1MxqQKTQCWw4aI6bhAfoU/ugaqoGpxwMHmUBCaGdC5
E6HlXq28zIOFjAklh7pvGZ12CEfh+bSXxn1SQBvqXKxv1hXlTmQMcPvCm33mft56
Vg4UUDwohdc5HPCdhNHBd230Bz7OB9pBomtrfhrV62juM6Q9z94NOESVRyXoe/08
BpJ+zvmFcvpnjFaK+sYmgImBT+D3kwRvaCeyRUdEvEMFVbPlgJd0qu2Y+J62ndSs
C4wsR4EkswHJu+hOGds00CfTIEdKTJVxDWpOq2dvCzktulebW2ThKGTG02yyQFQe
kWIggpaiz4iGloJagSa6Ezn+QoFhNja63hMPtvlnnijid/u95ilLSvNpG6LAJROM
dCtUXkwGofIt808vZTUwKD4bTock7ATlKlObjlMGFhKYF0+NY9WGxq6faDJFh2g1
czN8rcXGfhEXisRMCov2IJxenSc6a0jDEbnZfZwOFeLqisjKvakFSMS9LNW9Nkkc
0aFk/GcXQqMGKrvthbAE2vGZUpDu12BAVIEI1x1iI9XXaAcChPLZjdpW9Pp4dQzp
DCEUTPEL6rFSRoidHjH5L2L8NzB8NVmPuDkjW1pEFWgxt16iCq93bz7qWeolHVOb
y+go9EoIKcO4sfjwKh2iwuOFmgMDI0DT/DCUF8VmSVgbybme3Oug/2Stp+TdCIpa
lnHQqsHCW0/zuZMg7XmSuu0N61pCHyRxABAEQSBSPIZhjZVMX/4xrWVTKRdwMquC
pEBO4x84JFt/FbT2L+5j2mE0yGBJ6pAfDtdrAmP3qDE1+ILBVN1lz3G7As874nLK
Nx23oXPMv+/HTIvCKsO3m0lNWNN87/j7ku+2RaZ7XsBXv3+bCdaoOMjF+mf6ABLr
lWVAGz4LkHTfZJoYJLLmm4+VuTnyEsELdGU14iHHEKcl2qNQamjWB/pLQmYsC44J
DUBCC48pnIIX9xKExNFaGyVBkBKmMvtCt/7ZZ40MOsaNgo29RrJDZbywJV9XnzAc
xPOfMl0QsQtWf0LqA/ScDgPYVXPlbcR9utjQqDqhXXmEPR7l7z+ZRYHmO8l138ru
IYUiPHrCfR1gZMxHJwGNDUqMsjQfiwQ/Cs4U+C3rAVs9/rikqYwywCiEbHem7HSO
OVRBiokqTF1YgYctBO15eXF7c0k0xWrbzZGfQVvpC/NJA3n4FhHI8q1OHUPa7IPy
eVCmspc/mpts7bgxo6cp+t8mD5+GTK3lYICKVpdAnURmWSFKrVrrr+5vxebAwnQv
ltZM2WK+BdiEoNhBAyOeR6j/Xp5v9mo6QVrrtqrB9jfGOmxu4MJjUpuloDEH47r1
n6aNiQwNEh4wICLJxtZOndYpn9RPxFpRyFqPFid6X4xMTE7oO/GmLy9TPJa1wEev
0KPYMESn0gn87JGast5i34Q7ZshPkNAHQmA0LsM97we3rTJBMBfOWOuD2z9Wk9U+
gL2q/Zd4VxfJ6+A3SdvZYR4AJVSxkN/eEQDndh5E0Vd/7IljCatPWTZSklLHfTDd
0j+zILaFXobqTF2T1CUdKt2fYfxUz25zoFO4W8sn4i9o/ChowZrZDbOBX8ZE63/E
acHre8r16PeMWe6Db8jF4YZkGOWF0jHKNq2Umw54z0s3PoY/CnpKko42Q3o2/O8T
qPslGya0c95vUw1MsECnD/i0skxQqDx26t1pVhOqlDlRX3W0vR9uzu+RYJ7D00Ag
wIGJ3bCRjeIomSVCaXqdTOCvFr9JCxfCiT7WyVfUYTFKYNxydEMvIkEjPS55gHIS
aFJDJg2lsc03Afj+FTB3Q9rz8WqAyorxcahIBKUUIIdOcoBvMopfWd+OJ4dPv0V8
JEK9VNuG6Yva4v/AojRxa2eGSgfluNrmzJOdH7oCVtYYAfseHyzPOrmXIfTtwpkL
qmuJHcpS7mrhSE4NkhyoRjdpLlsVh+hmaY4Pd3HCW3SUtTI3VuRGnv7iwF3a5jRO
nuisqWQes/Q9CCtmdbt0KvsEV5gvAxyQqjbRvS7krghqF38rRHLywl5sF9qLKLxZ
Xj23Y6ucYlUAJdM8KOglqEHHw4YK3k901fnqOXAnUlFcBHgNQhUPaq5t5B4mxVSY
TVUg0XB2QKFBxX/zpImtU7ZAQRLP/luDa0382jVg/NfYRuBKVz6DL74rLIwywkyX
68m+/cpeVlZdFT9jNwCohyvBuflRUlWL9arLVKw/SLuDevb/mC6m0NCvtFVePUmO
4/4zCQHQjavT4+/HvDMHzT8mCLqRO/Hhe9HeNL//XmWGV7X9Lbi8pNCGTORGKMSB
av/FZmlwuXSzBF+tEGo0UvfPtMNC4K8oArSLIP4t/U35MEY4/yCd4WLmWJJEtsvL
2rpek8XqMPxfj9wCn5mmQeB2/pfH1sZA/NZHKv92nqG2mllrqq9g0JgkP4r5ig1W
p4a0/0F+uN6f06wKpThNOy9k1hZ276h4ZhqOCwtKlbZ0sZNwgJV29mbpn7RYrYH9
42JQ6vfWuMHT44a0xO+VmlrOzGkNAwvI3lkaPp+SmPEqHSkj3UnVQrrJ7T1HKMdn
Qtf19UyJzw6qRstHkkv8lWVo/n01y6aPyqIw7QO7LSf6MnUi9kG1xjlDqeyk9XFp
zIZaUiE9eUHol1QOSI1XBXC8EP0uW2EFtgR224OntRJr51jUxH+7kwmsYw6ua8WO
PtZhxzY+OtawpafIYvAI/+/qeeFWkuIlhN85wKO2rqlzI1ZtbqaxeU04hJMbxw11
cmPhci4KOLXXHLB2TsNn8YoJbAhzN9YkuV00ptFyvIh+W37E8bcJ+k0QVxulf1ME
HhPXI4ScyEyACP8MIi31qAhqaZqGmpzw5uaSxmWYFXtRzNzAtcaRJch1FtGHU9fa
xFb06jMbKK8/2mMBW9ibE0qt7MEtXkBgl87oP8/RwJfNEot6ZKgZD+eaZoBEzNwN
LQrAGvfIbT5lEMZlbwPSBJRf0sQKJ1sRYYa9OdG29OEnsv6zFirSxkPszYi1rxFE
uYXTy3HoVcYVfnT1I86yYU5p0JNIdSbFhDhOirpYCLBvVUd7CyFkFEEve/gzDgHm
+Yups882/X08rdkOuweqxocuVvfw65qAo4VjDF3+oyMjwgXY3zF3Ha6jvVuEYtKz
ZqnfDcyp3Cn5Jh0J7EbFjFBBkFHfaDVupERfD36n77U9UxVsHChWzxwE6N0+WkPy
7xE/WVxjwSaUx1a46LxLWF4yeOKzvv9q8KgafUJ2ed71+jZCmUwHS3E2IgL5MRsT
q+dbmomP6JrUD7y+EjqUkEsD4+SpxMqPH96QKV5iQCRajSJc820Zg0EuPSP5X0Ux
OgIJuwoP0dAx249MMVT1fbue4Cjj7WvXDA/dcxEIaAO+bBQStaixXlHQadXODtv8
Q3sS1TXeLncGswMr+Irda+KiuTOkUwXQ/M4uDKAFeatBXDqDwtEyDofbVP3eZWqJ
WHdrdf4Bj9BSaNufdUl1EWlp+2vZJOGvVKXt5UA7XbR7bmN5Z9ybjJsEIvDGg3TZ
8jpEVjpEkjVDrQVMCjD8h2o1JwR3hEVu37I8UbvnJs3pcD/p5uHGL2FfWiq/epcJ
rljF6yEBNOrIQXj7GYrE+srxDGnJooDz0lPb+kng1qyPwXo2BZncegz3YHzR/THq
OilaascOdFJ/IdnyJn6LYAcApg29uGKjV1Qz6Lju3CUyoJVzfYyLNP2LR4hRgDhl
9hRqpW7Mc9tueG6ojv+mFolo68YF58eliO/yxbEg0I+Mbw4jwLXNpmMuBAzuV1gl
6rRnMXOaerTTz/O3BSwhfscDYxKmekNz8/s4ZMuezeTNLDTWjQn6KEI7Ms4UT17C
dwDMbo3sRenMzJrv/6LEqHKgpG2fkFguJ0fKSfVpVZBTsCxOvJZRqFkRun6vF3c+
jka9ATNeaenJlRsHM8A7WvSpn6sQ86A9FV+8NmVRbZSJrS2FpJJdN3NQjMXBY5yP
EsoaIpeknk8BvkshtLWCy+2teXJcIYEkqI7Gfurbw1RMMG6bbQIAUZ/lkGgl2lJS
RZ/By23IUVPjJj/xJw49tPkG07hEcYeHy1ZVp5td+LnYlUOb5Qw9gHtG5gPNFRrm
CSux6+2utSfmF/EI2xaUyxUrTLBjBLI44SvDRYGUv6gYWL5cNUjJ0Bg2SSd2wBpo
n90XAJqZGqqjsx/uPJYUEa7r5LfmB1BV1yatDjTE03R441HpvoAD8lzDb9Gv/Z2Y
CVDhAXfG7vLlGxJpo/p8JrRbLPs66xgb+hhvZXWJ3/9T/esqGN3JlzK7DyWzuPHf
YD4OFNnGewdyjh8s0LwFa/rqIsVXhsQunJ7TRE/MGRAnOXyhLr7cyLTR69X2Tdq1
1b9QcZEJ81f2ACFJIyP/DCMIJSz3djTicUbYKbGiI6w7R1NcjTcPNa9+bRpBknAo
Gyxr4ofIrlNHPNqE2RpgCgfrEe+YRmwk/RyUpi3GLsYCherc2lQxuyxtDotozVSB
LZpofTNXTG50w0GhdVP59hrz1qgIwrMjqOo122a5A5OKIzQtkAqlRGarLBhsJl8p
Mde5j4nrgk43VadCwDA6VhPZ/xlarh2cG0HvnH93E1ZtjdFEZnHScbKHlljf6f/t
1eCXt8ye0Xvo4F3tHsSQSbRnt/ultm15xWq/CM8yZidPVCBNEYrob891LHRY61Cb
3gZ48zlOJBQtrb+k0LSEa9sXSTxpSaBD+OdO9Ay0/Ns5Il9Okmk3JgaXZygtTASk
AODiywNhmSJsUNzlerwfYvkzyq96M8kW3QCObl1gETeIk0vVCF3fH03tbxdYsv1t
nEERlYljBK4CprFmdqwsuWuqn8ErKQIghPCQz/8b1otjzevhseVafNDyEoBiNHct
x33ifbzB0rzmUH0nmtpZ8f5fLqqUc0jaxIOwFiHveJ2YDEuJCtfjxGaFxLLasuFd
x2W113fuWbOiArjswXjxr4wLxzxd1fcfv8zYPDSU/XC6WdBMCA/18/cel1+WehMy
mBzTD2GKiQNagTjC0APGt2qLNW/8u1Lk0D4o9pb8TlShK7WK+nG9GbSy9mWKTaHV
KMnnTZLJIzQNPFoaSDZaGjIzroCvcDrMKPSX1i/jcwsOn/JYAAeF6qjpjLKZyyDW
5U9PK8mhacA/u/YMvuwkdgwugKyVftH8BKN3lgW6TwCsLTo+FdD59LQP3eyIZy5Z
gfL2Ax8km0HFs84M8r5onljDZP0SpGrQVemEEHc0S41pX3CGT7BerGFf+2e4+yWu
EtNT8p17eGKW1ntuOApqiKVPf0/NuVXit771EE/72hCteEYl3RsZ7IU5YdRkNdcO
ksflH/90kZmCSXJeULUbmyutdGZ60o2oDPlJDzkdDYncrcskwpPwdtRM2IfUOs8l
YjY/2KiaVM4rgBwqNSqZuuK3k5TOa1K7v3jFgh00yGqq7MNeDbLejsLZAXLcZVzw
n9bGHDuVRCE4MjIiNEqZYoEM28tpniFCeConmw1uv4ST+DGHvklkOkvhnmoRgWHZ
xvDZ2ULqo/C9kE1apRBPdrAULx6nxrxQm8f9OBjHL4RVekoQD/4FxoHN6E3Kp1jJ
4235U5JGJLcy5F95bEPHK2iBeyTgpqS3cu+tNspA+hIuePIcBNW8wsYMWjwzCtdj
zGhAYWP5HJhkoVAFEznHxpGkkHbdj4c59mTUFeXPmuYhEAFmlF4ActGrMDoSIcoi
8zyNSbWLzmp8U2kPMlXopOq6GUUQpD5QXgJqjm9+nvSR172iqb+K6CJ7Wf25wFWv
jRn1Vr5geYntXpVBlPl44G5u8Ldsw5GgrRnLPtm0qZutPZ8DQzQq5jAYQ4evbLNQ
BXW1TWkLZ03sLc79uWnQwRMmIErd1zY+lwydJoqAUfoMVticLOUuCYmeXH76s/OT
HWtxhWoUat56L1z3orGJEc8Ja/dkUACTRza+TjmJYrw0LWrxicV3BYUPz7/h5/NU
0Ph72qDzP/vvF2/fPex51iESynSvlYKJGeYrvC30ZX8VczdDHMqOfTGMgMcNP+dx
dJ8awqXlP0S9XSBPs2INDmWOa5LTJorgnTNtJjSpXjvoVdCF0CdRB/tp/U9aVzpF
8bI3ZOZjktQ6MX50R4CZAjX8MibzJ0jARU2LObXzzDEMnkDn3NN1ByNti4hunHBI
WtuakeB76ut3fJgHbi+8DPQsL/i6qnEt04GPFrC7cqnZMQAgcwLtedqEZ2XQ+aE1
d4A7Bsq/cowUINfHJWlOKoXsPIUL3vlpGe+sy1rsJfQmRhKfaVAyBjPECb6d/O94
q5ngh/qFtIDCnH9bnrL2p6eVMp/+hlDksZzdcGn1gQaBYP5PnjP1/mBXacw4kvE2
hZHGH9WFr9nMjerjvoXyWHXC7Mu67T4dv+xQRfl9dGSTgt68oFXNzPM/Vz1dj9Gb
WQBq1eHrGVzQPupoL6SbCsd3rfijURJESZgBRjxy0oDDKCbrewDfwZ928pNpw2yx
eoB0InXba/384UegNjE0dfHWVA7RPDjQWh5gsbLPVs3iikUYHNVGx6D/l/7Yf2wo
xSiy1yvwY2NFy0rT2MHLWkbeCvExEpXzDmmMyfMtqhhjbHasK00DqL1D4EgjrUse
LVNbDsju08dJgtcEMVAk3I+pHjjzZqZjytt5OjraCFxcTRUMXETR20lRZRRBuJGy
nbVAf4FDVp0nVXM9AXAntAVOhN4XFMf4r00whhoh2omS3DCeAVNFnR8px2skg9dn
zLyB9uOJ9Q5NrekuWV+2T+ZIrxw1h6VXCwf8juCG1AR18d/l67OTkBbGFiTeZ9ua
PimT0z+J8T6fKZjVEQN5byj5I+5K0KFMOWMoN0RIV1mjRlMespS5pHYVWB2babff
rxAGF+Ylp7Poh6JFFaquR1MH+JlgaWM9xJtJyb6OwQR05kLQ7N1mNgz2zo4K+Wu2
4iE8yC8zMnJpbiMmyWDTqAG3c6opPN6xLRYc77YPFXre1FDSb6EZ5Xo2fs+lsOew
9ItFABsYKFmOEYEG0AfX4nXuSZWvRmFNVh0rgvALJaFrPwYoW9KHFxh0EwiorQDy
OuCD4xPxN4EF+4hIPwSgIbQletEvjDFPCTSEdR1ls0qk5YDP21Zn8FVi8JwIdKBN
i6Nnw1NXsS+6lixQGhVkOVsQUufUzpr+/xjZVXH/S1nVsbqqinrDSy0hQcPitEvP
unGSuNjblEbxgUrqmc0PzqOnLKUMq6wQ3CvVnNl2VdIIZT4ukM9o4/U99tqEu0J4
+1cdSOBW97vUQpALnP1V1wUfeOOe9IGzNulnPwquixigKqKkmuHw5R8W/vvi/qBt
tvvsqhaxGo1inxkUfyfuWrn/mwsop3LG2ccNKgtifKAmVOCf/g5ufBLqudhnrvZx
XEJfpOK6/lUfrB1QWWKE/w3fFp0tKPnKUkPrfCmCGK1hk1s94PgUJma+MOkmh2K0
/n/MczgbRrZ6/iazsrvaWk3VJvvsOIjc72SPgxBHGSYykMC67nvkFbuctdPJurhb
RqMd9m3nlh0fvaVViZ4CJMurN37iW/ZrX/r/A3z0M1U32qLaqYNNDd9iNdpzOSVY
cQ/61Kh7wb9sZvkG5WJ+AkBN9vJE8VRjIpz8reGPiQq95wWwTRxZo304pGGPaBRb
sY7N5zNaxjpl9VVocP3zlv7O07qgWrDDWfVIzXxRjZyWfrcmS+jmesKOiNaXSvco
IYKVFw1WiGLbR8Hf8ufSrZnWlTLqumdJrFOX8/Tr3sB2Renp7FQmFhuECDOAmbI7
2A50+MF3UMyVidb+9yzfYxt3O+CWyuXmjGcwAQ09fzipZKt8aeA8RdBwIpgYzUVw
xU2K0gdtOsxODLRdWgH20cDfOf46kg9Lu1XZKNIifqdYIJG2tYowKiyeLoBIDgmP
9wDC7QB77qrpZEYurvKeEEI6E0Uf3nERgZ1kZWFDnKIHe9hBRokER+8APgOaVLfO
huaA5wI3beKRnnr7fwvJ4CHt7tbMNZJiyap5ZSH/Ed6EYFIxIAi0QoDrH9ozjsxo
pyfSTMTaO4/BMat7hbh6M3crdfPZODq2dgXoSCkZ4jkDqnqI7cMHbQB3tlloZkG9
No36UHEWIyqV7BTwFDuHw73gBD57nUKzzhsv13U0FHUdl2NgNdKYnlfSSP/0wiIy
KaEPCXKInOLlC8nLawuDVDlsLWiZrrMe08nqx6h6C4LJGuhUcODC+CmPE0XPDTf6
Qd2W0fTCesdmd6Y7fC3tD5Jt9VtSSsN3gQKr2NGojlL4dyIba5nMDvYXVbUA+IrT
l3i0fkRmJ1i0X0ikhuPKfl7cDYhijvzXFFIySkyCgbaIXbhoA7GD6bks/lhaRB3k
UOrqi76qZFFRr8AQYfeEmaXio1bcoReuMMKyqCLEJkXpa67Xnc/pypvIfFPtwcpR
zOgFZ8PImd66WX7Xe2oTYzBsjtT6qJmay5+FeI/4msxL6NRGR+/DKJzwQTk/yPnG
FmJKa2PK9rFB0QWo3sxLsH2emp+vfAq7PzOWDvWKEDaVQgsDcf0uoM8TSM4PruSz
10adKcz97UG3brcluoPPmSL8T7LSSxVdd34lrhSrp4sDybMteQ8/qnb0/sVBOjT4
CyBiSqinj8jgG3qFzolj41dIVRdvEqcBIxKGCWAp/LaVf32JV9pG94Le+tHM7n38
vsbOdiHBsq8OtRasORlrQXBfH0q2cT9Hs0pQaeEMtglPVWuYJ2pMWCPkL0fNVd2/
lDHZ15Ihz7NGXimbj8klfy3QwJzNIdK1lf5A5z9NYYKI6EDbSTm+EGpmOoldvwIw
l68cYcrrth+Cdsp8YSEF9DhAXP7C9pZRj7do5Sy1R2Jxhoze18FUT0r2j7yT6W5w
TCQaWNIcQeWVkweR7RbeNrRXnKoBKQNVMsG4ZUfS1IgzHreawOY5V9IydH1Rnw8J
Mu8j6cI9hf2Irdef8R7X1QH3tyRMvI2pqsUlAbgWGyjlOX/1APhkKZERVhWiYu8M
wU9Hioc2kRHChRg4Lk/IQIOfvkC3oHxV/TbIOGLGC8CgRMpwiF8xE5OnDDGH23bQ
xVTjWWjvGj0OGoH/Mr08tV8+U8hmlGTjEo88V/2kqeY47Gg34jkhb8Pjih2vXDbH
xu5XW4NxtVTa0fJ7GTghqxZsZq06UmzzJRwbQPTosTXVNWpO7bBhdNoRlp+GFQQc
eQUkcXMi2TggQV5YOYvUdriicT7XolwXuuAnu/H6x8Jw7COFwbJNWcsktJDZNQYu
g60e6x/KZgiefZK9COD/7Cw+A8twr8kzRVMoMOtI6udxrzrVwa1lJSdyAjEC27zM
JCEL4Pe2uYGPgeDLp2qf4lb2AIiioZvdz4rM5ilukxJPYVPHbN78FK3k6DF1OjEo
lZrpd1PhEILWSOH5jYk28o3Mgf3QdpSggiqq77Z7dcFGMyxxQgE5kpwODBjWZBoH
kXMRKZYs/elzlFqAZtx0ms9fiu77Wcz3nFWxTqsIhNZzuburC/LY2gUpvPKUkBSz
hEq8qJpvFFWfte/rHsm6IiPxaStVstH0xDr/mwPbSokDe5+DDDneBa39xkAx9P+t
5kEkTIKU0zJ6T2dazS7hc8JwdoMpPsU1e2t32S6UIcCPINZHkTxs1/pCixAUENb7
8kVEqLqCAshrPIfkRU86Gulrc+0A6BewS/GH119RySkMIVFb4Qud2ilWP80Sh5j6
C2m0L3B/rwguGJvJAn47aswkHjT90w1v6zfsI8pJR1lsSm7aLIgYjYLAYLq6aBbv
QFsjrwinbgCLhyVG5NUUpiTuQ5hHzzhaKbVaJtMdi+5S6L14UBL2JInrvm0DR2N5
o4yexXsA18KJx5V/P7tbqntCl+5ONpiT2q4XuDPk0D28iGAns+t3yU/+y07ziMI3
rAV3+jIQSLLdy1Lkp6PYVtK1XoETTQJtr7PG3bXC8HXA9eiJ/DLa0k2LQdmbEe2z
bLSnNzbog3fXz9l4BYpyVg4E54j6uradIRhj0Mr9jNLf/1DFk7Q4tGBk0LHyiufL
NVpCGXkFeI7BmZu6BXSPOJmNROnv3sngRPMNccWj7+OTDtGRNIZ3aSefq2qcJfoP
ImhFBcHSVRG+xmVLHwgViscMPrHhT/Z8YjSlIO+0uH8WztucC4k6/JTcr6nBppOA
Rwj93XicqW7RRAwaTJpunO/ER2cUgQwRUibwbGxPlnpwE5sdD48u+WMke6ELWfpn
FcKuw35tlmwJJKKqxlaPbkR+9dwVS2arSyTlyIOaD0E6PehIab4GHOawweBMJnSf
A57UpgONXkqTOu5Uo2lTL01YTHp8VPQPpcIpzkb7bq63tAJlO8OQrsTQe0yTchpR
s1o0dwatUrd3YrAtrRQ/0yuwdeQNZfD+0QDn/nwZ2O02n+zxvOJoVsm7VuX6Lpv3
y6w+4QWBjmQGusbqkkVWsJ47QM5VgU2UfRi/Kfy6u9WWPOKhcl7vfie4CWe22gAQ
08nRC/wn07jlQAnx8KhP/nr+6ZgHOwxtEDD5m22Dty0w0tdkqXZ9aj5/M+L+NsqI
iN7Noci4EimXWNYArUs4Di53BtpEzHhFYY8gO0UtxeBtyX3wBubqaHNADoL3VwvY
/FqotbLT3g1TrM7vpnhaVeQzhGrRb+6G20/r5EQbJKGW6wZXNFq22n0Xj7zMa6j8
hHhxA9t2T3itL7KZ+yFLJ5Juj+StgEuYxD5vzvmM26uRZv8EeHS/umTvep/Gcyo4
Cm+MP9p5aKGekJ5LphyBtSGs07n8TANIzXoMdu6pXqWwot/A0npLvfP5jCULWAXC
iZO5tz9YQ0a0g8g/J7Wytn6klJFjsi/62evbcGvUU4+C2r9R5ztLM1dwKX7ctf4g
vTky99vp2FzG4S75FObCpBavF4iSvjqHGF0GicJGnLKB/72Jq+t222sxDYLXvQDn
NK+GSB/xrGmuT7OGhT3f/eMb31T78KLYgtuIxd5t/dolMmu+StA8Q/Bcc1SFACnS
QTchBO/c6t4eCAfMA6eYp6xyfI1XPIGGniN64NMe7l4xQFc459pPXoItrPuIIcpU
scOO+M/PHr0CMaNVlrsnBg08UlhMSP3yZv+g723BOOsjcRp5jUcZMrY8cZJRKRAE
SUil0g0+xHiFPoMjJ9hOZvNvAUg2+9kRjXykyfFzfgzlXH7279YlD49s6vQ1QO8P
dG2isOBqd312G01MUfJUPEj3oc01NOKFlPNJ/I/hAUMOxmhwchZRao5tOzQwiz65
VkrhyE6fU88AumANeu9u0VvfRxJ98WfI5iCnI9VUrZ1kekZUVDpfTJvQEk39MGrf
94vZvTpJJJdCse981lNRowd/bMjC6HRgIkrOadBM/6jayb8okPZgSXsJkZRYcL0A
HFIuLqHnfL3+T69vvkdQzeHmB3pH2mxF3aeF70Ak83DfajicZR43P6JDCmpuq6yd
lW3W5CUtQZ/I1rOkLer88TDWKZcoavZhAlImmmEhzH2iyBmSu9N9NsLxhXhDL3/h
LHWfLWlp0iq3VVv1QHbbYTTEDMiPHqeDo3iRcsCJSRupCsBgmRmDE062FZ6AJn7+
dq2yLVlt4FIcxFJtfzUnONj4MvYQw3JHxYdXntWX3NZUNpTJwXqdlf7QoQmTf0jD
ioLnW21NqFvBdnHoWrxUqp+/kyrqd7ccsBMU1nfkAQeI2quH3eMNj8S/F6BKQdEb
n8WQ9wyuUnC5nHqlM1BDhjvGxHTyul9e0/GgCxig4S0N2AxQ06pb3pfXQW6cQ8Tg
g/us2jH18+k3fe3Q96FGORq2z3kICitGylkoY8/n3OwOwSCDiYotNZU5/dw3jPx8
vdB8FfzyVOK54Y7JldYMAVpoxpy3xHQdDUM0W1/WgnDaCOEGvKEpq/CWClqm76mE
15B0tiwAMn4qclnti9q8ddlfAZy/O0f4TR+WyV/A4B4sLUmJB04GDjlgvGHNbNCC
diZIUC6qbVSKIq1peoe1skdAMrJ6ecbQR+qSRdLZN6CLWj6+oB6PGF2AbmMbhczM
RpmgHftQY6Xn0LumHSZRavDzVLyDRclWxTp2fL/zKbLFK0tlbLLthJPIBPjXAP06
aINq/evhJ3rnCAGv/CB3STFl7v6cNemTzgRoonWdl8eewyxMcrRcG8acStMhP/4w
F20r8LGaBnXsBm8bIOVrb6IRfE5gKao/uGZ/I3GbeouVrzDvx6BQXfxUM7mdkj9Y
w8ed60+phetG8OuTBnf+3ELhzwFFQje8qy2fPOEtxTjgHngiNaOJE7cpGVmKXYmx
BorWLUI1YRi9LSWnKfDC43EhPUgGvmjufN+XkHr9Kk7n2aa7y7IP8533Asa/Q3Sh
5zsSOXFqyW1INM5CWHmm7iOmEsp0b9L9QT0JlW4Ugc9JYBrsCIYa5eaioKA4MI4E
s2k+6LfAZsGlKZwN42KqnB6Vt4J+DUL4AT3tgCPdCbwzc6/t10jL0XLW5UHaswAR
mNjATJAsA5Z8buWfsV9L6LgZAxuq5NDXl1KDMfbZI1YpEGt6YZS3m7QRda0IBw85
MbggZVg7x3mQNuK5t90ZHwtsFbP2R8IxKyPWLGavPB6N5v8ldV09M4m48dcpe1FS
X9lHmwFQLYF+1LhpnmMXsPrk/rGqHS550IgEGQAVEmzZvqZRV141rrpXZwOtriSp
koP0/bUPJxQhIjcle+nd8J7MFArWX89CVsGpk/CFkCh/Xo1KJiaP8ZGU1/rqIxNw
rGJAmT7hyxLX8yPi3xj4WcP/ki83ILO9yPasmkgZF+N5xllmCTWl/hAYqeAbGHRl
1VN1SUxCKNsNXs+d5XhZdxvYauvR15PRciMw7e8L9mGDVH9ODGzIDmpfBSDw34H0
bCoW/Yl+Verg4Uis9dPLKGCKraqPgxYDmMPZIlyOoqXXtCGnMyLzoLZk9iXlJp2c
IM7ZD3pAy4qdNRhm5dQ+eUD6fivNFhhWE0DEdubNTyr8ObkT34d7lHvtfAFy4uB8
p/TGRKg3ME8CmulU5hKZv/BY/liH9IL8AlQYbJLsIN3x9x8Ah8LPrnuaFh/2UAYz
DVRUwkqpelTa7z4SvI9Vvqv0rv/Nifz0fLhLe7u3oA8rki90WKRkxYUhWP4WazhE
apgZTDkEz3k2yNmwME3txAmgzC1OCWNT3/NzfyBU4RK8pKpfUBsuonZedrb0Ls7E
wC+dvaQnqkXmDONHxHfGvShwQUaRV/Jd+YWscXjORB7qCZ/xPtFk6HAYN1OquuB0
W4/l6ZwHWXcKtPoJzhfK8vEI4Z2s0ssATTkmBpAwuPcC2bp6Y9XCtvCdI4LZ9AHv
63Jpyc8NykGTnNVBpG2rWCUdwb865mmp+S/M/vFYKbsuPlFqM+FoDQ5GxWY40Lng
N70HeYHm4uh3po9BMS+zrpe7J4JsMRYSHPaeqh5bm/yQviMNZv6S9VpVjmUoODy/
u4U5hah+2+gUB8hPiFM6lj9o25rBIUfNiNHabRxJY08Lnd2gllc6kWdpYnvd3dg/
LOBDmi5VHMyvftM4vWDgckNh1PHY2Dmc5yJhVZL2y1Yh9xf0Ep87vo1iTy+9Sfug
s4WRIM8xRtC7PyBQTxPxHgY4+l3E90SU7+k8W9ZZ4wDKXVK8aDFneyMSYz8BOJdb
/AKA3LpV17rpgEahMfOAOIqdXIxqNaRBjZnzCKDGvR2jWCjn0EJE13BUuyiF7Znz
vrI1gqMDb4KFHfin8EyZE9TuN4p5bZagqhz/aEvZnbrpguxs6KVgBcC5N1DUsQKS
lUbkE1QNbheHEpjBPrNwXzEZpOpWK7IyPcskRxmyniQQT4JwElIlTneKI3y+x+g3
AbYKgrQugaHDkRbTklWe+BxUCm/0+nEwPIueVkH1nE6bYGKw2n2YW7biZgZj/pe4
seNKM4BSNU4vvzf8uYWKf9F/ZUyMAPw1Vniaxn9ADbddDlJUNQ6G1T5wBq2A09r9
75+I63rStioKpYSlYaGXaNheqzDoiOsGHw0YnB+wm6C62N+bz5c6sUyvC9ZW9f5L
PNWMkBEpLU6xIq0Awj47TfKU+/wwRY9pc8ZXnWdOlczbDQSAN3vioLMdhWJgvI0c
7sbpfVGFquJ55nJV/c4xii5eDXIGkvjnHAJhw5pQ4st1BxB2uKab6jgdKIxHwQTn
4GK60BQt7egPoU2eXugcwBptNXwz1pip9jdjOsrUH2Ptx1V99N0hqoF4FLNusnWF
qIvfeJb4H5WGHtU3qFMVMjsKN18i22z69NwHtG/sqjclAecTADbxi8kX6sLMqtEF
NGbt6FNPfYlVsCLA+SEtfXT4XXOtFaZqlY0id7ZJbiyL7FVfdRTRpFlfA9Xug591
Ibh0Etsey2GmEUMeoLY28dTJn3D2xcpM+lhWLJTEW7Xp1z5L4jb6avJSBDdmT156
GUxwLaDpM4XxcW3agOK4T5ayIQHn3De8aNGE1E7RQi5cHVF8jddear7M6Nr09jYN
8geaerVPuVqcb7IKsQA5tfA9lJyYvvKQo8Su76TLXYPG619P4Pec4mYKGscrj43e
KTM4DzGhkYg0RPYcS2pW6lIKszMbDTmbkfjfG9OC0Pv4OGHxcfarvplbb4qSkImH
OBUXqahUb7UbjyHPCrV3kKZb/M35+xqy3a1O4iN1nQDNjUQyG78pGbijphZA2ucc
O/CYGSPf4ar8xR2D79bIjDvyRujxK03cCJ0AUHoxUyRGJls9E/MHevnRdLxUAAbB
sxZ7fsGviOXuOFFQiHy93USLKaxOOd0okm4neD6BLGqGCzP7eJtQwRmH46KTprru
iW6RaP3r+0apJZ/veW0WPOsQrd4UPH9o2/YIAZuRMneVqXjR+FI42bT00GifGyzK
k6TOZVEcTJj1zt2uSKFdXYByI0Dhj8cfujesfy5EpkmpsOSommcA+9+AoeWaf9ld
eOJU0xZkosKVJlcEB8L9D7sRbpkYOIaqeuL9tyxKHVyemlJ0ZUp25C4GJbOsV2zg
C10i66dj/qcnT0PT7JJ8OhvVGUN6u1cs9Q5VwSBN3OikacC1QP+/0jMuw9wCSjaj
27ik1qJSfcmF1M7vAZon3H1q34ObATcedRR6VDS81Rbk6jo2egS3I4DVp2GwYukZ
H2uc/59RYy48Z7VkIcDEbvhczD6RxZJKXEv+I7aj6E4pUVqnIJ3TrQk/oOeZ7Bv7
C0frAA0k8fMWwWG6sSaQsp6H4VortZtZo1Mxe8KYIFW1uUz5e6bIwY1q88/GwZVB
uIsXV0lqZD5vhPEhFlyeNJ+20iNDSxvErujlPDMT6Z8nwSOsZMrR1s8Fk/QU029D
66ho351fLzSqHlvF2H/MMWSKc5W3+tO6Bl64Vu1xmCkr6egOjV1kga+txm3HBh26
MHPQItaUeFa+colXPBG5Rm41uX3HKE87SrB81H32e+SsFCLaZ7NORFpJKsfHNUjg
W4EVjDPbx7aISqpgQHd6W+B3Sd+IbFixCa3B7xwNC8li0VTCxQN8ZuOFSMgrEyLT
VfS3FHLBqbN0XfsThZzShEoeZaL5kLTOw12M2BPBQ5iFO2lttUFKUM+EivEcIYw4
Z0P3RCH2vOD1RciZEdlv2062NjWaz0WJ7+X02YCtEWONowyB+FLVuLRxmvahkwQE
BIsQtNifucowRAP0rZaSIzqWz9QQfqappqBLcLTaKO3z0PxCqkhFebpdjVFRFmVL
1qhf/5XbpjBPyLOtmcnKCuBW+ibA32Zsqc9drLL82EgE9m7dh/PigvvmFN7sv6GM
RljOidHBCINnV92+pZctn602UlqNeaIOJ6/Fe+y/TxO7Ac6aiQbwVEeTOZwe0idj
hbMc4Arbf1pigBtsdbpQjJPNLolE1lquVSBjgq7hrk+B6eBVOJLfiyLZOHGl2dtH
wmJg/Dm9k5O3o8PcdTz7ajHSPug6w3zOjwXoymMwtj5iWlM3FwyJNWJ7POEJznLE
NFLX8TKyVgtA/hTuQsU/utzoZuhooYcAfIMIayfL5zwbqTzTT3g1+ps8l4QSj8Ec
7h5jsqpji3AjE5P1latARd6BFrSwoyqnh+sNsTlkxstFdjnt7LAFLBNZVhoSDVay
ZX5xeU1m9gJRAyOFoPF13a4HrUeGaFUsueWcmCNBfN1v6kfh3MkjsqfT/S7WrlXV
q5Z123uSQKYy8Em7zT2EKEle34hzMaFQqoqY1H1TVJ49t/n0BCgi6SfOrxSjLX+A
slxnKJfv1Car0pAn99HtWYnawnvbxkD3XHL0yAvRtcgQRAksF7A/8yVSbo+RAhTS
AqeUuXEPziddX9v9tuLftjq1CITczOx92ngcLQL0IVRrYzY4dyQpJhzWPhZZiDpc
UW3gMZ7gKTW7GookLOjy4yytS6tQ/U8rZYB0pmVGI0Q4Cz1eBHg1QP8fWCCry8z+
D3ou9TKkD1wdkSEzhFGWQeE5sRGf1UboyxhjW7v2Js43ee6eCNdxqf8jr294OI19
GHe7+Tl3WMnE8JU20TjwVf2cICZbh2Kbim5nPzauALV536KJdzn5VIWp8nT1AMuw
5m2y33hXASiWDWd5pzMRSi74fDDzUj4PQLNS2iizCCbGKOiUMylBFJo+BJfqAa99
7Zxdy5FoDvgK/Z4SiTglH79N29xpQ8zn7YhUmtK+09WrP8IyueraV2TrOVo93zPA
9lL5ZxsF2/iYwyeyqwHe8XLfsEIk6gWCENZ2+exzt5bCigIOhSEXMG1YRgyZO4Tr
nC2JsBiIQ0Nlr9GZHFzP4Czu7dd9i1jp14u7RKYyAOv3nSYWyA27pyeRnxOV4Xuy
yu2FM9fpb9Uc1OI81TKrAAcnhtyqL1AcDsJBMOyYBOJk/Squp7aneFGAaV8YwT+q
TIE+NB7fe2pHiaqP5Rwz0dii2BT7dMqFD0MSzxHn5F7iOeJ+Ujt2K1F6jt+JeVsQ
52uEjUUv/6HGMMlQOFVeB6Yt4hWV8RkZx0ClEmKgtZ6akycvVC9TWSI73ZXOSI4N
ScmeK9UkakbqJ87yofVaDHZRzrMIbuU0upf+YU4MTRnihumBFGi3UZoLNiGmuAj+
NlpWdr11FS379CNxcABEGNwnmrbfJLutjU6BCUJgD7b5OVfho9SyrP6l6pDAj1Cu
8opdp1EcVlAawMRgs/bYVpEqL/sS0lPAmWhKXIPsX2At85PpwED41IL41WXqFD0H
/51HVGdhehHkk4+3N3aUYx4+ijF0kN2tCo1WbJTl/8ZQtjj1W+3SU8sonMZgX12i
qWeYiLLO3Km4SsuoqtFEGmlLdJt7LlfAXmm/wnVLRd000t1DNneGbSAFOzfgEAUf
9f+RIlf3S3fWH+I3/alw/pJadlYD/dGoSeryGLuFHn1kxjJ2m59Frd6nAQ+Ushnb
nHXVsSHYakmxOxhdA8OrRd6FdgJjHPWA9LRoZ/WqUGyq6CgSScAHQcRpP4FVU7Tw
XZZvJFYQ21btHQp9So1z3EEalXlhXwCOpQuTD1x64GOZRN+RvwnqsZvseOmksi3i
2Nf9uzGvECsYxvF3gyuHlj/Y3qRajKmz4PGtNi3DBOmd2oZU1w+5swBd0cbXdlNJ
b9SpMNpTolm9gX7SQyrjZhMTyo46cwj0W/w1BFxhb5b8xQO14w47Z1pcSvN2TNmW
shhMAe+oQn+Jny+Oz4RI34zHzus/QYvtV/sHHEoXa2hghGLYGV/KKFZ66BL8TGfN
naPXMP1x921VFsoGTcz5xUZ3JbirZhn+u43Di/PIZ5WOtz4xAiPL3G72ZM6r5t50
b4bnvrVEuIpWAfMI5BJBrH45X0T5OCJhKKKIgiyr0HPAW/GH24ZLnLw7Oa8TH+Ju
smzdKuYrEGeEKWWawN154tGg+q5sqDTz+diRGpfvHo8LNcKL0CEq63/IRkDuzQPy
o/FbVfoVrzuAAdGwErGOuns+KqAVuuj9pKExEZYob+OjIUEm51Ok9W+2UOQFdPf+
CL25YSnTxdimnbqrKZqq6FeJUtpy8ycYyNmoUdXIw3QgrOtoP/pOEwaEE7seGIis
XfDuYonj1bSlM/7NC6nW6eN9KnfW5fLjur0cwEABmwdL2QwEu41cdNau/iGifM0k
RJ5/+n3ojs9b2bracDG1I/h4MdQ6R3dio0yYULiVu7mpVdxnHBzZac5toOXokIWR
49tygoYMwjG9+QljOziCY9kQwbaZkDxOsNu5EeDu3lV+YsyS0G8+Uiq6rKrGr/H/
pxQHaqSrliq8IhpT8H0rGOypBIdk01ev/YiCtNhYBwcjR1SiwPi2VqRFr3ubj4mO
fCdYKfnZEvtjCjp6ZJFWRDIa+iul1ZV6od0Xl6bmZrwYow8CwYhORUi7r30LpmDy
nkYrwdiEIWq0mWoT3Ukd4lW9lwgMtO8f3NsXmplrtktQzYcoFPztP5985JzqDVFe
o7ec7MSDR6mZwH8aGjhaEGx1ZqnAWoEdf6OojN9+yMVtLkAaTuFa8qX842HORCkq
nw3hoA7I8vofJuAIVSY9n0/FMv3hBx9jN6G+3F7APYkXHaCZbX+z5Wzs4oaz0/ue
o9tV5Vhk0iuTQ5FC70lVQ8GLI29X53rtehYRnH9hA1HxrPzUFRlNvOJeCa9W4UP6
giiTAp3cEHXldxLdbRL4fnXV4v8SW6knC2SHs/4zCT81jYFevouUoJOU6Smx0diz
fQ2o8n1IvslEuA49GiGkFH4jPRPusZvT/SxLo9cxv6STrtNZJW/P+n8K88H+5U+4
2EaMAitwnIneOo+Bs9znAVQrBwPtV0H+Wh2dffsNZ4gTMDQvS61MztHw6brhW09t
H2Pv2wDNjLlOBM4Bkc/EZKXS9fJq9dxPAAoIXsQkneRDc7KKjU6QBLAvyE7Oz9+S
za1LK5V0MYrMnm1ve/sjy9ExSI6Gegd/3P/Sfih5WzWh7CTaYWzaA9AOXGt90yq6
ql6jSg9G8RX9SjZZ08BE8hygmPRCpEJgyVVonlgFRfN8bBRFzze+lROcKNeXt4a3
rPhsysPdeKDnfHIvDKheiwGn4JdU+jwoPjkNtqb870CEphyhaZDoxI9m8/d63OH/
MSt2JTKfs8MXwvOFymTbWgVsQvbx8j8sWlBwHN0Zt8yLy5D6Rl9dGJfJusW+Uy4M
pMLssnPXh2UuLZyxYK+sY3rzrKQGiboJ8Ku4cblTlVFaH6RS3tI+XxuJLQnOimVN
8BJWmsP5XvuTU6wcen/Cd1HiMjoIAFPzLZ5uSh3xgmeKbtG6v8Q+6dIgdEsuQfz6
rDMbG0as2BRAYdmoHbySENVS9B7Bu8G0BZYx5DvS9wionFTLwGji9TAmN8cYIo/q
uLFstwVkWo9V2rtRkk2gwq1uly4XuX92Ruq7+oEtZ2neycIwqLNZ64SrUvE+41FC
dZ4h3eojfE5r5e0DIhK/E5y5wGoPOTpDfzo9SkAn/Z7ctKk8oMK2x/8HMWgF7wLq
MpC/FssJ+NR9vIKAX4fiGrJXe29DZmM4o8Wd+IL3HChcBkNYzhc6auB9BUCyNDc9
nJDZcFF+dp196lvlrMkSKtv6L3AffndSGd9sGQ2GuGYKUc44rgUMU1DXqwoZs4OI
jOFtJXm1Pp67kfLyIOpprD5DyYZyIjaBHxQrA8vf88dxCkpKsipdM3i+BKyPv1OD
fyB7/WGUVraqlBJHCTf68v9msq4Sv5UpdbZGl/RhB4y4LqUH96wA7Q1+NMseUWi3
2i3717cegW8FzKhAowwhS5Ck8d3Td5/fnBLBMRuhm/SY7//sQiuIL48oIzUtBlOy
lDQ795Yq72J/rHF0KPZxy3bVcirxsQLP05STivVN4Za/5LRzQLTfbvkKz3cZ0ebp
zyUls6CzKzMbI8iMaD6T+NVsCZLzC/BRLyJu5EXWqUes3XvfCMGd2NMTj8w8VtqV
srwStofbBcMKW9R/CtknSXXLSfAm8eynGUhAMkUBXgQ8MmiZlGYIfN1+33mdrjah
0HidFCQCRPyly0UnKVjj1Zzayv1SQlC331krtphjrxvlE60SezF/2k1tznD7+MPz
NSfN14vHcVeOnqhvGSv10dy7+L4wygifBDGLW3mEZsXZXIIrZhZTc3y1feAiMFKV
Fg6kd6/aJmAYXsENVx0v0qopHpqwZ0scZD7yKpJbG96BBQv2AvZJberxsnnUeHe4
zpEMlfWNVi3gol8jOjhHfZhl0rjDiql0Fqouv0bk4tRV//rYzrAQxoP7cUbAq8oG
6el3+dmuFc25JmEgzRAvE/hpi+zFtjtqIgw9ELhBhQLSb3OVxALTMCMZWqhlsMGH
+E1j1vznPRlTKci+wExAaGLtzECzGxb3zyuPFRFI2BabiHiSglCjm35yK8qD237W
m0rc1EOUneQ8pnOE058n2QkShOZeJxQtCJATE2bzdBJCkQ+PUAjZNXvEhkrPxBEc
GGuYAr/LkCck4RWNyioDZwlbdsG5Oq4u8CXTzpf0+y8E0D/uIhOeHe5gtm6d1jh+
sQrsbKMGlxqUatcX6dIsHZXzxZOQo/eUw36z9a+56aD0z2Z60EegzXzXNzpNGcRp
Q+KGim3chfbBsllUVpGK01EExBDL7lN60PQ4djygeuggISz0sZ6LIkif0PiwCqX9
c+HVA0CNZdzl/IyIZBVoLlNNl7AXPaDAqPogb8GEiYXz9mDxsfWJdN6/m2Yr2oR8
virNNQ/J6wifaq99n5s9XR+gmAjwTPXzuvmQ4C6PQMLMuf5POWOgIlbfbRC4WCXm
UHkAZpsHPZ4HdZps37RiWmC+5tvqaIESRH8RoH1c/FO3/TgpD8uZFZ4RSF/Ztg5e
LEEK3RoLiD/kYzTZAhvdGC5NltnhMC1In50Ygy6uU8z7Z06kYAo7ByvH4KsdAYdE
g0A/uNP9zUKT5ILmKnVpRNLlPU7yW2IaIzY+H+fN3+ymh6GJ8GlCqkuYavd1gh5Q
a2ZkqKkkL5XG+Cv+zaW8Hh3RyhXlJxVcpc8MNUDtE329EUp8bjOCiPpkt5gHuo2k
wgtGslhLcFJB1hz29A/xgUQljPYR2qVNccuHzzfZdICnGq0uDJA5wxzxHST+98Ke
1WGUpd2nnjpCIt6eXAkMwfGn+nwJEYC/4hjpd4wZpzhFhOGBE0OwX9UqcHrLQvQb
v+Y9tFsvnknweb/brIE07oLEADgRGn66g9UvJlS9Z9sZLKJC6o5uo/xrMMi+0bKf
benwqaWbqlg6pCxupqg1Cdw4DzncQ55PRxO2zT4KzWluEPPGtcIFBQYeE9TQ8bHa
X2tI53tHs6x0OOtCkKqDrDYSuXLtBzK+h84cMgrsK6Uwgp0Tm/NqPl6qCwW8tpwp
VOzypBiD3K+rcx5CRlZdVlgN8tLCHyItd4tBR84Y5Y6H76RQIcDJHng5rmrXXy3Q
TfL4YjYpi5X1GABUokzy9UfAf+bmpoGmyCE3AetBoS7BwSSfydh7NaOu6+O1+QsD
ailAiaG5VmcMOAlim2emCCMqSpZZE1LNTyTs9f9RInq0t0Ny+/AdCRAHwXvksdrL
KqVCmGczIdRF+CsTjkslUM9ADLSGKUioloMlnihUBwRPTUou4DD9nVXt25bsNeUl
81FdnIUqFkGqZd0ge50WmVqrNKDu1mWzFRXN9cMhGb8Ybo1eEffTIdiEXQOBtJ7i
B3QocO4zuhpN1iWvJCdPxiumRMQTNTwrKCTJpnMgEon6DmM8QCWM+PVk426NibNl
v3WCN/eW+GMeU47aFa4WeShkrT7ROKGH8RY+oMA88O+b3MYqQIvgdko3QYh13Z/g
Kuxn0ztp6MjPlKetvN0RYqOTKNVLx2qw88V7w8LT/1WE194Wh6BPvzewMfy1yhkt
wXPLTivKxIZ9IOn4tCI1ShxMLlougF+M2zqadSZ48wRW0eQNvSi24rr2DT8hQF29
jZyWvGudVy1yhFgjBqqyEtOLbF2u/LYP3pV6wvLltKT1QGQgNCvODd/M6B6t/X5a
Z1x5s1oH3eFwOt9SjMJF9wJlmQQfaPEmf6MJ5LiYIjMKdVMyBfvAPcKDAc/miIXH
qQDafBX0A8U7EEuRJ0moPl0Dl2vIA1Kq6Xs5g2BOfLpM7JEXnhPWQHQlxKlcvA/T
BdAUXaUeSTDiaYHuRHkDKyKMrDWfAVPnksaM/P7RuxnjFXNmPGyAKesgO65vqzA9
7Ohu1SDkqn93IiXI22BHVL09MSgeV2P9gqrXTaPVTPp7aPTwjeuDPao0zVwud318
jVUAfaNaEQoUqMJxlZr1X5go8W0VgM/4QqSljonvQru5iRSVk6s8HfDlBeGqLVMy
C4TN9ZpjnsW+0UKrsAyAQU9jddO9wD5Sbk1hxRzwCKFj2k3FtOCJKRzhQ2gRdCqf
QgrI7sAs/71q1Sa5rNos+LI3dOymESrVJnSKcTrrNHEStlzwTLomr0a8uo97KxrB
xQHUgrsn4xlqtX0HsCNLiI8hq0KCMyvSwDUxRrFb4nMmdv9mwNTNJXMl9ud9R0Sk
nOP9L93rwCA8yxEO3wU2FER/1neasEIyA9iGg/CNj/lI+Tc91nzArEf0Xf1GiABE
9bqoSntSsjjMJmyXiIOsprhJEIcaubQyUpQeJpe82EFHD3PRs/KfeqwZfBPS7mSC
+j/QatMA7XzUspDzQGShu8SR1dUzabXVCbKX4r83kjhYOzR0fRl07dUQ0ccSazPB
WoaUUJfoqBUIVlCQAZU53hp2dyWxmVOYo9r6bJeAmd3XfQyzdmNtEjvKgJhn4Kf6
ubtau/cnH6hp+e54eoqJeHYWfmpgm4COh7hzVCZY3jWNaqzplbwOMrwQzQoarwo5
p5enmE64Gg3oIiYkFpzqnrpabJOWFhKaL0legSNz94smWeEaUaUso+PLtOc2+Xuv
JC5dAIvlkTvglV6n5KTrxGZC63llVsN+z/+QT4jc4Wsx1qlXFv7Txhhf/8BP7iV+
k2zix6Ixq6Lnj3v3n1qQfE6J/DHm2ZO/QFjVU4GR8BK0Gp54ITmzwF3lPhnWSyAe
hvxmzm3BlSGpOToas7gekFm+WlSJ/3AVYA46LoLA7MhnBgYvHIxCqc7l+7nBsEzF
8sfLFgO0Q7o2lovkzbuFpdmxvDxyyNPRpZPYeuqJkM2U7JsPybCdilKBC5VkwsrH
Q6N5snWpwHP0WvlTU2H1MC+7XtOq26xtz289EwEudD6MVmhW0ukU95yPIV0yxiep
xjuKMKRkevtyu0WL1UhZHbAmIy/6e00jEPwaRGtauy5gIVciVrfMe2KSPd0CH8h4
Znzk5O8i4lEqgPT/EtgijUZ9FiNLzkyLayD6KrmJLXWdQhILtb13iYs7eniYPnEs
5JHsnVh6aS0v8hjPcGJNIPICLNgenqCl+1ShAPosXVNsKRTe7YOoxyRtrM/fOL6b
bKlACSJ5swSWwnVq2KakYuX8ecS4MVQEaGVeWdBcNO7Id/RGawRsTRdDrlZ5uwjS
eWcheO6VHpZeNiRxBs6MTkbM/GAPLsyPQ3s4/Zi6CFwIVa4XHoOy2HXlUH9SJRrK
OxknyvRnFkLITrgpGkX86+3z+9r4lMkb78twEie6R+BMzWyPA4zG9zqKequm4epX
KM/MR0SzG3BQQ6nX4fNn28cNFbjAcujYOBJqx81wcfePTt6SA3xLi70gVCPrnfpW
LlX0icMp1MMnPeGqluL0CxWvndnHrO7YeEYPSgh0FykaPnfqRO1O8vfGWdqToD7C
p/mDUWNbAyMoUXEL70jcvWyBzANx8enMI8FhjMtzV9Gw9jxN85yqdzo3sGJlrz2h
bQUkOfGLSBvS4gWm87HbIZzcZUqsdUBPAgYOmjlRKnavLPtX2/6+hC6c04zOOxZI
x22wOx/K4pGz5WSjW7+24g9IFHqRNcKNDqlZeUskhSbaojXeelFBBRmUXJsShRav
hmfvvoe72aFlWSRrxZsMNeMjd+NqWjcnm2jKTxG2acwl9E1Z6CDOEhj9ulUMuxie
c/nftIXDF5eeuStmQCpgRl8O3x9NaNX0Z87I8/abctVDNtpd5MaFihcaDyjyRC1M
jJ3ua1dLnko7Lk9gpnpdgZ3Wjk+vwiwz4cnm00IyB3uK+9pNub3WlAQDpPce3vzA
OdW189k1QZ+3L55pwmpyZ0h0fW3vkTdBgV4j/+RHLCqkBSPQNqckkhxr3+oRu6G+
q9Rwswwvv9+Wn+h8aObZ4nNMsfuHU1zByL3A8uVgxwWOYQoX/XffxWcnidqjb5n0
8L+dsoYt41gMZy/+YMlgyc9VoQUyVX9Jbvlm60jdFHQ85qbayzkkCBmd/ZXWneQp
SVryeNXrGapgcU0fph2Et04y42qMcgqXsU4HcBftyjJUSl7ONsYPKz6bpbXz5eRG
arjwRKkw3PnzS8AFNBC6Cjio4VNJbIEGi+bu9HSlZKYkYiUNWqdfFh6JJ/fYSD96
iHBTBQvgEL1VeOJiaq+CUzAQvLWyGvFlQ68jl/s1Nh82mVKZn0khAKBX3bV+h5gU
SKQ2oBUOnweTjTu1B7WeSJitWAQ6xdhICbcnvsDNnIycgZdUrzLUAy7hjzTB2kIr
H9pLB+hnJMGr17b1Fc1d43ZUBCz7O1rhk8k+F6feiljZmlL4deIG3Q4x1Z6iWYTy
beo8nQyn202OJk98ZFF+z1Z4hEQtKCKLS/KOkAayi0xT0gGSs7rdosRAhBtQ3vXQ
Ww5jdJbDZxiEyrHMUnIzriZaDAiENunvqPpra84HXQTG6V40AtQnE/tH/wHI0ESy
x0h//rVeblxwU33Im4ai/U1qm1DBhb2cnOs3biHmyxawJQWjslI+o4wJE6aNfLxE
6UfiU2sxgslYuCuAlxREMgJGQLnusAwONqbGnySMEKBpBsmm+XbjdXTyRuknBZlF
Yy5ymO+Lcw93JIhIWUlgP6FwkU6XzAhWK01SiiTFbSFabELVvOtnDYtACAm0MoUq
oLW3bgYF/8AbAbtls0ZPgeypgTJ10dvFhLV7l1GgmFrqF755NL5p5/vnxn+OA0i0
FX0ibCm2QNXThB+N2H8RtQvHgu91MEPpjcrSTN9JoGLcUOqZxoO+pY4W2ht4pk6/
jEqGcbZS004oW6X5aWW40b5XWE1uQ4Vs54yyloDQvWlKTzxi2LFBGT3S719TDnK+
soaXCQw1FkIWoKCSOLiWIUBTPznEH3JDaDlpJIMdKRkFK7NJtM257nzRIaSip6Ni
m8ezdguxRKxlfBH4FU4lejVOsdjCjVQ9kwSMsQzc16kEWmTLANXacnI+0M0lAn41
EL/yrzfBKOoCmwaDec8avI8yR6OVJRC0Vl383uPwXYxVEqw+wNEEoJ3eqMPJ7eCx
NH7R1ASJOL0tW3jdVUGUDPFTEdtsLvVLvAHsso2aH3XJvneQz2ngarGz01a2Tnhe
aP4Ao3Zo0ih4JN1zNEjCTVwQ0uV/4iQ6L5l02SsBFgbrLdt/eX7FcNNRdojiOw6X
N9sO20XA175Ezl7541gvMoy+dmOsflbJgI4QyGoUNk6H2cd5vvRKWpRkuM/snpWp
mNsKO/9WDnieNQ+FE62u8o2G5BVXwC6rY1VRQi/jOISdxMcmvesHxUYSeiXEOWnh
xukRJePu7ckI611shWaj3UR8AdIilWDge61UOFQ5v57ChaSI+JXaOlAz2AQlsEbx
N7veU0+rXLeEPkBeaASLkFizvFOUqHSTy23fZcIhgYTWCAOP8F2QoGA5G2z+wEx9
Pac33DbV80jdPxfL/z3HEyFJvULHTzohLePv2mo9r9PthQTENRt7cNiXcqYdvZUz
B1sPBJsCwIwf22OyadP3ERU64ej9G0YdV0V0xNtbjnp1F9Bch1K2vp16dHPyeJLj
eCuXPgpJT6fE5DBmrGZmxgaU+t5d68b25FUqMAzzdIDW5hAcRXLiJMhDeBzB2++R
FmIz4D4yxsWUfbhiVkqkqXy370KJYvRqPJvmdPxgR/W0FPwCgaeIVBC3nvVirWFA
yHVFFQBhdj4cH2TTUZi5ymTCHFy/iUMR15qVuLaxyUJJZJM3ID75W2zjKYowuZ3n
CxN5nbHgEKROHXOmxEtHBzKqiIElxIWA1pjK58qTEdV0twSHKbDqKJbXVfA8BPHf
NV2nmKcA0tT/iRDpBlZWOLD8/kNK8RkZY2mNfgKQjYB0C9rH8tVUdckp+qEeVsQe
c0nH8NbHfk7I/bJkMHawgvbOCAVj3QsHu4hbqVflsTsIMTQk9wKB08ZQMb3CLVNN
zYLmUAk5RXo7FjhDfmhmPrib+admbYty3myICDAtGCN/HA0zfQeYyn2YSWI0yxdQ
MgGoNJ92L/F73wSqhg49XlrLJEk4QWOcT1rvBcDNn7Q1TTmRZVFwTUiohK5gKAOG
gDum4XQQDpnBNahNVQrQB8JNpMoyKEHOiwCoMIOhWP485KSKCHZ8zIhY/ypF7T33
gqtk3OI3nZijGs1kK2ZjTmzErv6d8LRGKJHWHZ9MQFJ2FZGlMXrEtf3oiPIqw/ml
MEIAfv0ireDtBhk6LGBq/QVFHHI3FRGM0uPSBGR95SOfcWYm68KK/7NeiwAic+1M
2Q4nMbdWz4DdQV7x8M13hRiY9nP/GC5OpPobf0RMuDRTy4rb8v40lqYJx/lkxs4e
c3a2zMtipbbcSLr7A7SzJi9Yo4YimimzhzXGv5gbyObrkxsMuuHm+arMvyoJcmDy
ANIxRr0oMGpCUUcMgUva+BD/tYyOoUtKJ6iJrDygFeDxjpGe5dnb9NVsp9W/NIPx
1PbH+HapXf4lu63uCC/gADc+3ibO18jt5vSC7ovmD1uwDFPw8bI3fu42kvm9Ybs/
tqiSOi870YUP9EwKmsEAzyGON/rO9scc/f/GrUIw6GG2kRnaU4tRGIaQdrWAQfBd
UAdgl5Eokg4f2Ys2uMzLvaK7enOgeNsHOiRuK+2iRdlNmUZW7T4f/a2SvCTXXj9S
ixVtHIzx0TiQooZfDsNSrV7If1DDAkvoD72nOflj1ZRikga3kp8kZYw8Wv9tcRW+
VB9BSkAuPcKkfMgA++3JWN/jd1RcrFQlrkdtcCJ/efI4oRnavVO+2NlahSIp2IjM
n+MGF0fIQr2xr9w8eMAsT0bM2En4bcUF74BCJMsQSJfYj96tRnuF3d9hdZS9/Jbp
CBuR8gZPbNWjSi5oZw4Hrb+BafTJdWsi3n4+rcOoCpT6GsqBzkpoGjtYoY2i12Z8
yDNdvryM4zeD6F/rdN0J/UptT06Fxy/j/t+IDtBjD66bUq8UQhXC+ezinvVkHFMY
V4paFBWC8YZGWcIv/T88IrhGz1ae7NTvgVjK4MaApCFvBW79t8Gw5Z/vVlpZlVJO
PDE0sP8XpOjUjUtdgIRLbLiKfDkHHfiLRrLW9OMDjrJPvlYE+oh3TumDYNgv+tO0
OmdAXxbgzBcE4pd0yEy+8CnJP3V4bujJh7qpnqzAX/MEcGvg7UG94YacSLGmQ5hJ
HoNpjF3Bb/EomVd7g+RWoYuhk+Y7CiKcgeRBE5JNidk/91NWsg28uCMRYuaFWMt/
Mw10XX4JnX2y+52f7zr16NswU1ij7ZjLFOlTfA4DB+rf1n3Mb/bC3LBO5ix+Ag8v
KyKAf/m7CtSg7zF5ZGIVB58FkSEF9TJ7lhpyOzTaVromCq1RDZziwg4ST8XYRkrD
8+Ebpt9Pat16kaf18droK+cY3kqtUZRYQBy0VtuE+/fBzLG0/hfWlhuTnag9IOFO
Q1+7Byrf1g9t4X6jm7XuDvNs/GELQlEo1yMTP472xgK/5zJ/z2iopWXzWTi12G8x
WRQdgMcxB7Zk4rzeUf9RMG9FsVJMl8HE26NgHVnRqCu00x9C4FyUWNYtcuAa3LuO
ZunK1WWTiIZSveOoT0L5gMFmbPgQ6ZFZYGNs56YLaIjLjou2CbA4/QEP+yPD87SC
yf4f2i9toAbRgtjuvhi5L53yw5+97J/Kd3Syv4Z7d2Qzlfe8sJ63DJnS/Y694b1u
I6gfKJJXCuvEEJSqqROjmLLzuFOFLmUwISPSYELOcecFkrRZlTAI6abh+t7QB8i5
x0vxjxOtOY/+09RXJWdWxSncQ/BvzqerXos5OvrV4YvCoG8odhoYDCBtH+9T678f
eE43SEufKZ1keTp+7TKAcrmi9uU1hlBISaTQUpkpo3wNLityQtIM4NPREK3iTLlR
MAikXJhd4sU5qTui/PutlDYDo050im9ia79oPepsAru8JJe5y6UTXLOjk89zhr1B
qwCxxWx1238BbIokq0cbeIW2kx8uhTk1BhIS3XNXyf9mOiFELl2bY/r82pm1Dukh
RHuQjyLGRLSJ5tO8keJ+/WFreypDe3BUfSBugQs2KknM6YYsWg7x21DtOB5AnMGG
f+n436GiroiLZY36gJAWDrvwXq1YwwCqgEmOOeTVzNNaAidhGZIiruFbxYleIQgv
QDEpOxu92E0V24Qf3gUMDZWT2M3QV/YuQvxPhQiePNUa4n/UuhNKEEVstZmNcErS
R4XP4Mfz4JCuDW8Dc1X3w7wm2B6mwktcMq9vRzJDfURkoeFS0/6XWlk5//Sp8/7r
RLqcbrBU16cbCr1mbD4rXWeXbt91oZEa09ruxs3zcA+IYx64Ws8SVRQB4U38e6HT
XyqlHgQYcm3ktG7lx7Fu8mlBtJLKNKPUwmPELADS12UeBuinI0AOgmTxO79LdjG8
tPo609wuLUrXPB0z9VbJ2tsRp4av4iQkyzkURN90Z9MxUIqtLcbdmlQfRvpq8o3K
Gp99c5a4JrTk3uGI2OYIdN0SQCPInhzACg7HD4rmQgEAqb2zN1tqV9iKCVU+fcBl
skDdWIXmRC3INBKl9/DvYhjpvMNMeHE4cj6ODcJWdllrrwGT3qbyC3aTt3JG7lSy
bFR4fXiIXBSBFDQC6uGHBV+2bJFb7nZgVmh9Kbx+f5yi4WwQ5rpis9ZyHmk4sPuL
voM1UtLh59uy8j3WKuefwAVwIpg/h325dqpxkZtz0xWSmXZg/xkd6YYbcxGKOn10
AENNNazBV0uviDoeULgG/GAGj1mabZRRH5+vxYIBupCcgbiexv+iatc64dOiPPtA
B6uKQPiEEIxIZbYp9ZlboiL/hM1uw3I/CoY316wAgF5Bnukx1HzIRoMj/FgPTUxG
W/75LHlixFOYA6kwRlRWoSmFuaCiFxjBz4gkb/MFQg3ujvPHNxAYMgT1NxmPY7XT
VbtFradlRgBbA0jQEAFEas8c0npyOux88xiQRX1FpzVVPuO03h5WgyGGklijWsal
4AxzrNN4K/qlzPtutnRaxS/iTuz4E99QKK17CnRgDNJjg3j1/wfcnIyg+qF2Sd/2
blXp+rUVCr937z7bMHhB0XrH76yd3XPY3oQBB9bgOinv8yn5As5LE18d6Xp8hTwl
SKcilTRmE0owgkOMRl3CjR27s2nC0rnp73PXI6aHk/3C6lEtKwt+MAI1385RIEZA
Bkt3xtWOyju5nd986uQmevhpyRgKz2a3obHga1Tj8HqO2WiEQnWTy/j5advqnL/4
h1XprelQj+xzPaO0ZoqfQFwXDweXcV9nOlWmS5HNreShq7aVVfu3r+IC4nOtCFJg
pyZ7IQkbs556nwo/AHUB8217BuUelYBfAF+inKsF3dbDP/7TzeZdkrKvai7X2pCL
edJB7DnJ6jHsjj2bj/QsxT6YBkjZhooS7hdXDSHi4u0YL2o54aV4OPG8uBKaExg+
HM10ApS7MwcHWboFzzV6cRJz5xFWAitx3OlTyFR5FRqbgvFjNfm5oKSnubFcZnlx
9nGCINS70HGaVUgglnFQz+hxSygVM2t48e1LMhqDC2NZtDJ4F1NyH8QDCwbVfi7+
7oHTP1gIIQ+4D7eb6F9mRm5GAAYAd/qSn5DsMZB+0YHEaOIyoVS4RGR9+6NwX5t3
XRjy6PRZfjw0XkTY8vmnv3lYgQ6PyBjksiYJo0MlLL8rIgga3OCRMuBuGexeTHiy
2fHd+oOg8B+CqyLAzAUjgJ+Klh/BK38DXTDv/N2ndW7Tn6W7DHQ/3JJT56tUDa2P
LEmNHYP2of9UKzEGlrSPdUTTjYPB/ymGXQHE0CoLkrwh257ML7+ORGdYAO3LM1bn
5CKrW9Oit/H+P7xH0eIL13IsTXRPESM4oe7HnloeQfNCbkSB1i6RmhIqgnTw7O8+
ecxjD5UHnvR0WN32+bQrVYebSNmQY8PTjXSDxJUbOG/Xb9Vp9pPXiYBZTExQdmqd
+0jxTQySnf/BbIRgsFHqzOY+WYzatjdw0hZNe8MrK0a0RedZcBdx4CikD8s0GB9q
xlsUZK8ioPgsaw+9QJbM2AyheRIZ/WS689klR8VYLTo+0G+vB+qOpVUvi2vNks2S
jh1A83nqY/wmhmvJ9lNOjKS6Kn1EYEWoqWYqhXR4bk+fbftDcPvNvdxIXZu1qCV4
+W/zKdqOAwomvYlWM/AmLgIaR69vGs9uM6/wuhyiHBEDvSHRPUNf6KhIdoiE6CAu
CdNWIFcWmR3iuFOZm5A8mSM7MLxtqk9rf1jqsfNf85RIiOH+R8Fb77SJzMLSK2FT
jks6s1+/H+TNSwXNa0aGcSQUdR5QtPONEOzenSO9Bpa2b2JEd8aiDhxSrPBNzyPe
o9tws9YPTu9BYCaFWH82ux55CL3DpSz/oY2OT+CU5Wv4/0Jr0kCrt5gSz445R9KH
x9tog7VtTMG7bpKM4t+gmXfVQp9sRIWrlZmsboQ3fQ5Svqm508M5o+MaQxW0LWAm
MRUyK5FyJNagLDe+L/xMU8kpD5VE0+2+BzhXIUayOdrj0Ngu1UB3Ru8JL0nK9DTE
78PdBSFYievM9H5d5a0YkbNG/yBxGh0GOpO6oqSN0urIxZkfmoHv7+sFFgAMOd6P
rLuT0XPR9peP9DbB/7e69ibKJdPeQKBXyfWpYALQhuUDU5mTjAl6QtONvlLqJ2Q+
08p2j7asMUJlDT7dwlJ+wdnhCkw5P9poKLyqu62Vi/5/fuoOFGEUwKNGmmwBKm4n
xsvQ8j6ZOImqg8F7cQ5NDIXQbKjd78GUX/5zV8NqpkNrxpcJAPNKJSH74MWf+Vy0
g6ibIix1qhyMtUKqDcolUPgjGKI9k8JtdwedKRwIIFEjx7pBfHZVa2t+CbkdzIia
2lpoKSokFROMqpmPv5789D8ZPHCkeVmpCDIulkhy5MdOhslBNkpRyvk2/NZtl+FV
rcPTn2TJHVUqsCrHbO2EI6e1DrQH6RvHVY0gSMLsyWGTS3NgAUmtbgqa6/x2OPDU
17borHh2mBxODanJVwYZfvR67ZdGweYFxLH5DqiBT6zOfx0M0Qo8OiOEtgkHDp4m
gC9UGbhv87WJeTtdWtiSD2boCVAUys5S0onLdzOqolffOlCyG1vEgS36zz1lz9C+
FS1Su0oBSLBbO5ARTondt+PbuXeSCTPCfevD3N6Q4+cfWrEVwK9GleVsh1bl8wZG
S9UpWD8d5eZ/4Zte1J8XkPIwr0TmKYFC173v76OqLeP293al7hxBP/D0tun3xcVc
C64RI1HiWY9NTEDzKa+VN9N60lsDFW6VeApEtrebDv5FbOw9fNXW82d2cd5MD7wX
EI33u8qjTn50O1rHe+0kwADS2QpQ4NTc8xbVCH0rkJc9eOj9dxbBEhzAmUBccbF+
hsblvE/8mysT3QQGZMG6i9g5lmNVJ5SgCI1daITKbJxetsn02PowfIWEf0GxPPY5
HSMk/fuFA98YHp3vqhG82iHS6iQRBquvonHy529cdTMRslr6sJX47eHexnBy3m/D
/zd8QC+Kr/+ccvofDsy17uSRy0ljNJK5ij4eHlQP2Vxa5oTLOF38MZkR+5zSyJHQ
M+rKt8fFxKJiVlyg3PD/V/mGHFbuYzqL95arMilWynR94gpQDfM9behvLnqzA3sl
TmqpUtMhu8puGQ4uS6+8HVPxpRBHn2FdVp7fOHHYExiEoByfDGwYPZFRRIvtQ+ew
rOOGu19XgSOVHqcN9M2kXo2OKjvKpcsxUGpM0FbxntSkfWSGYuAdNEzoY+SuLFZ/
OrI0ZL8TF9ciA1u7zaYtXZH7Os8h2P1g0It1Qdkqm2P+QjsUdt40XUQUMSTe2Iec
Pcmxrcl2XA/tDrsd8dZJ8HtkfG3n0mUT3ikHQUFX0wu7ZTr1iWhn8UbpF4AOttcr
CyKZ0aC3BpVJqj2iRa6fncEz+K6AY1rJ6g+wBkFbzPryFj9CsC8Iu+k5pa0XTocw
E83P4VomNcF4isFjjFkE9CXgbqk/sOMjJlCef99RUUlMXqWOv9WgLdGpDNGtv+tD
3JVaxrFE6dX7f5gSQHyrXRPLUlBsqjPNXkQOXFMf5C8Pb4yzY2inhygjkd7Jitet
PKrrfQBB5BBe095htlR57/623YE8Smb0uZShjGJq3l8cV/yEgHXxcWerkSy2SZg4
o9FEZMAxj0gv+4/dW0VycBjQ6tmPUDhKSaHmDOLmVEvVnMWQLK+Hf6ih3l7AQoLe
B9HLQBdkcjdCbehqwJdyRMZ1le8Y3dly++EnPYL68k9JZ32e2vuQ8ouJRPcsGzPb
XsStJIJCfzodXiNO28xCsey02yruVijWWkaSOepYmSJJG9qi5KTTU+emlM9uMhBn
HmPx19aIb4dde7DJWlu5EWDukcAPGorX0cbTEsC7Wn+psFTwdQR2UoJSq8xDDyU7
euQKTXDSVEuBKvblS4DFhtMewLhAYjz7WR0jeRatqjUR9pwPtiT8cC0KlUijyPOl
5rhSoXoQfhSC8NSnwBmtZmomJFp1pUV8Ih/G3MhNKMqZ3ZJtGZ1Mc7AEa+wSE9yh
nlRPVLdhNJ5++ViNsCrO6sqIONiGPhr6Fqf2ibUVjVOsgIOYLXZ0wepoZe75UR+z
Vu86EhuD64VXWqekPeTSIT1o2eEcMsZTYe0pz31Z/Dx8UHAPu3o3udN7jmWVaRY6
Mlm7nh9mQlHEpUAqoDBGlLGASOaw0rXDco2rNyT9rqMfuEwJAzkaohhN2HLyjKKX
mSeqJibvo1Pu59CY6dkHstk1+vGuOO+ucQ/NukywWtnZ7tQVIuw+c9tO1hajimV6
sBc0QjNc8Hg+NiXtdl5uRTLEHIF4D4Gul1Q/z7bBUU/uigIBZKhlpDvQFE2H3j/D
soG3OZJjQjdCSE7qR/5O15OcJH0ru8gKOd0oJqFmgid6hf3WGvJjiP4ZaBAN5H57
3QsubcoddaNWo/Z8c4TH5YhmQg0O+SbeJz4AuzNpGq4UEjf39ukV2lS2IEXCBKtN
xonwbOCfa5pnBk8R1AK2VKuWHHSWmhFJD4OSJo2yoUvELfVCgLZmNy0LL7lGPG8o
KfNKu7bNXXXe0IEozg+JYgwuaPFbdRiemIFeSwcJyHMmjInHnnw+AHWjoq4TrrVc
ot7YX1AzZJCO0mg5eE8uAtrmi42RErwgVMgbkzhFR7Na4KXgZ1iNB4Pry94l8K1s
4MwpGenPk1hAhPrqWIjja3KwzNP3S0SqZ/McAlj3nRb9NpvPVJLWZStA3EsC7S5u
6Pqq8bOC5LApCArM0Rvj6JVZ407yEXkOEUkMFW5tE7ZDz3CGFdEzmT0fzUTILpnf
LgqdgYkbtY919S1j0D/HPOeuAH4ks1ka5oppz1x20nrqNxgHa3ZsHs+AsRrkZPst
iRWZOMwggvDbBHKKq3/NR4vk9Be4G/qx//RDDcnd9HrGwOXCDnJN2L50BghiZyFa
ilhl3WBNqoRMtKlT+MBwoT7hzGnIq0Epb27TkMSAKWsRfe3G9ZLhqRVmWup2xFGR
XvN245RDqtVwNwSUSOKpmDOlFpbpus9JmERt+vTqIkG4siEsLBxQYRIko9XHumfQ
9lrFhUzSzlhqqeuQ5LdB4W4gP+4yG3Z+vKrdTUR1/KPFQfsxoq9TPFt8PrlvabYK
737n/OFQiek/Q+Qn3ZGYiECTU1+pgIv7H+QK6wJeqQlZPOrmf6E8LAiaJ+JE4i2k
3gA10ZHRltvxW4zLoXtucNOU9kVpTtf69eiYm9b/Q+lHcX5aCreItOss852VkDTk
lNeO/3OMIWZA96Bt9onD89AXNibHL2DrasucXFDWUq3PUSI23XpxpFsWX7zHIsIK
JOK6Fx7A1/9bVdkQ3moE+xDxLdITjcPx+EXvbYxLRDzLWgTnLJM1Gczm1erOvR8+
ABBr9ifwfcXwoi3EFhNnL/NI/wU4w1jInHIcIn4zAQtPIBQpWkAMDNFrLfT/Fpy3
tC0iEiuI1DXs0j/9emXcJO4BPEejG4bvi3ifqhB0m/nzK60m2ax5NiZ+k4fld+Cx
A1XQ0VFVnZzeGFVFna+tiUNeBB3MqWtrVRLVJTbd/TmQwTtQNzwWuX6VUFY9+KjQ
Rtnm39EXfHDyriHz77JdLfixReSymKn/k9Ts4pLxQqbcI/dK/YV5oVOmNokE2b1g
eJ9TnYoZwiZd0gj/FCLAQXOA5J62fGLjSon4Lxi6FYG0pKiykFU2SSzjuGcDzXmn
L1LgWUOjDHjGXZRfU2/AzvHUOtwz+R09Xuze/3L7LpqdsuC+r07kdL1/y3zY49eJ
9ugMCU8+iLAnKUqpIVoJQnRABYnhrKZq9CvSvtjfvGrwQ0IpQRF0DyMzpECRSIzE
ngQ9b3cvzce6qKgUbiMa5DN73fLfeuAQEJnaDZbKU/kw1vkkAWp0N7j5RbSLr7GY
KGmuTvH2RMJLajEPuHMJq911XNNytCcCj5dA1ldcRccAUjHsAf5hGD4XTuJPtima
gYgZaLUkUxNFv2rC8Th7wTspGB9gLBpj8pLXsgL3cbCQspmCnC+hd/gKcCLsNEyo
W/7sNNVqelIhErM7GR6JkGnV0FOWrUerA/kyZvi97dljAp5bR0nGO80dLMHztf2R
/4Fny83yrmncqQ6sJpgCybmj90QotmQyJB8XCoJ8b0O2r3SBLcW28qiUUBASi+IU
s/3s+Ecc9uUE6rYP3Op8ZehPPQsrXTqdcNXZVYtHR++ZBBvANot6clBTYPweKpjd
7Ew3Du39jA6kX+QoXI3A2mBu9T8CpSb6Db/SSWD5yG8xC7vlqy4FrrKXhL1oa4OJ
psWt0BUsTz3m3WkMuSsB72zdBOLFDg7kKdTonVBKgOv87X8wgm+2CooN77+f1LdA
69J1FLonBuUahCExndji+n4wooa1IfSJT1jmbO9vi+DXdY/MhWzpqd/uv/RifhF3
cmof3uVP2bg04QL4vQZaUDGeS7OpE869t8lz6ZpOhua2w7HHwF9DYrqSLW15Mnpc
2LZU98b8a44xeIXuLzdttoJapeAnT7ahjK2igoLLKg6Q4IF5JLIePrpq2Qonp9lA
pBIDoSRRrwLgD19lOU0QnUKolY7tmIdhK5efG9snTe/vZzxQ14IXozq0CbmckqWu
ZUof/KsQVQ/X+S2xfKXM9Fhvo2nuUNsYaownEabO3lizT5B+ZpGfYMdhKMfpo90L
9mapCanlooXsEW12pzyc7ssMr8jfjweveEV4mtdIB/iLz/WkIrLMKrWgs+FTsJIY
BYUk3wdYKgarIKNMdMYyfZWWte/RoLoTlc0VS9KrnVM44znlea34K7pYI+WsC3Pz
277ugcasb8AHzUVr+JzpM6Wd+eZu5PzUjMfuFmgSJBb5W/4NKhM0zT9GRL8ry7UL
syfw5ZjUYlbz4+U1hFbEF+B9iw2Ex/GyoOzhHTaWScqH5Q5SMCCyfrAnNTj2UA69
hDqfHTuMDhleeVNZRJi7ZgM9IWiVGmAeJ4X64yXD9g6H14C+sI6PZRfjLZkrOpCg
zBvYyDgeWrN13GrtM9dKUWfAJI420Sn/NoieAW/EPVPPnfo35sSGiZg5d65Toqmn
20FIIHoYSLDyP2GPS5G/+iGSjNAVq2RuuMyRR66NHJC/iKE4+QfPxJZg7LSB0Ovl
tYeg7pARbOgS2i+1lpDJa94R6K5SnY9MCfREalDE/XjRtWWY5uwZbZR96AA6jsaZ
fvCn5vBen91JQQFYMBSTYTD0ZkNj49cwcaoUwXSAzgiCqVzqJV8CgiF6b6EXPisp
jb1f7q2mA7xDzC5oUJn0yEGFAnbOWhYL4qH4dbx+0vcwOpwZRtTIA9pf18wBp2Gw
z1FIzHf+mNDZrmBxIj0DSRn/MPiaTb4bgufriC23ibv8Q41E3/P/NTNFUjLZ1g0r
Ho6Fas8yEr6CU4JJEGVEd9sYHD2CVkRHC3hi8S8cfZ9AVtNE8XW28EUBZBkk5l01
auNkdwFHaJMYflQx63yrzowzB4bi1cVbFvdoQmHNxQauGExl4X7LfOTqBiRd6UNV
Y8aD6121TCSyEVnGAdIX9UPrh+EcBDNUznPlclZ5HZa7IYgLIkqDvMpPXhhqiJv/
vA+kA7UB+GihFZdJwvk2mf9krjUWOSXocuNJ26W7R+bPZba4wKDXhHWSVe5S9Xbx
qgranC2ebxXOFDFZVNyFhZwRgjKbsK3M9ByeFjFfqWp/xTnkIGaUF0zj6TCXs8vI
EOdlqZftYH2i7bMuEnvUhZqYB7gTCnEnudBGqswiGZ5CgGzjhsGKdtpQ/AS7evtQ
MagSuNOg/SHKtt/almJw9aPhWAAlcLPDDjhwwMKRp14Tzgc981lYIKJm+rq1tOZo
mgr/L4TUNYeHBvkS4dNV/iQYWt1hS2wwTwD0G0fxgyB/vp9d1ehpF7gMY1WN5re3
uVMl6oJAyj0+WfENzXEe73gMGrkje1iJWzraEBmItVGd9xeDg0ofgAQWq9RCMr9X
Uq2vbZF1PhOH8VqiQwF/Ciyp+hLCMksGKC9FCBWWnpBwIRsYu9Idxtqen/3zzdwb
ofwuYMfAsvtOrgpMukfJpzJHuDCuGFEmbZS21yKhZsyizJ+LeeIafuI167ZRaYHA
fFCuAhjiB8sa2PlcqTgP4BwK1yIWmlWpPzGFlwd68zbQzR3BAioxDCC4J9CeV5yd
iSkXIYcLpcT/4NEsshSc64TjY1g3vRMi/+pPyKizlaRm1N6KYb69vbvwNILWMuvZ
xT84Sa8WV95SAx016FVXnZoYdZYl/rM2lx7BeUd25UKgAcVgvBR5C9F7vZOZphHn
8dHlX88lE/PGasPgPn8xCv5VirVyfeH0HODCQe1poveEJIOKNX4nW4Z39/ljdqi5
OTu1kwT1+i/mxw3ZKe60OLnPoZ0XvJRCMcQkR2gNPyE8IfVYQINwe7eT8TK+Xkc8
aLhYmERdDoWMrAGKpNmy3h6Ud7cDxMcP5j3mMMR8O27+dGT42eQD63hUqnyoEX0H
PmIVFNZywyfw/rnEq6QEPTRf+YrafYiq0gfEIy70gFT80EXtQSemNaOTyRWRpRYg
E94SPWgqQCcpnVlUNoq92RaGbdPkn0OlMWoctsjHmp0twDSeX/dC2Pr5w03Xur1R
ibJoY5OqZUZwgsYu5SbReqn/alF875irCD63KU3ErXu5r01KGy33o4Arv4JU93St
93dtEGxFOXw0YEgvjtFwAsu9zmOhClBIarWxnDULBNhXWiN3S7GntAZ+VWhtPnNo
IAQC+PyGfHRtYaTh17UCPPP9nqmSM2I2n7k6pzr9euO2JwqbnhcFhOF+tQUVxxkX
PSIKrW4m3QmqG5hrddziRWp4Jrh3fzCT5Kbfr4lrsXNlGK9GYBYcsED/BrtZPxlu
6QvdtIXc7TOmUVNTd36b9oPgvhaKB179Gp2XiyEaSX7WAIB/XWYXkMV+Y4zcQcVp
ptnxEKOidi4tal+lGwS87TXjongokted8cuxXl8oXCv/mj/SoeXSTvS1yl5f4TFB
QVkDveCyJr9QmwVnKlotOe6Cb8vvlI99ak+mRtVmQrtDdsvGkSvN2XV4X00qljb/
u4Di8fsqv2jw9ZAdV9es44j5edFmb0iR+TcvS1buzLBWYUthXGJvxsRwK3QM/2Ih
3B695A+t8St+8FPktV32mrB7CvNXLLntLgE2Lhp2UAdPuZawAgxuV1B/xpSudTUG
rpqd7pOvppYFNdrBj1C/d5J1UL/RPNKmurtnxAmq8fGA3nxQc3wVgu3Hq9LniSm4
ZRKCAln1kdINClceFEYKxNzQ35Vta0x2tUniTO54GBJCqFnF/YLVKwm9SGY7G6Mh
M1px5ZNrYu8Q5uyvlqMSOR4g+1iiOsuXBmoStRVavfbBckKB/C4snYNo3uYXj4zR
CoJXBYukwblp713qaJvoQc8SBEsD9k1bm35rTD3uk2t7eflnR3neRuLxfHmf0qWr
caBJk/SmFTtnTU+gfti9JnmhD+UR6+aLEZHtgGSZp4Tfx/JqRlcEVR1H9aG0HK8L
3f8mVrH/HwT/yA7eQ6OMOBygxbKLtD+mh7leRizjmDTgmG0pFrTexyRzjNBrZfD9
SamV8cx0qj0buhBSZ20tgSMpazF2Vtz1lsUgzuNk5AEWEuuxsAY9zGX4r5EFI4pf
25yhaNk6a0/RAAh+L7dOd2PBcWZZn5kKHn/evcKO0O4QozwG66yqsFfJZqWtS8jN
icLF/O29QgSg0UgGzWNfzvUN51lmelz3ZY5yTJGeLkQ/c4zvue6lsTjjSu1nTLMv
UP9vgS5kYIHBzFjzdeGkb/oNmc3wqaLJRNef7W4xVuo54sj3JtP3giSPxU3Fggqw
SGcFNVfoOnPO3CgeqG6Ij92Qs4S9S6ImMQsjd+1knnGLAtN1watVSWt5Jee8vdr2
l38QvLrDBd6zuIimY0N0fwS4mvoGqWOJ2mzYokFSpYnJWD41fXn2IZRqN/j6rkG1
s3any0uN0PsblNFdkdjTsQ/fY38GaTANmULvOazKPmiin4PVb4bxc5bJjIW4inTs
BQgFAxxID2X5j1TP15vbEIyCnc4al9Iam5mj7LKVjlu1k6vCBjopFrrFUiasKjQf
xSwKbSAWBcjpYqGsUEC9l5ry4s1qdrbWPLazDZFAkbqcsqTaMF8OlpqnNUo+hgAT
+EVzxyIgO84/615i0inp4RiKkFTN/6SrVBXBgrYDjXYxH/JixtGKBNuGbwdpBDPs
cFJ/oIdZMMTKt6MHiO5d75omMpfou9DCrQYcJTVAGhaNi1F/BONDkZeknoZbjHhk
yLs7ziPzpg0y0aZyLviJWPWodS3o1jyxonSRVl6Qm4dLWGBbIyBkEPvFTThZuJME
64QXO56cTDO+ddDBRMMNmeQEJN7f/ZOqJinvXF5fYWscnCDrlDuUedlAxBdjrgOz
NjWxdpEoT/+ERcBxymxXc0N9XD53gBQpHy/2tRzqYLdUl0wcQqjWRKPdhrkU5TE4
gWx3XD7c0qszNgMg5NiNOIQXmw03W5Lw/z0ASuYNrUWAJgyhSK1PKkj7Wp657SDo
8wSeenD3ZUyGv2qdT4wHoj0p4uFcletR0vvnSbjidbT6AgRb74y5qBI4IjKXUDVn
Y8qCNr9oaXqi9FAJ0bQuDHT9vNxQ/81BcdTlWFUQxHkmrBgncZ1jUnr5mvFIKOuO
Z1GGdICPO5JbCwpxsJju8HTbsbL3haTppzMowTnoVvsAOI6w0tR79Gc3tX+KIMN/
EtK1pHlO/lKGRzarlnNbaNyNepEnSw+F7Ysa591aOlobWFu0ZdbCO2FKRhBc3p2S
nDDAxRr+F1LCl8Z7rbvlkNVPZXvO47ErJeuB0iw1gbeuE7OxA+T2WGIR1UN3oYgI
zG1eEcIllEvi7kcZXMBS6qcvOmT4FXWBR+Zpl3LlLMerssbSKGE6UgbucfPIGF22
6EYWhR83zahZg8VXIW9KcX2chsEGhQELuxNqPhbIvo0+Szrkz3dS83I0/jpAsdL6
8FtA0HnCIwJCCfMDjgqnOvdeQOCi9HyuEoSH5c7PCbSejMdO+uQp9MQ0EidmG4r1
nAK6W8KIX7tAYcyBaqMAPqxabiSYh4/FR0w4lglDfOR1N/wMUAjzaZ0o//qJjHQJ
67WdAgdyMGwHtD69QGhMwASODVcuZtYNzT2ikihDxSxrU8igdKonfpTKb/p08kJV
r6zvd0f86Z0py82FkuDxbmJBjA/SeGLoR4llwK7vr48pjQczjQa/J1NYkvZXzDHp
bKi5vJjrZ9T/ecSIGi7F0kzjNLu8afHRDZIuo8tiIdNGawG3mfdSRdin1ffP3H9I
undCY7KSF1vHofbdTtj/BfaxSLnKDjultJ8V9W14SKgv3Ra7PAhIQQuaRz8HxWx6
ZP9P716WDMAhFr6SOMR3yP/8CbD4UTiExCcPZFgg4UdahX9fQe8xKsi0vCpYuV3O
kNPXcrcOIGHqzqolpG0rySPdl9LoIvGdM2WgROYpkXDvQDHvGE/f9IbwyHzZ0dfV
VgVsVC8NGU0mPWY85hXOesXNAA7RglH0g/AOU4QQINiG6TAy2lWo33D3oN6JHMC/
QDopMAsF2/G2vMvtnN6Pp5JEpKags4TuURPnDZGEE28mLiDfKH5L/7iq55AAwG0Z
kA6Wd0vby9Tl4i1Z5wZb6HrOgGSi8uGGZXSOcxZzd3laWx5zwwLfLECqvs1GETIx
wBiPVXLU6U7Zx1oymAfFhUdAaooQ+2u312fphZPlQmhruMvNhUdOiuqX25tDN+nb
kjiv8BZgqHC3YenFzaJLsQb9T2qk29RE0FFH2PBc+OWKMk6z9E4zsSSQXC2RypR5
Q88wA9TumYWl12FyjgZILZp0AukkdpXYVKruQGYbj3PleGWzsVxB8SH90pOlM9zE
iXFA33POYSR1+CVpKiQPIHTKBROE8AUzBCqsnEB4bOWkxAW4YK0MJoyr4yvj/8gq
sDp4BVOJKNyisc3JMAG3PnLZQXXYzZUnJXQt94VlB9S/q4fzn1otA65pLvbsbeWh
PeGnhiEGb1PZUiC0CZ+VACcTFNYFbjw6JJ/xwONylM9qQIoZHYLNtOpZt4ZDtHNg
fl2NCHwJ5aWRWyfG+EQBWVw6hu4oOrfCH/c4iPXwzJPyGAICIahqCzDOhBbrutMf
kxMQtdDW3FcGzLH/piL4sCjjZrrSzf1KrSLFb2mOtUx88pIu9HbraXGRmcTWk9xt
KUj3pmk6P+IWYXpZGkrAgtNi8xVQGPmdWdsm/zbQ4Uv8MunIUiOQPTcENXJ8MSvC
kDPKDlJwCgGJdHExQcQZt+sN2oHoHlhG4t0mKiVGkoEg/8xJiwQXb3vaJQNTitkh
oHQ9xIaYGvGIUXpqAizK6oCmX6y0KY0Blp5T5YdbQyrEqXtY2iuZHNZnBEMuEkxu
ial4603GQ6VQ4hdsmlhYCccYRtRQoqj+Z06sbx/qu9eITy0ruIleg8wdeLMK86gi
7+ejjm2LAGhgPrwObXB4ZalW1WRsnOPYvewkTJ8aPgmTapEVCFAZ4m6cxVg32ifw
Na7yU31xvjsXzSTnemAkQLQjqvTVz1JvVycZRH7J0si0Z61EsQf2hbEA63FmVFoZ
PJJA6mF07IEv38Oj9RZQVgHwQJlCRubdKtRGnMLa6UoQo/50fmkyCKvw6lt/cLbd
AgB/sacKppDIU32j4U6v36ouozezxUVdh5wDvWXrj3ZmwjMBh4BbW5W3MvjHyUK2
QP5S19oWPi2i41JxqC7RwTIWA3fLsbulq8arDgsohDUKqX8qDGikkY+kReH980SC
9S9jcR/Ea8Xu7FdqWa/er7kM3ZEizL8D0VEAYa6bfp219VFj/lsx13MQYKivj2xw
brYAG2z65IXR2HTpRhOAwGhCit4cB4J3bPZjSZzJiqJG+B/TWiln/LaPhpcftXGx
MAn8etoN0bPWZhlTjpi8yDm13jrRXskDQNLjTPn7pir0FwH9rjTJ0y1YHU/CTT/j
EAhySP/U37SJ401WpjwDPdKEc3dbAWKoJHab1zlj6sbqKdArof+8ACBOWs1/MWrZ
KP49RxG+USL3n+ypm4vbbNsFQLseHYhUkcAmL25TUHQ3N06J8me/rMP0s2Moy2U5
PRfPzhS7QKJ4rVJI4pIFOlkJta6fxrjkrosuC/8HVfRDDg8HeTrXkHECK4NQ+eUR
bQdyP61h8AxHddSmunZl4160OakVkWQI9ZwLJ8pwYXB3b9omkWC5Br/JXD6VaNVk
JeiI/S9+PMW1q21qxm5P8vyfhZcO8Nh/3rkuKjuc1203KuaNOxzflmaiwAjD6Yix
3OkhZ14LBT2jE3owadNwXvrOtjIiYmmtYQiroLGIGtaaJDVXQ/pg8l72lSuRt/I5
xV1LnX0/Rtl7ybZTfpdet6ZsLccLzy28LyWz1viRuXQBIj6x/PFUA9bJJCGAV1bR
aSs1d3yqKaAujRol8h+Rs4nUGkR9FfE3dmk84E0g3RiBUCABCehpVXJyH+GYDGm1
/U+xgxePB7ST9Scs83nKOgKJ/n7DHriG3AG0r7UmH0WuA82T1kkA8tYyRaaP9W64
cup826gCl5F/HhSgr73d61ptcElvw7P2rhKZ5TnY/JiucNB5V/eV04qHLA2bVLC4
kuszgYVS0Pmtdm45P3aWmiGoJdKf2R0nBgpo/OeBB1kNyWuDWb2bR4UGKEMVBrq8
7ulaeAHH8LBjFIVy2FonKtq/s5upyM6MRgXaXQG3VRSyL/XoNeLO4Z09ZpBCcxAH
c4VECArWW1sG2e7P7TW6U2Xxlb11Zg2NozytXMQ3kaZ1yBunSI8In6A80dJCJJm4
SWUaj4cPRxYLICbjj0LovqatVur9tm3SP+1xg71DI75TKio16iDCxxKqIoKLyema
hK5HRCJ2frBvkNda2oRfMQeI8X6EUy5N+/4rf1pRVPuajyr6KTLKU/g5XtcSMLBM
HSFIaF1W7bSuR0D9HEFJdtTq5HUza7OwXeSJMjVYIBIMYF4Q/W3kNZ1eMaUIWzFp
FftNQmEqDSjsMTVomWwCbh6XRaoW2KP5Ee4BX2jwsyjzDk7J2Yyj6CkcRdWfpeDu
Xm1cxvAYLrIk6UTg6VRZiY42P6mRg+x/j7UvEqPX/xhkmuwjNyCvS/+R5cUp7tx9
dSFNI+hb0flEhzYal5/keaymAWC1xxVjntCZPsnryCRb7FaVFr3dGLswecY260BD
VxyX36bpAgFUxn7IgJ/PY/8fXRIMDWBt37a8rXxXPj53FnsWPvHvIHmmRPO0m6ek
c3bCtqSerfzt5ur+rc4CatJ2Eu7CSjrFOaukWaUbIvS4nUlS7yIpw3BSMMoCmgU1
EvRqFNvuUXr20WsYbAoBmdCuNLpTZAS0CsWiPtdB3z7stxddx8gnAHSb9ceK1xm2
N4O0zC3Soku0hJeUo5FNHe6nfDKD0VoDtequo3b9AP4U1hfqcVBf3Qjr5Bx/NZ8H
1MelsiNH1udfVl4PD0Q0rvPSxFfhTyYMxWG+30VMW3e441lboCNK5HJbOLM9rD+2
6Jx8FVsl7KKicybB+f0Y8n9cVi8TBzuhtx5CrNllSLvZzqXzHqnI8i4+35Tzex9p
0wxCiXv5E0yLuymfYwu5hkFl95FyKEySKqtVQwFgkzXdVHGoOsMo+SjuMAdPMLb9
+dPfIKgEdGHTBklzxYBcYXZr76W4PR24p/c+czyj+bFen8NsXUCk+estBVKh/kRS
q9CED423hE6zcqXtxlaVolQ3XVxXCu8dOlfb7NE6slai320Zt/FZfb4Ar/yc2xL1
zAzqe2m7jMjwGnhNEqx+S2nR8ITyYmxtqX3PR2wMQK370zjU1owvwJOUHBPQAVfG
LNCflZSC10XZ5Vxq8pRVcFv1dTUEkUYrWsqzX55gvuTtOi/MDZb18X4+hLm37fF2
sMDvExpzd7LirGRQi78VTT4fhxNFfxRq1wUhIbG7rKR8XOJZ5J1RMscEXor04XK1
HwHhsIwNnVMvYeAVPyq7T+wutbUetNVvoXME2MZZnpM1vGczRh4bff2o6/lK8987
ozYlnM0hj6LpSL9dwSfF+Rd1jnxJSFqXa6pBKHb++VuAK99g9GjIVkKdxbN6ptFK
f6gGvkprHa7JVOxvu221gJAfTgtX9MZ21bG4pefR6F9BGoQ5gz6G53DdSfj5aru4
28YRFgumF21k7q0f1lx1Xm7F739FWLPPpRiOpbm/dJzi7bMM77jPTmrwQG2Jsfps
jv/3ToPmWzOVBUGYFHW7EierVQijCxglUeaDDRhGVA0V3m7nCYwFyZqgfRlvmbpX
JIlVpIrdx013C9bWV6M+7Dqw+sdi4tAAASpSph0vKlTkwzqZ18ZHYLc0svtFjEUI
Sad1yI/0HbdYmNyljH7pgRLkIJr6DkgX38PBFkEcUE0+I7YZvVXGs8gOF2MuQQjH
lZOfOcKMAw5dOXii/lhBBAVuxPtbhZv/r40TjDbFm4ukXnfCQaP1jYLSwfT8TOxV
Efhju4JwexzDzlYR61E70zrUA2S1d/ghVw7v8egPVU4xww0QElp6OGf1/Yl+guzO
/mKVs3m62bKqkoQ/543DixSjYD2B2brnL/PL4iiUeC17HIFHL3Is71j4CnM+2JQg
iLnkqjtFOPTTWddQQzLWI5iYqw6Af8vvO8BED8V7wGsxQnRx9mJawD+pSne6sCze
X6NNKO52iELx3VxXJIPjarFRDhjZvboQnQF7Xj/j7BIGpQOgWNoGQrPiYTqM4hOj
PnxMZAPR6wDrzQvLXMaudVLpoM58kMPtcfuT9+0tc42DnAj0GIPDCmcDKq/FEUFQ
01/EInL+uW6zSKzl0uTWQlUT5Y0/lBOwW5h5HCCAdd9rV84eZL+BU2B9NtFzAJGj
tucOd4OyGv8Bg8xm49U6r7SHeFA/WJ4GxidEm19JLOTk7ZlYPZAuTtJhYqWnqHdB
wWPCh1y2TqFYcnyQBGVUvYotERcPEbO5DY4CyVbzhTT6Ti0fYwpuiGlYHbVVG2WK
KmyFxS/Y6uve7y3QjY6seI/h4wJg7Odad3JTiAYVJxM/P2dhLNz2HoW+gd5ZOerV
DmEDYFg+7smktwG7/LQxM0UuhuB/bvh9SZTBu0GtGWADnU6/zXn1Y2vKnrFA2YaN
Xqk3JJcyn1a0IgPMY4mSU/nOuQB+U8fD61YkMHdcyZjTWAzoYyeXPhyTaT05+K0N
IE1Sy45T16SLSNybdzJZr91kpRFAolWHdym+jIHZYpucoYkrp6u67cThTxZYpHtt
IRHCsJo4BmA+DwxmrpuLwwaWh/VqAkcG75aDX7S9ifPUFrGdQWejEFoBMWskGzVd
g/SePJYYt7Nv3AfbloD1X++pi0/txRtpWxeJuiyLzPtuaTCN8CQBc8K5zK1pd4BG
Sg04o/11GBxdB7N6wNxeCjj1Dn6eZgg03kS6IffNFivRA8pB2si3/Q66B8yjbRvX
HP4PtJUtFZ5oSXsh+cCoMPTOUWI82fuy+O72AVJg2rh9fkFnwCTMSfJ+tIzwXZDx
Ts8rxbosMMt3CfR9onG8n6TBSLRJWaSlPZwpWrYQ9Y/SQpM8WZhNObcqpCMzrbtQ
1LcwKv7x8n0I3fTs743pZubwYuXmBjPaeQm/maMZvzYvqR5s8xaaJrfnoPRVi7tt
LFTq/abSX8lxP6j/UlzwHxraWd0Rqz2Ep2sDOVN7xRecda51YxLglYvzQptGXjYb
75z3tN4pFLjMUDJ1mPduZ9qYZA1lPAleH57MUGOLGLaH7OHUOvRXKVoOlSMA5gzt
GrqmWdydI8ZUmG0/mxMCb3GTkxDgL/zkSkPeevnrx+4/jtjgmffetafvJrcz6pEh
eHDmHRtYZhsNfoB5ELKOD9o0KCLkjuN3JGutTTF3ytYUtsLGMXOaKnvr2OF5myh4
Gro97vDqJoVThEgU2UMhHck47A8hcU7zxPcHHwkaaTPjcqUOrE3FAD912AdJGmvc
AWcZSQyOmqGstE2VUJgfxRNcK5t2njTZanBVPLOjNEwe6iGSKX0Trnmhk7H1XJkW
XK/laIufTi5FLM2cOke2AjiBHQCJNM0viPNTAvpknMv4BaQyBMJ8er7+jLNRxe6A
HkeJFOEh73sH7lgJMG1csCmDAdht8Dtu3WUD3Omn0ec4GTibFsosyTWqb9ah6qKp
vSu3N1HSwwajrlySP5vzV8wDKnM52J/nLLI/hUEIoyNrotDsTh4An+LhfbDPcjk7
2iIaDRcFqCCxFmL7VWjD/wEIkrLzu5UHoLVMMvhs5VTRBktcwOkJNnGhitkFzILf
udrLQfF5XNM+EipoG7T3yJeP3Estd4o6D7SwIMFhJ5MzEa5rMxh39gv9fhyq3T+Y
8XmwASHpZxiMudpSfN2BT2gheR37QGzX+t++Tfdf1IN4NLO+CqAOtPHDzI8TH7GQ
yUy9djAf34X9mkYj3xReb91QD6F7/Fp6JEKyJdujprU3uymsyYl2uJXrI0n+kicF
XgNpUPnUgzBpym8mkRaWQLUnntBh8zbGUm/Nr5Ov1PSGuOVlWZuh9TqeO8p6Ewky
XwDjUva1QP8crIv8H9SWyDQFYkI+aG1U2ZVu5f0AXdrAZu/tqNXoeTwRwhrBYqYd
0jOjJWRv5MGczSTaqR+D1NPOir/huRd+kiztgWqEw3qgnAereouAoxmrP3ZSEs/c
THawQs5nFlBJiga3CNn3UGRxcxrRa8dtwjmYFH+YDIVLQ1PaXxj+9+sMB8V3E16G
FLWt+ht0d+k6WokwZz2BX4L06rRhbtpsrMFdhskbulJaViKyq7RQZZ3yM2SWlLZD
lpxzzK0djaK7JpfeOlXah184ERLh3c0/qtcd/V5cIibT6FmIClmephsaW9lQeKQI
yKokH85rLoNQBF72z23d5IZTMWJNatMck4Q2BxcCQDeQ0Wcjnv8ZCK76Z+d/D6zq
3Cq0IVM7oAAYyoHw/GR/b4sfOzR1ktAnTFlMnaIHIv5rwZWqLCnpKvGu4BfDFvp0
g8qLf9OjgIWN+aCToI6RRsqcKoFVKTHsiGl/p67mcQW//HNqoLgzY5TilPT1ySE4
9Ol0WC009hbt0t1e40WOweZlGNd4SMPSkDa+wTXqBMdtsg8sjvFX4vur3rklu0Bx
FKALFWqFQcMbVtJsAKZfSEowS4oYrJZT5nG/0Jw+VLuBjYXYjq0qEBtzWURoVVJp
FAc4LSOyoSj6Qd1GFiO2s/kzci0C2lbkNeljpPAUNFgkhpt58XAQ7U2EtOTfbu2b
0mz6uYXia7Vx1FJz4VOblt0tOxM2VdJWys/yYmdX0IxL/UZN5uBCxYz/I1v7+G/m
YPsHLz3XhbFSDQ1HAhtTnq2pnl7hinaZi1UAtt+YLWF5ff96nz7VjYhX1ovPYAz+
RULhP+5c4+h9InESMfg7GILBV4oSj1HCJwK1xYfJMPtmDpsRhleYxRSmSJBW/zKl
ex3UHp/GjSDgzmJSptu2u59YgS59tfLPcefqg4ESqjUWjDff/8ga7YjcqrYsDjuF
3PcOmC0y9XzIM2+639Qy2bIGiDX9LcDjSqO6fxWwzDSCZ4jxtg5Gu0rY6zjepnro
+i82gq3vJzpZWKGX8f9hOP/Zfx/aLBRn1VUiv6VBooFLtL4mM5z/jsayjNY/523e
Obxo9mOi2VJ1SqV1KHTLdGRfRsasnwUkl/YlR1ATxvmzOZNr5LoXOpcCory4hIS0
8urkJcwWuqxfXhXR23ogcZ33T+ZYqaK8ltd4nMJs/NDMc5AENdiwXx0f5uG/9FGf
qDGztGBmY7I57aR6UOzNw4qp7i4w6FI8IfzsDgkUXyQjwBCCgxMLWesBhdtyVZ0J
IDBd9QTktxvewb7cNN0htfR4q4ZJBVIzVYa9FhUdEW0WzCMsG6RsrFTV2nTMx0NR
xX4BP7nhTQS9fsuCxaJOXI+Js5Az3jy5iYtsx+mRpf1qhSD7KFBDbxjbBqIpsJoa
N0NVx7zQoN1WyxC8Y3UQ1p3WKmf9diB9YQrnNM1E7Pd2PLHNwiUVvRTtAvTjx8H3
Y0IR6W5Jej9ilixxRVYNKTe8rX7ktFUX3WC1JeMpzir4Q/dso4ZUEpCXbynwFAEV
yukFgBzTngi8BiOg+oO0c1aelYwoRzU/nPjWMWTM4Vls6esVGIyKvt/EcrROrABH
8ceMx4DjKn8r4L9B1KK/Js614+zF3SLpFNrX+CEAiTW5BtcDoow2QeN2RpnjVfCX
awzl4Q9RcMfsAuNnvbMnBs8ZqfdFTgVrfPkW8RR70HVsYtJmm234Bv7iAPjlEGhx
+GRqTp6U3m9TnHwGh5beg2+pNjHEz7QjRDxFjRmt0VRkroKZQ9jppBSx2aNpzbu2
X2W6eE5+a1XbddqSEW7hZw7vArfvFTr1Jb4QVEejre6ycRJCP09uMBiolXF982yz
409kfgjfFPSow/D1VQE3oFWcs060qak+Rz8j/QV5nG8SAuLvaGPP9gpG1EMrqHVR
qEZ5EkkVZWY+yltx/RXeIvRH+SP/89CAiJCVlIlpcpS7gmMbhCyIadUVINgmH9b6
ujRKeVijHCwba0w5bMLRzwJAm0zznomuCMeS0pPOwmAK4J6XwtTUG+v89BJcuQCc
fAFH28Wqz4R/U770e1PzAt5zNANgAzV6xbB6Na91nJbuTZ89KXwgw+xv99rDjkTv
QEoisSzNvG0e5INUZ2XyGUTyQfBR0/9SSHSHkPpIXGX9FadiEyy9iLNRif0tjQW7
w2di91Q+pwc2126HNUzB9y+GXEIpUCF+7oDmRLTwRim3dPkHXY9BylERsr2FRfEC
Kxm/5s06OEuojuaGFAzSLqH4wwBGRVo7WKpPwzZ117P1GBZ7RhYi4ImPKkaR4kLf
JjFgX31KBBkZP20YPQ3sVGTg9PndSyAeB/Cd/lQaNe4reC2DVNLX3+iT5pdN0RdV
cyECkQzQHO/nos621cCnEMQ0D9dD3NZ6xxmfZif/EJw2u7sNxBBs4jj9UZeG2jCz
XES1J5dEViBrz5b1Da7Rc6PQ1pqaWVZ9VrBNrRPpTpU7YaLx9riZWWAAONRxy0AS
sMPGtrHuUE392st26ovJ4gJYC9Tlj6k20dPrtIGcPx8WnGMzg0IUhpahITCUn46/
RO+vXGfkAw+SNzzLb1BWFvw8BH7VdF24xR3IN2vAZ+WmZ280FeQS6RczcPkUvvlL
WWFlXhAOKZOcolXoftSWYfwXhl+JxJoITRM7PysRdKQYJ79Mw1GyM9kdk2zmq5hw
exua/DcnwFx9Z8Isyotvic+RJYNkjLikkI4T2LS6Qvikjp5WOQusR3qElckvb/5s
ligQQafM4RrVQx85eHk6t4zbAUpHk0rOPv1FK/qmsve9CoL/Cy59kTf4t/71gbUG
iUlikh/c3GhUkOI7nKxyVrx1yumYyXo1YvRQaIeG5wAbv45VTUxmIqlCcCDRTEmj
UT0M2MkBVIYsMJOEhwECQy1K1ZSIikhrgdJKMefXqN1+c2qoOUFfl9bnpe9tNrD5
zY9nKd8wV1IWVIbUrM/hQr3q+HCRm8owbGvvpQJwi1Xpuu1D0n5TKUqih+yaK48y
QrUBP7asfZHiGC/cbnJWOwJXy5fOS2LFUg5U6K2B1fKJVjn7x7V05GzLtxj5uJVG
7L4Ahyb//C41VID3E8RmHyd/F+nWhfw096fguuqvVF/RJAMmnCfwObCC0LHeggUJ
PZpu1Se4QpkxMCBvmYq/SxsxdCWl+CPq8NwINCTpv9lVzcGzxlZ7KUubNGk9ZsjH
fY6Pcol5r11JVHVk8FvNly9Lq6/oa/ty1aNnqG+zQKDwyIumrg2nTJ3X+0XxMLjM
1NgTkmROQ0AViSadywheuNk824NiAgB5g6DzGWoXUfLfj+MHXUSxDSnYVMu86mHn
cJ3CojoL04dXwy+QZJpTnRFJt090d+j6CRj8L2dRab20L0Zd3Doweh8I7jyFjj0g
Zm+UmhWeEXiqZsxQKQsZFtHywNyCEFAdst8TGw+SroOKiRggYNUZJJkQGmvfSsQp
83umMwaT0/OXtqU5LOaf4rPSX9BNHj4vnLn813xkvGIXX1jxKRByk0h4uwa2ssyA
p6uGPiydr6t7nn7ERZDXdAOiAsAEbRoyQV+v1n9yix8CXDhuNkhC23dBDsBhPUrW
cuyWbEta0nR4Ul8bpVUAMfhgWm49P6rZbiBub6G3KqHXWtF7mb4SHHG09CgU7syN
jckoLG63U95wRZH/ALHd8CUb+RZqCgIhDp9OF8TLOQA49fSV6lzr82COGQFg//5d
KvkxvHI6D17YW8N6ymcMgUQD1u6GNGWOSZOFjWTFQ1JjC6IYOthpqewOCwtclDzp
jdUMV3qPvKuNzGzoXMKxVBRuQayYt8TyhXm/QAL/QZv7Z4dgLfnBb5e904kGIne5
Xr72QiPbUhE69DFdmBh11V4c0sLiAYo8TLshGkRqBYwZML6ZWxCZBQlQ3UxoCjeA
ru5PdwpO7ICM4mV60I0uNULgEG7s2xhbmITPlr29b7MzjjkZsDiaWqhd8Z7BrAfj
Xdmq5EpVxzz/9cEwMjQn9BPfKa9rmZBWoubvRJhv3hmOWW7Ph3crEu8oD2nzOO9Q
Cu30c4FVe3NfuI8XFVUJ2ovz9DhZcMksBVZS54cjCsl++ph0qdv/aRFUGurtA1Pl
e+XLOrvp/I/0v0ovec7K989mT81Q/kqDvz78y9uOF3W4+IQWpepvlk2W25XA8JW2
KRPvfBCdVeoAsr5Z8LxzvxfaeNwERIGYCbfNHt4yPxDwMvNl2EJIU2rofec8EqpE
V+zFuWCPnhZQpLNDh0LqutS/brdwLkWdH1rcvEdfgFXAohkTl2Z/LOIEOIMnB8CT
SsWbklCda0hZKCSc0YiGnpHo61H4Ae1/9OFXSudNrpjfmnlenj1TeHd8SUWAD90G
j9tJXGhtnR52998g4BjheHIjcBP44icXCiwoSqwlS/U3fgP58mMqPUbCTqSNi+4I
T9zLzKFCWQk0siqruGDC9C5YAQZWMtZ0wJGJGIctcF4dn6CwN7fleOux3JMdYm95
sripvh8lK470HKOJNZR30bwa2QKjeuzFyT+JeN0XELDg65/lMlEcmZOq3cc9jbOK
BW692sDeuZwSXMYct7cIWjksZLU6mBwPaFU78718gIlcVtX2BZJrqU7cil0Wihbk
GLj6ePK7rCPM/zAD8KZU1XWmgdAG8mEstFydqbApniGLjUTlNHW2V2Z6CNcRMbn0
v9ZG/powxtrCHj1CkB2jrenF4PGvqEEkOHWTy+VPciQq/rUqAKKp06dQy9rPvwEJ
F1zEgA1BfhgnMx2D4FRNlCmIgMFpdZqnO1H1qfyJissTb360yAPvZK4pqV29s4Tz
IJDiqLECBWosPDqaLwezKb3RIJmtj9W8za4ke/xKJ4FL1khw178aR+aHQW+uIn1c
vDSQdgBChXbrOnNL0U/tRx6uiXIB6fMr23yDXLNmbTBTSZq+l4PPYbRmc1abaQo1
rMvLlRQ5tf6z5hbDRAlPJ7Gqo+jP8Vu6tAUsaP5OQgM2gImVM7xn7kP8L+ZpM6+j
46bFjS+VZ4FpgrZ8FsQmnhjfPSJRj7KQ5JU81OqcB5aL+eqCCyMoVn8rlALLETCv
gksJdf32p1zvXhJszSvazM9Wh+1tBpOYSsEPT7+FjP67REBcUdAtij3rO9zX6GOK
bzmy0McaBoIoqUB5SVvnHwweoadPbm2hZwA/BBPTFMzwdoDtAegH5M2Wom2/9wG0
+e8vMzk9AAvDVD1TQ78Vom9uBZs6iNkLfZgOkkxg2knzRJWo46xmFN+/AeXLKXWd
ca1LRnbXlnAHYSE5BQXQa7T5UIv2nW3CUDYTGKf36rAdgy7h83D0dQBBKT+BEcFE
8Rjud/8vAof3xuUUkoVJlgPNwX6ku9kiV66u1qYCNu8cEpCbJonp49PHFV4myXZM
IetM7H8beo/WLq5cVILFuqmBIvF2aUFtME/DF0K4tYw6YUNIqZiKfXVbo6I8zXTe
NFouo9jjFh1crTMOs+azpu6SzwjpOgagOhxjsdcToK0KESbVYx4tUTN/uIWsLk7a
up6CFVZ3TAvfXgr7+zAfS0sdFcr/t8NnHAqV/DLa55+W8xu8oXwoX9F93kdCvumz
BnW3A0NV0h+6wRBYjQ/6aVIRLFwLCOcwvU1Jz90GkS8abdogQak8aRJyfHGd+l2M
57QqiCj+rew6Dk3DZltphdoZCwNVTz0GzNA7ycl2ryzl46xMkwzL5xjohCVzdm73
UOAFFBh12Ei7ZpHsKhVNgtVzH7HDUb7Q7DABPjEASq3l+F1QrP5Z88iwr8+iMmmI
XtB5Q4q0CO7vOZw+WHu/Y6Fy1NC6Fofl1Sku34qyP+12zLJuOaNwVZT243SAu+ww
M1Hvl4a2wd5Yy7kMEUgbNeWJ8m7BXtoG/o6niFuCW6LsI91FYrDLkfbzUNhei/Tn
g3ErxOnvfwQVo8AGbgVOl4dLpFcMIJY+dg+Yz2bqdRJJddjHG7Dn1TBLTemeKiXV
m9T/Zr5ZLvHOlreNB8xgrXzXcdWdnvroYe37Xid/14nfb9wBaun2wvPjAi8kVMZ/
VaPbIH8IiCRy/WvOrb0BBKUIpfJzrX2t99pEDe783rGmAQ0k4iYfH7+DL4IDhbqP
XhneQSBgKlisqYDBBvynXw7/DSEHiWZHnIqcH2fyU+To0uxAQm845zjGsawSOiyL
TvoydLNExBW/GhBPl8CNf377EHuJSTwVwdldLE9EAEa79kctKzfBj/yx2WZJif7O
Z4ybBKbXZNhq0lJTNkW15PZMWaYU3gGc6WGX/8nhHYWmZrDbHXFpItAWEKCFxuj3
dvtcV1cAz9BopeqgDSBa0IhyjaO3AazdHw3D7LPMolIOKnAUWB8lGGZExhvXxQ/Q
MUSO0nR9QgkB88tIfVQB+V7qNOTm8ynvyUTX8NVr4iaoYD+u0TUeeIHHtUF1tZi8
KEjb3BSJeyyt2bG1LMvstqznLKbbBjIn75+Ql7Hj7SJJbG4LUfHTL0e1ssI6tiN8
fy2IUk8WkmNz1hiMp3ub2fBRf5yWn3TmGNf70yVN3mZKTLR26OM9hd16WxwKOcj2
JfKbz6hGVZ3pFkpe9Ia6llViDA5/R+pdZbaWIq0hdAZOvvhDotJ6d8Az4EI52NIw
lZf99m51X+GpPYUXUrp6mAKQ61oUtxJBJjb3/3L5F+fllPzzP72ZUHNrzHhfVpCf
46mkIbJS6fzt3CkKnYK+lZFPhPOUNaw5zThgUXmzr3SKwy14sl3vNS/b59v8Pkpt
Ym4Ge8Ou9wdKHopeFzqrqvIZKZewzEJWr9t3jKtanlaZ8mHw6vYqzmuVGWGdQas7
kX31UbJZ38BaIeur5lzHF0HavbSWEGw5na9CXkjvcty7q3pU376kSU/ng4c6u7iP
SZXh9ne0YdI/kHxQnkZJopmTaTuzMb3wozttC5XwF8eqVGsXWAsw4LwtyS5f/LNA
e6FJ4lI7DKifEuDdxEkWOGe5hBvodmQ7q+VzIbBqBufvY7XzlMh54WIGkAaWFJJJ
tyqSOMn/RYedKtu5HqeT60aKCVQGK6huN+zpl849PnZ3LNcWewLxfiCQZB+63EkM
F6NfuQYNanq8XrEAT9a5aL0G4LZBbqNPMKiWlV9KD+KBWJua6hFVT9xvAnf4LIbA
QeIjoHdNDC0GKlTTVW4n/7fAHiVTI3SZuXopNGVg3kDvfAj2mZ2VAPnaUS9tnH50
7rYKtKMJPhf9UVGWKOYmTlEE/cTL7etEf31IutSuBTIK50yaFRT1PUyZHrjHDP4X
JODPz/M5+BIJkTopslfq0Vv3o5ua1AYtVrqtXFkwd6Uoz8NWDXDlQchf3+iwe3dQ
rYkeddsRngX0eDU/7fxxgalNqgZMvW7XgwXnQngXOnc596ltjnx/zc0JkSDkVosp
D71hS0vCZRkH151okUrB/wrZWxXM996q+tobKzIxKsWGhN3S2Fo98m5Cy3gmYytx
9zFPtxvnmxGvqlGq+NaLe6xXSte/qX1M5UqkZn4mdxHWKwEtjL/2Ojf7XJLhHYg8
uAqL+YQDuHCuYv8+1EuSlJNNQ3rVTlD2JjUvNXanB5TRij2GboByZhBzTWzZq1Wb
NL/x92hqiwiKUZYQgTSqUmKBDuixBvIj7bMukrsvV0lchMev6sRhJhh/p1kwmmK0
AcsDfOqCh7s4Id8GxhEEmAOnLkLvshpoAEa7/GtyNMIQVtrm0Ce7YLJhsQjhZATc
lgkqObpx1V424GMxqt5T3+vv1RrGXKQ7KL1ilanbqiZq8G7UhCiX89ygW3xVbj+F
xk9PxPHBWYJqbWwYSTjbEQZnDj9wsbd7ZoknN+Nt+8i49aEGW12wQmIWbFkFmBBx
vRMWN1DrsEHlh6P5pRYJXyjeCnIU8+UfPfCjOwvHoA3wk1+pbBcBMiaGVKuRyr7F
Y8qpKi1EnQO/Sp0UYDGsGSMZkTg2QYgNoiJV2fId2iqUnx903WxgtgakPyCHVfaa
l+VV+AN09rrdoniZyLc9HQkFm+naN7uDZi4ZQztUUPo4HY+4DT0qFNKMq6//DCGN
udaxlSfN/AC6tzh0m0825XVInEcVeRhUiw01RFgWmYnV0HJFEgNcVdiS+7YXqnRH
H7CMylECcQjwgxH/MUNI8MoHjFnSDzdEC86UTDAkCJ4pIsdcE0dRe6QmxbK2/kHH
K8arjzW2xEExSQq/65ZnglbgCp5xhqnsG1wIa3ob578p6KvydV171vy+V2h7wzMv
gUTZANNGGgUM/pKuX932z8SU+0Lkht6q7dIZ4fo+QStJ9Ub1vnvrsh5UjWMxMBVM
O00ydU2VR3VA3FYgNFB3aVNcTziFvqD70cW7bvt/uBaiQ4oBkKDKHsal7FWckXv3
3vr5rM/HB9JlIyCvCMqZhApP+yUfRnr3xKzNIAyn2H/bmLjpVF2nMfYKal/WdfCA
grvgQlYHne8MdnqW8p0uJqUEnUUWKVddFvgRWA+4jfNynORCGVNHwkvPkOyOo8Lq
Mguo7ryV175RmfX3fLpCDR99Bw41B8UXIHpiL93cIdL5k8Zt9BW0Ihe8qhNcF9mI
u/Fa07fMTQsP2Ts5i3wSINp8oLJwEk5CrYZdIuIZiB6Rg0j4/KD/T/QcIs9tWLHO
aPCPP/Kwc1lK87qhhcHFck+UVGq9vA30yeZFfnMJZJlEBtKNL2vzpSZfvmb+5174
s8yLZjzuDuO2n8gAkYfH6d69ah9FTCk9JBvMKx5M6LcLhAkNIxrwvkeSnkcKKN/u
nb1+9tEAU6NOJCchcjGrmPTxA2TLJ8m8vCZTTBE2WFeUo7zBFALAKI29b/wlaUHG
vgpdVNw0WuvWaKDrD3M6EC2QDuYcEWu/qx4CaHWIFq3Xzq5BX4jQOjk/lNRpgh0+
xEjp4ldrN3sXD5pfU6vg/KAro8tgO1hzzafUGiqPOraEipHemTALED4ogsDx3GyQ
YduCHPZ+WGla9lvNaHzGNpyHU+jReMFlyiS5/YgYe1Ka5JhU+kWtfpXvkOWulNc6
R13QrX1G8yjDeRTuEwAIujlk+9zqVvu6vb2ypeCfzCZjo3wibSOowJ/EpJQhjoLU
W2mp9q/dNjgLdr5/1XI/y2q8kqDzcCcpJG5Oc4rDz26S1HQ2sGkSr2qidw3n+Oqn
cHOen8zshAY2rDyvnGsNryjUm4qEYu4lxsgZPA6AFcItnBJhINpmJnd6WD6D26eh
xE0ppBQtavjdcLmTvGyynmaWcp95/Yl95nR4rnMJlxRnP99MPp55z2QLf440EkZu
FuFGGGcHRgMqw9/AY7jt8JoYzjF4qCYSDj4JNGRBd7AY8Xb048UCdcsiPkG+V41f
YX0FMrBlOydKMq5q5SuDHhuKbebgZXETTt6FI9z8V7dXi5dqY9yj4nYivoarFXrM
Mguw+4DtFa0gSUfr5982JoMvBOkYTwzWKb8tf07h5z2rMYtjrv/YSeG5zzsLqHo6
ejqFqfpwySfmwZeohXiCWZdp4oJIQY5dyzvzLV4P+2GEkVBaaeII9skGtrSs5vhW
VS91aljhoXOB6rvGss0B6Gp0sLVPjBwfPa/etidX4Ig8c71vPMCo8gv2HrajmY4b
ME9uRSlrE6Qmff/C6OUYVdMTi/nlveEQTr8VxlA1Ft9ADWyhMU0P2Z1O3I9M4Km2
vM/dgOk+khiynxt1T2KpJLuoKGqHPtd5A/8JgagyhefNIBzcfSXUxh/EbO525qMn
gankV7GP5L7SIxkmO6+5skqsYiXv0nWFgy90DVaePVavraXrNfEK2oMLVlSNvKs6
ZfZcvpDjt84AX74Z6ETyeHoC+lSeoUsbgfQIRdyiALvHaIClSs6hZyMI/5vbxheI
EzWRNdPtO8cFJrQcXCcUy4RLQOTbJmVbjJOYk72B52qpl/AYHreWeuTE55FsNrDG
BA6Oe2iHs0U1ck5jTKUnkgzgspRuMCLBAQkDm/YogFmMFX4KRQGkXHr0sSplM8dc
uNWz9mcWKV5O1VYu/5PsDRdemV3p62497uJohXPYxiZnp1mywcyPNxdCp3fcJlCJ
4g6Eoa/YJoEGt0boo6c5f2rk/xrgcb6VoLIkz09KakoUCJG+JZWTWnU5k9p5KLrB
+M/G4al7WqeWh++QAbNhnbOox9rM2Ipmsk2ZaiOuQQuNxvMrL5cRiCEU21jCIASE
K/vDHbFFG85I3jq498SOmAOj6ZmgR5vfyc2cd71voXii715JQAUwVvQlO+5ejs35
yHgUwK1uDY1pweYHFQKi6Kdpkw89TY4dblt/C+qlzRRkSaIeku/zn3aHUtNE2h/c
ArSItZHgk3OzN/rUqsmcU5RdIABitfN+LlDqsGmRcScImk3LhOKBlgPJ98KV84Cg
HOBvHlbrR1RXZDHsGbun2vDD0Lecmsf/PvD8Ynf4v+Sws9xZUBxK1DeKQeNStBTJ
7pU7h/5fw/GUq5Ifw5EC1Nb63CxMf0NBT4EEvOQzx5QXusNkpDQ303ZPih5adCB6
tbbGbdeSjoqssYHbx1bF5dzSznXBFmsVF+KE2AzFFTJ0l0/SyG23qXUgrVrlzSSD
hrVnSWd7GTDErWcDzqap5I2cl0Eele1ruOXxXTrKh4R1mqAADTgDfpaHTUiKAMrx
lUeDIuRkFM+V9YlWj9Yka6V1I5CyEutT6Y1ov9iQmHWMNaad7g+HT/4zK7jLDZZh
Dw7wdArWfQnA9u8tr7+aSq2tMlUIRRHiE3R9xboa384awaqK00wDUfOo+kFPlJpQ
p0W0EQjpEmpDSnAP3tv9KcUy93mtqcV6GF6fzxFVHn9ANgdkx18NgHnfnijfHXPA
qQ3KLmvXwv1y39SCOgGAFPDVaJbdqbCVG5x2rAe5NrBO9GKxC6/f4nV6mmZo0FSt
WJgcbpKN0zPEtG+QXwQyn/mcPgIFdimDEy7mMgfULXqOOZyciAQbOFNTPghVIqau
FVp73sf7oI1rpTh/xIsUVVcaNAJ80ehUqKCe9vJAR1zFS+8Q6o5HlM2xjz6Q0i+o
WmWSfeMlhhgEDpgvrPXNeB73qZ23XCnVT6s9/q+Q7jAs2G/uPgNXHpsDu5Z0LzUP
n7P1NbJm2Mub1XtU8Pfrxj5LyALCX6X8BER4zdQRFArR/EHiUINvSSGJP7I6W9jn
xcNsEcMjRsqhudqKsq/KVEaOLP8Sw6wehHh7F4L3+gt/8WcV6KtU1+aNnXNm4Pyq
n/uoto5K17poRvw34nshPN7zgwMyISv9CoL0Gk3fVdgmhYMQtXDPBE4scg+mK8An
c+UNFpKNDnQhKkGiENV3HzgX+AEgLQcRJ5L3MHWq57P+/rQ/uvXmLqP1ubLFh/lG
fpGti4L8CDnNq6vm7MuYinipTZBfWSFNUD7vtmnHQPvYLU+hROmoUMj6ZyP3CLjD
rNvDS4dTQ8fs/hZw+4+G3T3IUuoNZueTUG1uh7LNRVDgxXsbxfxy0mFUWECKNW0Y
smCzUCFyln33DjixrLiWM0KDUPHYV751UCyGTldPUVptWiCYnjq/UuX+epzch8aG
luIxvk04iN2gclQGk3rRD0C9jsCuF78FkjXzgG1u0QdDdgxVI3NMcE+ktcmPXxhr
fCA5qbkJkgxpfj/QHaasz9ubz8oQncuPIjGy6zQT7HRbZ0KyQ/KJzoXx4VL3z+oS
NVmPWK/aS9DWcvqDVI+Ofyplus3YJpdzilws61b8O23Zi5hbRGhCFdq18aU9OENk
J4BWx4EhmohFWokbtPjlcB74nJQs24qfne7NMhx7PIoMcHekAU7ZeKzOITYbIPhs
kTnuysBAaBzYtDbdP9F5jnYod4h+L2fQQrzEmygVpffmbP1JG90Z5Og0eBkT9ocR
hRGSiFYJBF4soqf0vX8u6O4H/H35KzVqjq52DVUf2kOHEt0h7kays4+yTEBt+VPB
E4fMuQ9nYZRiPxHWGamsujh3I1wrJqP3i/ToCcTiJywch6DrhT0qtCRbV7zOK8T5
L2OQrsuk9h9g3i/vb9I9AtKk/7Cy5dJv6NxHE4EkPaIVesMi/PkVz14/67l4C65a
R4u2u5xaHSq4xzQ6Gd3N2gQfH7xTffvmDzgyUVbTLz6d+pFA484QmANwyueA5sYK
RC07h+HDUwW/1UjzhFsr9QTl1uiy2qUXCICjBqOXkTa25Jfs8fcAhC+0EdZPXdvx
0GgI8l7FWjR6ZY0JZtI2k52e3Evld77er4s4JiglLvLyMe4+h8NRvopsCs/r9+bJ
gFnrs9aq0DfXjC64uQVTyGIIVq3pKEQ+sBVmoatuGvGutR4qGCFmlJNwhxTvag95
P02eTljVA7KQTMkOpl/NurEWN2PgummRCLfjbxcnGsPn95svxeGS1GsNYzD+b7l4
Ry9DUID+CC+IWHULEDpbNjSQs207DDxBEkDZRdZ6WbngzBIKJA/CUSANJc9zimko
mZhntJYmSWr/94jyPMuCjoaq5kL9488qcw3R6dZ+4qXB1aGv1weONqYNikBJ3Uou
HCWr/r6ISNPDrq/Nf8Y7O4ONIooxyBMjlEe94B8CKLwYMr6O8wrkpOktzXQFs7If
CkLLpI/+tM0ns4I0QjrJ4YboSHK4YBSZqohn/oWCITNYsRzsQ3ccwVUdb6Zg5nt5
x6tP2KWXPsXG5rsVQkMx2YejInOe8jrdV+T8FZAUC1qpakUpAM1077KeAgcaKps8
jYHMaCEcXCE3Kg1w2st12dX5+Eku8i+B4ZPmofzMfm6lVt71poUS54t1oPQ8yuk3
jU06v/w/0phTsjD2TPMx0iogQtbgggZn/l6RTG3Oz8t2E4d4OXvRAcDP2v/kywWj
iLDc2MfmVm0EYSYV7r0deQ6/xO0FatP4VNDC5S5U8DejTTtAao5ZfGEJ6calkCqa
XKvD1hbZAudrywKRQnbW6pKKyom0HXC7LqIUC2cbImrVmIyFMI6Jr8SAKXax093M
nPezebuYhcYu2zcHt5ySCS4TYu0xGRewzJ/UeNSfS22hyyzLutEUeKlTd2Lxs9M3
hbpX6TlVAiaPC5SgYHGlAZgK98+4gs0gifFyetweda5zuutUUVc2psM+KW0NDVaa
V6wQPH5kJjmWeEmaeEYJg/A9b4xXQQz0wdjZRFgDrHYPa/Q6pO5M7Gdm14F9aQSS
LaIxQsPylt9FCv/p1ZcAgHDF2vyxgbZDDtGKhf2zDdq2D18a5d+6NHDWxwnYpejf
FiHMuz3TLqCJklJ76K0LEeCHbrmpkVS7/5yc2rnNGwSuZIVZ/eLDfXWtiS82xk+Y
a97iJoLN3Cbdoyc/hQIWToaigY+OcSZ6zCoVlJVC4cDmXcSQ+qr7xRHYvL2EMgGb
QB0hN7MUndbyCQoE0OtFKYgdO3MxbVzdN4ysq7z7evuZJF6D1J3M4lXt4OJV1YRH
LFNwgE4AF0w6gjxpVdfI+EIDMgqr9vjC/j4qoOYi+tBRlBypMkYQzfJ+iUOkSbF7
HVQ0U3rkf2k6BPsukkyIPGgtRKs1LfJl3ENYi1ki3z0F0CdD1IChYXhbaoqfRFqe
aFOIJiuF8EI3e2Z8D2GeieoDqFRowcWOKEVCc5QRXFzjV0ZAid4XlF35LpcR4yFp
BwfNuVqeRNaHuVsy2LgBgD4dBZux8+embGlVu1YmnxM1lDuJaaZcBA14jjgkeRz8
dxuimjbLPySTnhycoiExsJAZqdAzkuAxBCewLGI9Yue1NuJr/OMtpTqvSBokSivJ
gFjgGeL1ZLpQQGLnpbgsF+GQcPscKvQSbKSY/4ZyucDeq7Wn1ZKUK1FRpyYyrRbc
vGrwpCQxRDxgawjxKn13UjFdPxqH29Yxgpi3hJ+WYOrOF3AxLxCUh1Vo76eK3mjq
25+8T78nU3vcVWA7PU+Zzccjk2hgGdm9Ypxjr77MwUUtF82b7HWfmNSnP9mu5yfX
b2medrImqxDYGQ3M1WTOLjvtFM6woHH3xPXxYTDMTT0/pIDUCKKSmH7IO7iRDIiq
perOkqqabd7X1c0BORDj7hBV9Lq64zKU4yzObGkxjvdcGkbXl9eXok/STigeGOM9
f5AETQzgIuShMtXWPUBIFtJ6rcTYDHXpd1XOZoV49ll9QJF33JdNhEHVnr1p25Qz
cQvu7vytc9Ghgf2XmLwm9/0RNlGr4Lb+yKdsG+F92a3XmRO5Y8Dl20/vQiO42EwL
yIkv1zQwYcm7bfYrlyYCWytvAjHkf7A2yrg0oYPtV2lKD+/6UmZ0B82mcVucbIvS
5Ss9Mz5zyD9vFn0qNX0jD1slDTEofn8aoBrs82bskohS5k23TO92KIKytSkocAa4
ukuKXX7ivKH3L9YzrmxuYQ2JWd1JVnsCkbubZBtQXzOBBfwowlM50CZxBJ4aR9KC
87tsBeR/+LibSks2nn/yN8UOZFUTcwdt/jO5P/aYqtty0tJGYeSK7nsWSzgl38w3
FgypXud8Sve03u8NoYbBBmsz3tgCvi6/cZw0eBtvQfq39tX64gqIbM36kDIL22u9
/bpLRrSMAfZJhpe6RrPCz3s249EYpLzUF6iiFfI0QGUPs4Uk5i6CXWyRX7ljZdXz
MXq+LJBPwiY1OKmrW6ywBqTarmvQPsD+eG4FVGM/5e1NOpDnMJiARtK8bHLAUplm
fc5fk4cCxFjQDH8xqZVC9G18UcVJvmOM4ECWuwmtseNkn1WDzfEEKxIgUskSXfe5
9MM5qHJxwbmsrcPsQSVRZzjbH5gB0b8DllvMutzlRmLHi3SJEqdaub5PZD235FHK
mHisMlBdEaTOqSVgIH0saGoHm4RlT8em+CAUunmTR5pRkVHDmxyYWxS2+VflqTge
DfC/crrKQ2sK90zY56SwO+dDLD5cBfLilg3ShaDZQE7MB46aNscxib8DeesgEyZT
pKrcEIDQPRDu2+MCfjlccGJY9ROgMIVg2R8UNM45/bNtwlmfUJvI+MJHZXACXDdz
eFj6l5jUUhJCjlHRu1t65lQa1QRueNf13cwWtkxEep1riNKu81S2TW0OzEJws38Q
eLVytIy2ZwKGQ+bNVmLTZTK7FW4Ht3D0NSRWGaNZgXQ2yWEQknykcYd3UdB0Xkcr
iAu/ra7JTe61qFUa4o9SPDsnRIEjRB8aFV8vVWVmDMQUoqLjDlg7D7ah6llYsUiC
G29hn0U4SfQN6FOhLKbEcNIQMTFmihfyQzScDrNov1XknFW1A0Tc71bQ18ylx8dr
b5J5Fpw+pZJC+yjA86ImDYBfPGh7+g9/5Ym85SE+A59VhDk5yPxXRHbMxh0mcqBn
ewxNweudA17g86gptYfPqpw77nnh11jwZ/Y+7jbJHgZSOsVOM5VBvamJU5s1edCs
otkJK/Toz6lB1+/llldq0yIouhtncJGSz0XSDUjne9om92eEisIcQcRlj9t6tY79
6CeezSS/gexAqjUKxWC0pUyBLyd3LYkXnt/WGiC6b00V4399X5cKZBRXA+z00Myd
42B6PuNIv0pqsvAWcckL2twn+0pm2RIY4TOxvInZccZRew4s/X8yfc/d+KnZ24n+
GYP5gEX7MrMdvLQAjFlEiyTbqOVACpRm8ErQkVW4CDKBWWGkuAq59ZDF131KecNY
rbPwwubEsTrYKh3Yf3I6MAXM0wwksbNYsMc/dNOG+wWwS90uoBXuNVfknN0Ga4J8
TNOJjVnBdEK6dbTBoJuYM9UtU8FsOCqB1svxstYcT386RPKSm/Se9qudE1W14yWv
0ViTLJYzOX2PgRrZyPN5jB2Rk8p5m1RZbGoeIUy723ca8li2zIOsFpyuKGbgoZ8F
CyN5jP3euqn/Skt+hsKR+j8mnTHjcb7Lc+cBjJXNWtXw8eN2UPyyv77ya/qn47ds
0rWj8DPzR6pIm9hmbFp29DYkphHGe+FOa22zAbMPNB125ujtFyFDlYfqxNPbHYbi
E9cZDmZ7gwwWPNzYNF5u+g6rF7K4T0SmGtSsEeq5RdOfs74Wc8CkvrMieiTYEDk/
M6cZdReqqT6Gi3TfDuZpQd8MeWdgugRDUnNLm6qTve2K3+jF3kkTl6GIbntvTboW
9ewxBipzr/XPbrbjGX8H4ZAUk1qOK3oSqTbl8XOfKIek+RPRvIeDHrpehKNM8fLl
nRE2MJob0Tnzfw0tcn95c4ZxQA2cz+cPZwd0WZCrL4+Gz1Otpm5RUWqVju1SVGlB
4XuJTpXsnkb6i5mm6009UHdlJIa1uwTGeLmjKy5cBKf3twrFNY9QjqkwYgFA4+Dk
f63fZcJbr3JJLvUD85LH4RqPGODk1onRGQwk0Er2iX332thIT3uLQisIqsvIyGrT
NXei//5RW2LU+EBeA0jOSNaS6y0R8ABhWKlfgNVWCFDVrqfNEwL4qSF38AQMj48L
AasUbs5ExZlek4UdijWeljv57paIHurQU2CI/bHhSDHE/NrpXWk7SztsBw0shEcc
cW7SSGqtncfAp7UqbbxIb1vJRjzwTVqQRkWbmfoG+lGBeGzbqp3vz2G1fogNEX9T
LxEr2JAHgo57z1ZE88PgFek29UAyoe0A2G7LHZCBeWZasyWq+onKg3sxWoAXTLNY
w47U2hI0nJ6x8ckMEy0veYnaGnxc+dA87kYu5C0tlgP4ulocpIRsR/FbTswghaBt
h+CczSFnF3d5jjvrzm8F4XwdrtKgwO82oAda+UiguZ36pCULNHwpzC00j8perr1/
olOlW4CdsYWZBzC9ARnGwBqqRK3bd9ZwVT7voJflzENYvq3oRiWJmPHgZOIvkNxO
pzQTiZLGixd09Eay+dHn5AsWnnS26SdazDtNAq6KxR+4N574/8cFaWLPGaTLb2lL
nzXk9uMU8vIVCUh7WtKiyaNmirGazM7kCXtfSVPXxoxzvLRtxhMj9Du9E+gO5z0h
MLlWUBJdJK52SSGPr9WMR8i6AuCZj7iLe994rUt5KAq6y5AE49eMU4p+REYNeQi9
XdRqiG4Sr8do7Yqq+daMazOCcvZac2YZOPgoUK1SYpRPi6fntlmYwHMjMYHoVmyP
pqM61J+j13OkPNqeipKFqrwWgdYA3Vhvd/0Pd/5qBe3dq8neLZy8A3upDc+hzl5F
dllUc+na8u7/9W0nVrN9FsF57xl08C3XM/hVPUrzHrnjfIC/Qz1mVibbjSoCFMIh
WSNw1M7nexmq+z93PQqgk/nX4VVohs2wdZBy8pLo/F7b4JIbE1B46xBToLpSQEfA
634IF9K1mfnjXRotEzje0y0QjKyr5Hu3nRY/c+/y4nVWhL5uwe39ox8ukpvNOczr
X7dpVQXrBrcwCJvqr8M9c8/tAUJAWjd32HajfmhLnOaPdPtn7xQ6oaPraA1ABeGn
sgFMmKEeKO97G6h/j98A1bWViNV8zhaFUx4AbfFHEyGtc0wSvcHcONde8AJ2RK/b
PxLsbRqt72B95rgy4JF2uab7y73GTuCLUqkKVlv7vcsoka6DmL1QIthQNSslGLOc
1LleJRBmPXODCK+E1/3i1v07ZzO1RoIvjP0njJZi2jSgbYheOsqWhgTH0uG86ot1
iKayXjW4rNbrKj938R+o0fgwAO2nDeEL5SZ6ay45I/EPG+ZVtE0F3uBc/vZQYtm6
EDVjZUyhJmVwDYC4sej5D79EhHvkeRNATP4gl0OJoqz7TN8OA+OBBv0auV6n9QKj
orfh0rTtegUMKmPdlqT5W+jO21j+LdhyOsV1YF/cJE44Or2Ts6EoPEJccLJs6G6L
G12u4/9aVpZ5pC1xBo+3A/PVZB5PLaavzq58rxsLOnPqVOjsCEc6QVOfDkfoI0GA
U+ocD5kx4LMe8Y2WDH32w8irGNM+R/bOrJpI4viOXJhQW+3v78FV0DA5OGPMIB5i
D4FdY21likdRPI0ueHP2ngJ6EMAy4o8+GcDE+NZS5h23N1jovzqNaYpYXcDdyigI
XI1n/kkNVwfsFHJgrBmlqJ3tTQ7IEnPgX9LO4Y5y6ZL6c4UwlkU/I1GVmSgq7kd6
XhjERdEBtw8iDW0nBFJeiZDY1YYczIDFOtQREAIXnBoTHrH/7pbZ/4zp1QSISCak
epD6k52g9bRliQLtkewUGqK5aiS39gUyvhLDcfQ6iAl0TPJyQ2meFYjYsN9QSO1a
JtwThdZ/5HXaLFb9Qg/m9dvYltz3is9A9xzawB7qP9Rr+xX9ZArM3aKIyRJAciUf
gcOjhjGrX/BvARJN1i55Tpua0eBD4VE86Ppy3YgsKSm+XLKMs93e8ko3vROIusl0
OXoH7l/q0D478FZ7bOcwEs9kVgCgQ2cTafn4JdVgNlgsJJoabkooqqQS40ANjZPo
pNfGopNxKvfx3Mx2ubSztRdNzm+L/TV4qZbbnU67/7HxgBfCaKJrWlVLEcsBUKlx
4Isl9dkPclF7expO4Pz0+Zcj1yUdjRpmydmEeMnWg31KQCIs3Q6i3gLnBJD7/yGZ
9YFbkG2U3XZiQVL8sDtSfKHkplrdI9L0whp8sWWlYtXsusmLAOM10R8f13n6Uwpn
oTnoamPjvdH0KPRM9NmOofSUeKuiInTLn+bNsUByIBFXZ0sIke9Oo501aBxtx5SS
oHVt18LCamy1cM8CPdg0XS3FU9Q/kbjmMJZdfTyc4fMa78S7GS+0S/NVsGLnl3Sw
QUjUYJ87RxB5RoyJPjXUzfaimDCIn4ffyco30yFqo4FlQEWed2ZrZtu8qBYRQzvF
IYy0F5CtUkFcipbU3C7a49b+/m6IGBMadafsGBWhNCIAK6VeEHor3YGyPhY/oKTe
DpeCCfp0pyBJ2+05T1MJLPbSGAmOvRH3fqxTLAs3pzq1DRKSDoxAwJuNWe8RNI+z
c5PV1BhtY2QanSmcQVynrUWUtNN3Qd8TBLfQz5zvRdCA5U94Y3YC6zDiltimxuQz
Arn3YFSguPZbBL0uH8vEasc9aq9UbyFtmMbjlh8dlcvHuFrSxLs/KkNAYIaHsDuL
0indX+FMo7A+dqIhamlOOz1w1AWtXSDIqRa0f8ld64mWcpI7KvKFVqI7R7juzHuv
0dO0yD5vDBXgvbFl1gqspmJHrFrJ/Wwd7Gf9UsZEGtD2MF2uIVhvsvssUnaqaxfd
00SsDcaX8tYc5QHmzJmCQr/poYjWOJ76SxmGykoKpU2Bdhur9GMalkW2EuXGPyWe
zhGVAq0ASt3CKhihkk1J0Raen9G946Z+ikUYHXBApHcwYY+UgG6EeYeR/YhFGWrd
gJ3i9OeHqhVS57uy/XwOhIQtJE3NT6W37Wh7cM+Q0Txfldx7x1GEjf1Sqt6bm+C8
gE3s1gQDUzHG3zsTebh0BCDHBjVbBKO12EMn1gE5ilnfVUYXUyCEmbJgo7h/wV0x
ud/J2lS71R0OCTBkiO1ZLGy5FnU/sLE8rtMnQduE6gXlioixRydCeTshHAb/G10t
C2tZMOnf06/vpBFbiEO7dtNFByMC51V1+HOgDhsRML53uv0oQzSo6/jfHAqqX8VS
h7E8T3simJQ1Nn+J1ybyzEf6FqfFp43+jYSGjLDUf6BcOGx6bZ6RWB2+H0bPKKQ5
XdR0hswSZP7+K0KccEafEjbdcqCtinp2QKusj3HtQWQmmAQJTodFRiSoo8Hi3GY+
kg6jYgRUJTl7uEUP+Aht2ySoJYW+RWDTSAc1Bkx0gVxOG9lHiDRdeeGSDep2pRC/
+O3zusJaJ7CM4+BLJmH7Z5QlkTNK+pifZXPdWNedcX+BWB2M6bhUk/FDmLrcBfLM
h0GME6s/WVewGqVb6MQbePIZM7UFrCSTju9QS6NGv5wHi4/V2RQMqxb/T5ykA1ms
ALg1xdleLQ+7gGRd6cz2GKZ8juauPPynj7YS+vhJePSMVkzyd7W6Em0E2G74z5mP
/FVKfPWupxs/INCdb45aDE+ryF6G960G3wmzRs/43EGEJEeAkdi8tQL61GjldOVI
Xa7+NxZzO0/Ck2MyiDy6mu5pjioNGmCFeiyHoYShsKbQvzeeRrVJHQfq05noRkEC
QzgHHtuh/qLXlLgof//vLCGB8j+XzuMdV6cmM7Dfs8XfsZ2DWi4j/oZp+ilQjfwm
EtDHYTaGF2mEYzwJWpXBYl6m6ki+av6eb2UNgxKXP1HwddZmriLNMHdYJe4FYTes
w2lI0VoVc0geB2/X/jW93OIXyttOurX2OB4dXwDej/m5Tj0yqatrl5k2O6p6i7Bp
0+PjhHAKbXiwnPnYlweRPA3bykz7eC7uehLWTjFmKpAvmAFyH/k1fal4qRxZBDhs
LrDh+Fhvb16nXaWthTY4lzD8+RIfF8dJ6fehzaI7ikHQHS4nQJG9hxnvYUmUsONU
sTPPHQVsjMWaztbrkA730sMWDUm/YSMYRyMsoecHXCiNFGvN9Yt7GA79nsRsf6zR
7Tq8fguuMf1w2xY1C5lVHlsiS4U+GRAy27v7BdTZvhAsuDo3EVHH4xPXQ6/DVZQF
OwMPFLQqlnfJacN5BHHS/Yh0+z5mMTHG3opqd6IloIM5K3202b0oPY/5KuvtEaFD
Z/Osw3GdcqxQZDHSSG4oozz3801O9Ff28ki1sNshjynOtKNJetTtCM62cV1+ElxQ
RYIyw4Z8/B90ft1o7IVnqEJ5ScbRJX5FnMVurbT3C4yq5SUBcEBQchE2RrNag7Rs
Rp7gmWOcYvTLutcpZnehgRUlpMKwFtlVAAvCm5TE+LOj0QJDfPaZNXquXcx7VjR1
/C6xGB2mwTBYwVrtdOu3I2iRL4c8Ruqby9eXc5UzvJ1pViJ+xrqVKX9USFYbtpGo
bkcff9wY+xmfsozFgGaJzFhd1OFxYexziaEoF/MJC6yLYt13svy6no1gA8IBWbLX
0KSrGdKIzqlt+8hG9BNbdfuAI/gNVDrxziGQzyH9z4SGwab95fQ3KoZVs0H13CWl
HodPv5MM7czIZmzP6uDQSMx/TCluPtvFNDX+nMSeEVfqeE9ncklJSXx1aFbdXHQn
xBAESgUCbSlEOqM6FPdLytcfL5wCIzwNiJyg+/jkaTHc9xlBRVHvDYNE64uwSRzF
ZMB/zVz1lVxpy0TFX4CwL78c4oFx1mJA5hYDpJp8s6zUkJCHd/yEQaqVnRkbvUBT
KG/5WQrny829+0ZuPYKpMj2H/j6mNH1SaIB1mCtoy3Uf91Qg38XsUGy2J7MQYa/X
6ApMXmmUE0/mT18oxnbtl2BcseuGwGaW6iOA7wYH27X/+boxS7+EnsZGUzo71NQu
Hz3CcRnT0GA15TRdFTdYo3Bz0pFkJPv2o8d0h7V0A5SkURjwJ/XKXzxFs4j7kCe+
qYq3RL4deQfulKDPXBJpZiR9wV3gJpoqHG+jv5vwY3Ly93Y3t1sISrfem6Rl5NEL
wEL6SYUXDHVODwKJNTl8Jwf7NN3yVzBzkLXL74bCUGniEKNBRnyRBK+lP99UKoDg
X6+2O80L7jORhmM+GRxAwPJ2zzPAkZZAP5KoH4m5q4gqqIQGeWr+AWd4Gspbcrl7
Tc/9GW2nin2tqp9u/ukTCuYwA+65cl7hulnuJrJEWgPGyRfa9kkFvP7A0Kgc6SV1
mvkERS4zfnM1W09zYxT4E6IIa+qhz4ce4ound2l06X6C9Jsp3VmMvbBAA+Att/DQ
oRVsu54DCfSIEyNjKEb7uoMmK8gnNFt3ELJ8UN6VrJyrkePPM3XIi0uj4+9frVZM
V+BCShXSr9gW23rlZSd3lpw5J8dHeDkcYYFqLHIVPJ0pFMXeZLQj9KQ3NAC+lsPa
ixGHNlBuvdSGgIr5TGLupM3VfkQViTvNfEYtbLPEnt1Y7Z6dgrN/lMJ61JzEPx2y
qsqx30gklIoxQsJd3EFXlkDLIo9+YfjUa2qrjOxblD7hONNDCku+Clkqu4ZP1Qba
Q40akG1cCxGlki1GZuh/CR0WvFG6GsXuOG37SeEz6kc4OTB1P9jFsfF/h4WD1+i+
oLHbhKZnM7yxXIoD1JaCfyEYmLfVhcHAM44B0nIlYWi7VpgiOGXpv1COHftKnbMK
jr2xqGlF0QlwyHS1J2ujbthwRNEQ8ORU59tuFLqYKvLPDHq963+qkdY6v4OJIFZH
fWO2UjzeMZu2v4nuLSYsy4VIf5eE1Loo9IApZrjeYnlvoyy5Bs0zIGSOe3kk429x
67URbcfws+2P2W8OIS3s0eSlyDiIrYkz2J/BCu+PzADkSTowEqTTy8AZdQ03luix
QjMgR2x4cWbcZeME3fcqFwGud45DpVZGS3oCsQvSO2fT8si68+mIHwIGQWgUSn4a
dW6yyqWt6mv4KvTzXuKm8KC2fF2zup9LVuL6043mbdt+WUZQ5wwIE7+thnw6D/eL
G8Fcy18Bx3fxuFE66+WdGq9Kl/OA0vdytvYHZD+ni0a8Gumsy7LhC0K8lQx8tyBZ
Zb3lvqtDiyVfDtCmScONF907vCBXcgw0w9g09OLVUG0aNMSIHelqD3tMvP5WpPYD
B0aKypU6/h3ok6RMLM/hjMN+VnkPMYN9lFVAlTkPaEpNmVoXyVCoFPbFMMtGkV1M
bTgWH9QwnYmLAeoKKO6K68HFyTU0hjAIUtDESfVnuvrfZBTyDCfp0pKdo/vPGMKR
jc/t3xMLP2D600KO4vgVt4BtFzcYUzC4O20v7nVRFaLfCTbWQQcizRsDM9dEA7Hx
O/ExzArEV+j0bwrEH9s725Y/CGkFmmbTMCFLItYsiLv1y4E5pcou7eu+IV8x1A6g
oh057F/0/iDs0U3DH7LpmWAW4BX1Ro+CGvPgeav3CyZRWZU+WIiuj6aha6+wDXkp
ZEvRozFiRRzMMtOCGZntUHx8b6T+KQILdhTGWp+Md70m5mS/sMyLCnZ5lk3oANnW
A2JnAcQ5odfjyoiqhc4ono11S+66thwEFwMyDDuNnmcP6IlapEfBh09u2rdALZPl
84veQlYP0deEnvJKJe2ZTxw8tAMlF4mAGYrtXTwGHvvEdj7xDlk/ZLKNaWqVDFdQ
1c33IJG4dT3MsckNxoWF7pKbmb46n1Gd3R5S8KkBN0EAv3EMFGMg0RwflfYkHFFX
Cjx73XOUXd3sycAe7CcCof8jkqoEVzmY3MLioLjF8rlnJqGJQfp93eLMF+Bgz18R
Lj9sphw/pzvIPjKfZ5nzVA4gDU//T1m8BldmMv/ZE0ghhfYDHHeUDIh8klqHwmlP
A24FSNz3+KNaIBuWi+nIVhN/7cPngUGvZf5i6kmVcZobXy+4wxXMtp1xxlwF1F3l
irEUalxw4rcrFbmouLMK2gckoPmewIaOjh+jlNweB2VKJq4II/nE804Mw6pg1rm/
UtFdKyDCpjFslpCqbE4bJWp6CMJqHt4bVQrmpyfmwTjC5aEeNaZ4SwOJI8RtlJy9
HZAWhvAEXva9IRtd17xEfRkjevKj+NXZTslZR1bZFTAucj5LofVDuMWeczNpFb5e
5AnFaBPHZ7fA+EbSamaFMW29KBlGDaU1NwmDAkaMmtZN5sMZhn5suzM8ja7cIEYq
LZSSS3KjCzS8PrRya/xVWs/VOuKcEL730maEWc2pI54p0sG9dKrSAnlOhxqIX5Un
SUSOhk7yqV34ztxe/yE/qIpR/kcylFyY5xbYXOGMG4x+2RN9YjDNn2wQl/8F2d4o
rKkkEaJBqfsPab4mqBSB7JYQ4Cu6zsHvLgbAzHeZ806cILGAH41ju2WwohZZizSO
4JOsZ0hykluX2WKKdp7HcR1aDfK/2YC8r5YvwYAGusXBMCZqdbRs+SnnCwMRy3kH
JMFN6+5WyyPhs3awfweBLAqCCf9OoC/aoMH6omqhJ2bCTchpyuqt7kR91EYAvwRO
k3xtAukMe/gyU/1bgrnMmyQXldaXQHL75jj+Zs/ZIDxA7VBJ0xvyGUkWQyQl2cw0
StL9/2MiTuksrZu4Bc0jKM7OPDFkonZnqaZUgNmR89WE8XC7SIopVP0i6iQZ1w4J
LH5BQMZv/IUqo1bp9LT5TVFu4vc7AWutMwAudJUAfZnwAxyWPNfuPCVy9sWM19vw
BZr0eHCtqyALkOpXCfNA/Gzou1EUAq00EmTsnl+1LHwgZ7LeHCptJEgEmhIT0D3a
koLxKpaKHZudH9HPzbQ4bSn4Y+B+8nBDPI0zPFciMG7Kj47fOv8RZ5JwnNzDGZOl
f9CiZxPYmcg6ES21FqPqbn/HglSU6sQWbqjq0kHG/WUKIDuqmF3yr1XwCFLMQ26O
HDBGWuxADLBLZPD/ebWD+LhxrPuXPMfIkWjPDwWvFOtfafhuwolgSQA5f6oVYsRx
LZ7K6b8e4RV7/ONUPk5gvqK8H1gz+3BBQOUxENu8l3fiFeEYzF3d4WPgqxZEg/YE
0JVmea7+dR6FtpLxBaeEsy03ldekfo7GhiimLcX8R8jFwbbiqfHR5Vwt5yIslIDY
C6cB1jz+38Ekdx7wOy/umPA6ajr7GUA8un0HGPbb3TtIEvxB3FS/RFV5Qbl1aEGj
iVzAu3RdccfdfB2WhlBi4CkRbisqxk/rWozJ3QliqGbgZV6Z5FWehxb6qudKpUsr
GROiIZ5lgMxsvJWJQjXHJKpVjH9Gd858htprSh+ZLRWngMsAr1OfadNMuZenBY8c
1wgw/e2dv+4uj5QFX3Pbi5bNGSYybkBlqqQlAsAMETskRMmHj6QAKOye++e1ckda
6mwOQ6WhNUf9i0pLe1NtsNdEbfNGU2pbE/NLE/jwMlqSJrnn7z/fuQBQ+Ycq3pKo
zXNgnU7GNMXaDi6INcZNlFPsIQyHfpzEuy6xfy0Hc/HvTAHw3LCIWuWd8BHd7Ap3
wBAq7o0vb9ebfJ3yvNL3bI4PFt9n+3WBW9B+gXHiEtfhuJkx55TNMB1koXU27ilb
HnU46nJrMMLFGPalKqSVsRDohhu0ufBHlI5KEXr/nWc64PPhRR3jbbyVMn0Pxw6i
nv+SnctRTDKi2HL4BvXcDBnaA7jopGmb46Dhu072QjgUBewrksqCn/4/BI5wARr2
l32dGcSisuejOC6ACS5qs7ckdB03Bf5Lnwfl9zVMoYSPFomqqgnDcGeUNTZ91lvC
6f9QYIzjBti/W17IDsb0uGMvDt/N+/ZsLESrEAdnXiSsinFsnqCMgr4bpJ5HU0Zh
6ZdRhZYTToqR+CNqIzmiCzjBJ3h7MRT+Vszm85YQ7o4uYaZc9xrrezIMzc5q4JnA
efSZKY0dPSbUyrcebwClvXZX7gNhka6jyvGLf2HKiH18RnIFUq2Mgtl87ZGlUfeK
qgZv9UjJQhj/bNFdlh625sxrur6JLgUdiuITh12XkticWSTcbryWfCPEkLKG8HbO
1whMfqFXE8rMgRLReb8KTlA4xuqgXCmxNGsS10E0qHgQ1kzBVJM+WwHMspAdkdSb
u/Njy1nrK2iEa737N52BrAc9lNNc6K2RRsup/2CHbNaHwD7/Co+2fi7j978wQACh
kj6wWxqiwbvdIKxNzwpwUMMWcjn6tgFOSM9+4hyDfE7qgbYugha2h0LSrhQ2NNri
yIj+P7eKoMhMojW2Ct5KAvG+6D9XtaMET5462uFbIUXBiqf9D36XKl8hQuzzDsvQ
n9GrNIJERnDfiCG35sft7n0vVHJiPUZ4G5RWcI7Q04CgXOiOoua+bxQi1pet657z
qiw2Sdo5YRbRajQSzg9mB8LslPB/MqKdN9icBJhUrBc4PpVlrQ/s5kAU92kwYyyi
0nmvEyRbRKhXNanhpZFjX/eyFdxCAMs7HN3W6mz5xIjXw0edHYwtq8Ngo3TwzoQn
iHRQD1xPCab9lFNpm3GGwAA2gaPfTrRCanN3l13PrDDvtQD7Vx5AfMOM6xq41zHS
GggI/gmNqLu71tD4BwhbvoLEvYEG/nuMWWQYIWux2Bi94A15D7fIm3u6XHle65Hw
FUM5w2KuJOb1lZrZ8dQeHguGVg0KBxQYh0x13W9Ix2FuJ4HpTHoioMx7tqodRjTZ
Kb4s3IUVZUpD7ney8AgoZSszjrv8TvjXUSNtifiOhNB+1nWU+hG5B1oXPIZap87d
ILYtfM8ruCZRiYejalB3a11STGF//MbitNj8cwke8UneyyH2RJJikUrgA9MCSmPJ
lF5vhErZmnafegPGcdzAS7ezw+8mjOya6NHAtLK54ruKU7liPpGtLBL/0FkR36py
3WcZWFo5nyjsdaw/DFVy5sihuC2ElaijaIxgP6f4YGPS1POgU5bxEmVnt/C9AIQG
EbnHEgrs2zih+P+bHe5v0XgzNvqgjzMcJFwc+NCGFDiaYrT72GxSOcA/w5ayO1dg
WRWBpSyDvDF9Kwn/gWEtcOj3BaPvwrN1Zy49jNQZPa3/RXwb07+63owrzgSYMhzW
scWYJzHjKzYl6w+0MKz51sNuQXjf2t0f5SaRX6+erT0/wJbpGWLYCYS36xQyUrkO
Ub5wjt0Ovk321MRegyvLhdtefPRfiY2b+8leBDca6Da2G+aXU79eN5kaYuZSpG7d
mpU4HQiocfS+uLb/vVU143P66v3gmwJ42Vm1Or3W9psLC+ADkFzbfyPsxxWh8oW/
U/rMc5dlj7iFI2bgRi6ukRMzar/R8vsGVJAi2/TU0WdDy7lUda9Fdk9Yn1bwrXJ7
2UZOVTh4qK4BOM/go0XLTlvJPHoTbNzjCuqna4nF29J+LrVcNAh3Le1djYyMws1K
L0/SuvWhY2E806/gW3Fpk41Al+TKJVbSvjsN4eg6oWmpi0IxQcJBJxnVajur4d9H
bqa7qdkmAilR3EZLYPdteU7nZ6qz0BzaiDUBahXvnPzUaRovJYwEise00sQkeGn6
pFEu1229PPveUNV0d1p2Tb2RpYDyuD9zkudXPq6Y7xvNZ8eaEgj2a4X+rxuyhoIw
4KAAXQ1G3chpu/05uG59OljWs4uprr+VA/TQL+2YQvVMhsZSxJAkRGEPjRXT3QUU
AX+6jhF+dj++s9UiNkNtcprNo4hxIMDAPLeXIr7Sca+GeCNxfMdo/AYM8E17B+zM
mbru/hb8ZYvdjX0YZI0n464QCadFyZVA7ZihpVwi6wGnAp0OXLNsD7GD2l/N5QdE
VBiYFkI4mnrmwbaLA5U9md6PAd4A6/afV1Cw95PwqJT9ZMQNsSoxtR8+sNTcTOSD
ZBpeRf6p8pdmntltx/WdEc3GfmKIiIXYvSb3Et0M9Pixnbfyzc1cx2pUNbtrqqlo
6YYGlyY4XLpv/a8EvuCB3ZqVMxpthuZkOntOdFrIyhoPrPxxQHujtKCqunclraMX
L0gi743teIJsF/aeFvkARVA00+UE6hj3etpDhhnTCrlE3HMq+DjuawidziU/7IIV
Z/Y5Lyy4dKMa1XRlcUOjMVsgKFhRJylWcP9NQRNVuO8lmPC8njtk5JnESNW7wFb7
PxcQzpsAj198ZJLBSUrhd+PXOmEZxN6L/MiS1YdTl6rk0+RN7thc3BycxGvojB9C
Nxy/5t4tkUM6wI/0Pbi6ImTBLq+0KKgzw/ZR7Y7F1bKW60KvPrvPjHeafd2JQDX6
iJ+IDpqLWBa+9kVcLlK3g0TQlNSZ8m6xqcnabk8+yq+VPruaThUxWZGHBZm5pfQe
kIPosLGe0Px61gttPwihmWw/84RFawR/ncACufwHb4vv+liUo8g7aNOswLdf465x
mO+6ujxwIxu95+J9OB8KE9CwYoy1xP5cZTc5WKf5tnssrT57VKChQhO6HWK6hL2V
UXtTI4zFe9Fehqgq+r9fGXlzHpdqwsHZe2v6DQOvwyxPYLH4NzixmsOVeEWAjE6O
3VWeabUhK+DNjSXaR06om6VDDKVLqqhASvxdee80V3EqwbR5y0UfhRo7FAkCFjOF
2m/4rfuOI/y32GVyai/uvAIMf6992CfMXmdJIn9VmvXmbtvRlzJiwzUnImpwAVWu
3HMt56JfydQylJVgU6SGTpQbmuNhImdKDJSvPXThh+vdADA9y1VepJPeK3PNwXn5
OT/I+86dGAaW7u9ys/0C3LIdLAxgc/3UNMXwnZ4e4yN2/DjXJaiZC3vJtmkLzVfq
mEzJ5orykyMhOkrm26e4ZfdgUyX4vDp6lcc/E6Rwbx9/ZGaKv00WDmogSMfXFgP7
nsr0vpZAI8fHfpaH7ZVkzlRkbxBgjKOgRGLioC4JaXoQhVHBhBH/1hXFYQ1PVInB
1pX/+m92K208fGE9uKUmtIBVd38z830AVHoom+QaRoV1e4zm3rEapyG63jpzd4pi
F8r1d/oqJqQZjIZMSv1oRTd9pomZIgEy7sVfu3vz2C+BBz3+ZTcAa8gX9lE/LHiv
soVxkHL1elggzyYpMHVvKI7wJvlT/erGTwxSXitYnY2Z4enVxcoYvp8DlNlta5ZM
VA4bofP8Y/jxSnB/wyK+fjJrTWlnVLBtjHnpV4Ay2nbpTlmcsfRb3VqNoUQR6q/T
/Ij8FbqlBy279X2airyKy6VZw/M/+OUWI9gFZNwsp8JbCld6cDAbY2JEtSBLZqsc
5i2NI82CxixGoj+ZkVLxd3p3jnZELyihs+t5eCvd9DOcAXJP6D25c5UDD18GqMTP
UBA6a2SJm75reEzuIOaFH2E9m1dGsdO2IQ7nJGrt2lq3VrDW6gd0IT6fhWLStQjM
W0aECXdKVLCp4Y24GAkIY+mCfSK2zfQ1+l60vlbatcMj63SozorKap5ov/B2HY/O
JP7xFqrPpimWKComcgoySQ5fPgwFKWTH5VuENqJGqG+nmPIswsfCGSfNi3s+/GtN
DeJ2am8Or2EYCJyMGgI1OptxdiEdDYD8AqBTFI0A/9vJ8j+maf+q2SWFeKkXaxV2
Q3xslethcQUkOyOA+MRtpeUOrelgWMRSHWjbVxWmO0+fZW8vSqFEsYHY8N6Obh6s
WasFTNJse9otbB4GrhzC7Qi51Gv5L+FnERWAtGez+4IgHjTe0RulU0XWH+KQ6vuu
uEBSAC1ingCCvMDTeMLHmL5snhCbWZqpVihjtmiZQMhlOKtNHIRnfr3tNTh68lQe
Ezchylw4Jp8eMQtVxEcHyBMYV8Hc2+9R/TS4Uicm2IZcHbxBJTiUn56VPBSlKKfp
304PNrmK5/EWVWWRTUVmuXzPPhn12Xivlv2jO++MYdeLjDNG+UAqcVPoDnWG6D5w
E3aFox9AF1JWHqhb4Phewst8AoiFl25QC7/DBGu9M1c3liWzpcg1pciW9Y9BmZ32
jjl5yWDtkVxhKveVlX7hqscZH7ygo7T7il/UAWGdsY0D5+2miHJAQSYZ9ir1IwqK
/ZD3FXLfsKy4QhgkhQJCbK10Sjbw8wwoOX4MzBUw4JEa74Q2uoO66uZQw5NvErfV
q1oxw2chPAi86BJ+oB+dffs8F7wJQSkWI4Ql1YQyFEqa5sf6xQ54+Ok4jOwGKuWq
rG5I3/UGqgm3hxY8Bxnv87X3CrHax5gKe6hnz5jy2avuMMR8Vp/SUlxzGiHKM5UV
v+rFL6LizIAmKdKWbUPflYz1fa01h2/tSZzsnayWgh4nqpuVoTQEilhhoQ5+iGPN
HM2UJ77NuamnDOaAkpIaLVEntsq4nvChe+Q9KdgiY1LKS/qnatoqMNLSJCaaqivJ
QWDzknkBpF/2KMu8q4z6sLjkWVMogVeBR2h3NQUeDwgIaJLqwnh2ORKl3Gv4phAL
4YGhS2oj+7GJQhlixERntS6AGv6O5uHjTYR8RANS5py+UPGVDCOgD7I7qYqIBlmf
6e+F0nRoJC6d04HCGiAoCpK0K7bM/K2jlkZZ9msCmQZRTdlTqgFtVX70g991Rtc2
USwKgDbDq0CX7vHclb2sHpsrUw1N/v+2SAZ8+nkpWuGhyEzm7kdnVXVpgByOIWXZ
M97zMoQDeUlEAnMn2rIWUSmhYAmaIor/IMWXJILI9TKaTBdG8EbKAgnjTcMuny7c
aFUTneY/FIJy5iUynTTMHbhHIdE+//nZ263Wxl2zdeVOf1J4g0yiYg9cK8TqVJyb
NeEQ/WZHEDYvOx7xNij+OYWCkaNbVAyktwDQxQ9jK0E7r4uhtNnlRt3zChApZnPX
HldZnt1yF38J+Ve1n3khSXYkbNlzkdZjIWqSt670JOkNPnALLLdwsM+066CuIPaF
P1NiUhHtJTLRyEbVA2iGe7T7Q5HGK2ic/Xoe3kNJGjYEazEPeqxNyDqnfTQvH1nq
9TZ0+z7j7XWfdzuUwu+KgTnLxuXDVrO0x/GcXEgrCHjFH1L91zFFtz08LJ9cz+ks
OvZ3R8nWV7GFgBmiI8ZeIp9FFeBQqlKeWIm4yJgaxmHP2FZHJpyXoiagwhk+A1we
qlxo1LuT/olRKtde9rGXCiEy1t39hClDx1FuvKH3Vj7DQhqJPiNJR9wDpyQ+YE48
Ow8TbcIMkw2juxv0jwDv/QAkgESleAyLpbj4/gqpyXeGlzspuwgAq8YwBscZ+Na+
XO6AtKYWcu/hOkLy2MqF8irMhZuYZXQjyLUaCS/HnpxPpPLxGzi1BLQcrjXvNdGk
QdzV/tRNFclZCLRH+wb0dd97fYn1UlydKfPrEur72URjkSIZ5H7P2Qvz3+dd14cw
1fQW7SGqO7XxXJ0ihK1JqkXXayjXr78kKKJjcHqh8EEuDrPcS5PuL6x/s0pwmas8
f2Yc7gsQ2rCK69h0oAeIm850hf3/gZQOYFP0LoiZVMHUcnVkhtJRHFuCN6TFeCIR
e9CaJs/mmd6mh3BiCd0RmptZO7SCRbBpq8Esxc/mWyXKW1midydYanmc2dxScHCR
z12eD6x31gr+9vY+2QYeYdbfL1dP4gII70XS6zIGhkOGlrc77NStSjipxZbnQfO+
7THhGoTeX+LA8cVHPDtJ5CxIcuNXeJoUEE71JYKsVY8xviLJXbU4BS5wHgNc/WDt
eywetZomKVOLwKJh8L5TlRsZJ9tRdmD2swr1QnX8vpo/el+SdvPrnxTHfuFDTy1N
km0Fy4rP10PuWMRcvzfdT9DG/a7XLhnfyvGlaFSROsOYIg4CbijJdTj0s4ct/J0R
jcAIby9palYzp/EagOxB7hkcPwm3W/QkppLpJ6/BxyZe9pN2h/FGUh4PJ+lRG8h5
6cnQ7dFhr7FhBcGfPStuZ5Xfhga+8k96wlCvGpdXlD6iUcdJesDL7G+JfPiQgUru
XFUfxUPRP4qPJF6cqFtx2INqbD2PRRBgcBmCFYc/SrHLOrrUl0P/Id99o87KGpHc
EQAyJKXkBltAPfua/ISBoELHUPBCBFZp8HnY/TTEM8x4W4p6A45zAmL+Zk/fBXoi
0mnKP24sUFPFGYOiAP0KY8T/eXxF59/ttjuPeYG6rAx7qUuPS7vuBZ2/Ek2MZjb5
L7b5CW0M5eEP0qEJuRYKaI8gjGr80BqxkygiWfhGGAPc1eVs37lWu5UHW23ucMQm
A+aTBt8wfzKPO8VXqG3iz1IQlwU17pkvpYFEdtG2KLvMzK92u/patUI/WNQppfsz
Y0G04/apm2CP+iaQVxbeWcdoz7CFGeyI9wytz1cu1oGtwFhrfJBPEDzsArt8cNit
ZXN/XRL0zYkWX3oOjB+kxn6s45849sgFtY5nuFKptDjYcktROljs8vNS1zGTIsMX
ngm/Op+Oe9vrBxwj6Lk+pefpoMXP/GBtDa7bApaYr0nJiJZeShakfBFUy4kH4Kd7
Ai4BhctxQ9saV+apScu12jV7fpgq4vOTrB4zzmrnxPXhJuhIccu6J0tQ4rgXpULO
yGnlTcB4j+9YHZND5KugASWrUaV6OFOCzwxY0VpW+j5p8iU7TEMxHdD3glPhgP4L
q0Zvr4ie2b/UOTCO1L9mforXt8gv+RN95aWgprnSiqqXnGu4kzH4m13Fdt1PpORH
n0euXOFDR0G8HoO3e52dOHoa22IpViG/f05UZkHEXY/zjn96vo0+MQrDGmvt9HoM
RuFkOe6aQB+p2zN9jx4VvMfthZ0cei6z9wB+RhpdyJGj7hX0DlNnYEQvOOvBiDDg
75jLUL6RgfodKxGRMACi9s0PYKV0pbTfQX5fk4lkYBCvR+VtQj9FlCNmXjFgHOVl
YL1FNAu6yI5KpGj4zDmFsIrJNx+W69Dzv5DPQzvkj6zl7adDDOeXJ+/SnUr6gnnk
yST811sDd/AR+4dD0kAOPOGWL1ELUJt3nuzUEeV9QgloaX5ex63tokg+/7JWJ9/O
ZTeWaGF/jdYjTC4tkgu8R0ce3EKA1nVfHOyyqOA09bncyBBZ+0R8/SCgyVDLJ2M1
37TxxZX0Cdh8XkVo7cwPyrQFPrBVGzrfCBHnguHbHGI2OozKX5mdOxS9Eh4OCnel
KrmvSH5aM1wFGdPFLy3bf+hVqL4zzyPuSyiJVdN3NQnA339clnVJ9cf9Vnf41sEW
xk650NkvggIdwLt80U7s7xuFlVUUPKhi0l1LfreZ/E630I3pKkd52fzckSTLeMEH
OZHVo04el35CBXKowul5nv+T66J4xPn+pT7Q7Dn6+avIuQ47WcM2JKSkvQyfU8qP
nUV1yKWOMWokOnO+fLXuq+NqNM8FEIIfra6t9JAw84D2LF7a3iU9DHesNNaM+j0j
jIiOYn5lLpFXz9/9MLOydMLKYGd7RgNJ2YGGomwToYHKCQCuqQqqEFZGbJsjiNpJ
KmL/SnN1q+Nh6tVKgN0BEbDOPzKtoDBdnKzAqYwZAlw4YMNiNpvLsec+6Z1zbL2w
m3kx1f/xbugceu2VIQI80CTzHSzW+NiGeMwjgVxGQ7dwynW337z1PsAKCmnDnogq
FA6Lscn0vlx6CttL5LaCQsCI0fR/NwwbxHtCYwo+eJP7VG/XDvUQ3OZhylJzYmhl
P3zGDc6elDHCP9LAmkhU09+k9WL4xNQT21xQwbyyBQgzGsZ9aA2Sd1ilz7eZHDT4
oRndsVnL6jWuCLGhGYwXB17cMHr/gTWNL5wKl7I8P2HRyJ/qw73U0loTTC9nJKu/
d9vfKCj8UDxs1caZJ9Uo2LA+NXN8RPPRDQwV3SCoKoaem/PXNQ2WiSmQpmGOTQmj
JSIvukCuqYNUqLMZAdBQeaMKzmbh3uaw++OFzlcV+YD0FHC76RhL6XsnzeUi0e65
zCHbqmKBYA1AjXlApSlcb1+o/WdQDTD5kBaWB3us04H2s91AuhQ9z3EdJkERwcYr
yi71u8wD3ptUs4r4O/5lpbMq+VSJkPsmKsy1pTsPIlr34a6s4PVH+7G6a2e+CdjT
FC176KF0BXAwjCFNdJAnu741KASUXE3W4vK8hWmoo3AbxCJgkpqyWm85jZr4f7eF
yUQVzuTYbFT8vDDp4oa28mZBPAAZHDF049LvByQo2vuhILS0hQN9OZ4tWiuOsdCk
ffdrLoGtn6xMrrp+adC2N2Iw7c8nWrqtGBaEGomp3HhztqsaBrPxh92HujbIPJ9B
9st9QQocMgtBxiSepOEn1T8BQReRAPUDIcizsCRrQQOmD5+/vyr6tXNHBkJAnmo7
8eX7qwW2OvkjI39M3btDYKm47L1FZz+dci5DtswPdd6DM/iAPTnKBLZzKMLl0vib
TNrbajQPrnXgyKfmWIO5QeD8dgoZtmVKzdCyl42C5FRAoN+L16laMuIH0Z5CEECT
5Emx+om3NjfN0XReFWMwbq9+656x8P+a8gYrx0X3YWwZpkmLufT/ZlaRi/oML2C0
N8NaB4bV4NlWOeEu6hvNudzyfpMbmnqI4KlgutgRSOwQcJv4N6MaL6qJhvG2HC+D
QqIPHUwI8Zw6QkCjKaoUr8nBP7TQ0PMdZUvUq5EWr5PIocFdUE7RCPJrKnEtVr/c
LhmViKQ05QiUsJ2qnQcfA2HJMuIU1tMkH3CUe4cwbtRz0j3Ps3eygGXdm2gsHjGm
cjxjyesr63Ux4eAqbxTqMg364KyREwlNPDBqVsXS8Wl+F33znW1rk1+rrTjdZt8o
SDmj0UcnxuN8MNnjJdmFLarb2LtyfBJ5icSPM7Oubumhb7q+qpBmj985GbI3L1g5
JEORpo84hp9z1NZqlUFq0KlXC7VyMpUFwgbeEYNc/FolOYjHnvvw156dSgzzOEQY
cbrNnLuqzlLxIolitC422LHVoloRmy61Fv3oV6D+n7zFaDMWHgS6KpeDfLyPziLJ
omyv4MWrFMOGFoiJwYoEnxczgiVlGcUOJuomiq/1ZiQUtet8nu8myKCcAWZZi9r1
aRDC77rW1M4irzztCfPke4gH8ibi3womXG4D58OC86pwB2oSJ8qSgavhlh9NE2JJ
8v52K1h7Yt/7cy6970mAiD5FJpeoIyC06rG6PntgYHcgIJ1Zbc2gzacCi6wFifDI
zKfpuNRs0JeDGsCHHyNObwjLRHzk8YD9iZM/oCFC3AuM3lbqNld/vXwA3xMVWPsf
afYY7moDeTjg0b4Swg+ugVviI04RfpdWKzKi+g3V4A+WBgnx17Dws85XjT+xs0yY
Gr03ATgz07FCIRXTj2NhNM5YtqWpUasTSCYOFVOtXhihb7wT1j7J+6nqqk9KlCyN
gM1ebj2CzNV+Kd1rOVTa5nLMPCgsM1ym+aYaL5qGwMF1gxYC7kVs32yP3BLrJZMR
bUquk1sXkG5LAwAozyJbyiP4UoNwUgnfmWmCClJV/cduQlDABmb4IUATKP8c9GU5
CuH20bwq6pa+ElUOpGWxlUyWMbqnvYrySxHdpFJnBiE0wpKL3091QhZUd/eRBGq5
lq9MOj9a1MUUTiD7+g3q4fKtqkxXp9c8xtJexDQyO1Lk2EnrOSWx7cZ9xHXXHl5n
gKM3V7MHRq56k4AxtuVXOR7fmH2UEeJMOo9Tatqktw9f9/ZPstSb7t1OLtA2Gpln
L/oUsO9tkm4l6t0yXRWxFGMP3FlItPUMQeW+qkbTH9/00n7g/GKJoO+ZQQQuV3oc
pitxpoT6slYiUsbe0SKoe8tGy1FbsUxWAjqJZu58ZGfyHtuzBZotxy0syvXxIfYx
1QjETIPRbnNc5T1ytEPLHmSJ1aRY7PFTC3QG/O6qG0eecjJGREhdaJkHcLL8qNF4
rqQta6oS3/w86nzJHaLKsyPsHxSoysI7gO64PwZ8DXajM82C9tNFU7/NyLPRRTBs
+9YWAy/cZ2t3qOgz1UjU/JFnL4B0Pz384JrxVuI86KzgXwq5sLNnINXaANfaO0Bs
GVW9C1HuNaMFBVGHeIqSlSLi1AtOkqclcniHh5b64TpI0UfnsfMDXV1ZHqHQ7WoR
vNyP6RVD8VL3KhOMVgzWyuPPHiNoODDoJFM5LI8hYc5w+Q6ew/2sBD9Fuo953QQ3
UojPSdExcxsTFIDCF/SA0MRGsTGWasT+SnXp/0T9SJzpzpGo5Z8uXTf/c2q4/h6z
0BDIhhpk1jy5BQ4H1dvaVnRTs8Mf4Umx4PoUar5ycHd+R9TapfHgDVeD2lgBjHDu
vv+GYcASzDSBRKwNAHKNSxwpTYub64e6W72LP/AKdKgLDxDtsUuW21Fg5nkYivVv
kW+CDBO5PQxy4rmU5IhcNRv0r+YYYx4lFc+gZgAQukMJ8Oebyi5izL20dMbOIitB
fJsWVrujj+aBLyugTsOOthYMEdPfI/+qF3j4MuF1ePCtDBjuz4smg5hDIfyUmBHL
OUGv2oYrtbDoR/1UlmrM9VpXGijf5zXzBjkykfgfKuu/512ov47TIADKyfiXj7gh
lyDeZNmiN6wAArXLV56MsBqDinLOcuToFVGNWkQsCsFgq+XWtW3TzrM4jGLTXNQn
KkN/AimvNYN2REDmDBYwxEBcpv5mPxpBtklmyzZqtDsUiXUWUalL46di9a/qSgCM
idxjj5uTDOKY8K0LCdZwm8n11Mar0XWxuHeSLDNOpsSPNfoaMAjwPV3zNDFNu+K1
4lU9wjopPw169Ho0MuPDxE1J19BVxQnfC7+4crofDcVmnTNxzEezuGkHpSUFTgfN
g1ppcxH0Ni6kbjzKCBcBykjqOxf4cuA6dL5lQfrthF3pHJl5uzbQAd2qq0WKuVVQ
BoSNNX44kgwx/b2CxqXAed0jA9XWYP/P6MjPjz4ruMA/SQrypREfBqQXfWVwqQzA
MNyA9rDJ5tkr07qoL9hK81CzGdPu6mCdamWGjmmuhfz6Lbl9aT7vQi2yF/tprck9
z7+6QSP23UhbIdVAinC9SIxF+oHc7VP+ygZWf1K+YaVX0Ni9hsDrCEIZuJQOTOpJ
wOZN0SHNd/7nn0ZyvdrqVJgPL1n2OGD88g4J/fsR6kAokKedJqOcwI9ivq3Bu7bY
Z/BHcaqQqc8MaswHT5v+qM3ef2gnLCJMID8VK1I6fo6EpizXqZuqkGGVAoTFs/9B
jSfk+HiUm0ncv3wlIITuvNNFKKdB/N+uwLqCJQ27jD1OAJMsYKcX6cT4z6VEVFBQ
6CVOgN1IymyJ6FeTFRAjevdzEGKYNv+PjLoZ18AvAnPCo+JqQSs6sYBlJw1o5pfJ
8cVfeKZ2JUhVJ0Ek8Ih0hzeBV9+T6nm3nrlbxLnvzGrcobkbiuz4wNCpL/vLzZgY
qdbziMhnf/FH+mK+F2bMTGQ/0Uw7VgYn5fd4hDFwRJS4W4vUZVQLPzW4gtofAmtx
06aJyFzzfO/6LIMYFc0iBDZqPcl88YYlcnZrzd79nIHNynJJQJbEQvOK3w/cX6se
ebYPsCZqrs/7JaGG7d55xp0Tz+rlnCPwIwY6pLMx2ojOJ8QBVN32VAECxVK6d0Zj
cqXjlqAxSQSVtYsOLsmmBsjf7FDQkbUbfARLGcB9OEsD0SPWE+tawC06WjTaYvgw
Inj/+DCSDJ9nFwdbucrZvNs9rNDuYptFcK4EmsuSb26ob68nF2X1aqSs0jQpSEmf
+0bkEK/o6KRoC3ecWdDJP171HOzwuGk+i0Uv0W4qrmK0i8wMa09ZrzZ0rkvnGPKK
T3+uwBOfc5fy34OU6yuKjaHKyeNjjuNJ2g5+IODQw7a7HCpw9pkhc/k4AgrZx9ba
IHi0nlteKp0NNneoqZUb44S6A+QbYPmnlMtAZl8z4BzpRS40QieS9A3501g8i7JY
vfy7+SsPFG5Y8f2XlLrXN+ZEda5a+PIp102YpnPCt6BLhdKuh1ZdSSR/VYxfw8ok
7tu1RH9BmZo3VSlTEN9F2w/yiSbXIlyrE+F4r+2iaEKmrHFBOsVli+rA7lfbnnRq
3uHpitEibWJ2IuVc/jAPICh7I6Zdc3ZICcDacHfGRdfLdTB4l/8HiaHk8ZgzVYQ1
cH5dZ+Wct7xy+4iTU3TOKMcRMo1zWfkqlGlopzfCKe9J4xk5qv/JZFyJ0JQm2Gc5
mnHy5OdJqyym5qQOssy+dFIPaTYheI9IGolaaTRsxEx5sqP//5vjUMrllRcC40cq
6LFnvDQzGriGsP9drinUj/MR0JjS54cOotdKjmUioZdUxamD2VwzqpZCOx8Z8HQb
kyDT+Sfo7mlJoDouOjoJm99oxNqpHeW5E/jYa3xjIpxB87RMbLGhe66eUnLXy9cW
o3YcyrJKmz5Ql5/4//dosOzJtdtiBdFm05gDzXHfsOrSRpOs8BZVsfURM+DWqjJZ
P2TTMZ2RZ+vSRbGmNVikK6+Whh6iATpJU6VJM768P6Y3dea2mnUkXCesgg3/mBHT
GY0R1vKEe3H7sYYGbj3WnZZRza912cXguElEpkfvhGafKGR0bG/DHkafSqOnovcq
ogozbUh86jGTIXQbb9G9SLAybwbqI4xLb5l3qboWxc1qJ2rIO4B0ivTZQdKF2iSA
UBODxJKV+qYvMwDA5eSRNRt1Hr1APnQZyfSiRu1HzpDZEtskjtS/xkcAL0yiTZjx
zQLgV5GI0lnoBnq91gCrgY0Suks59L0Wc/YETHkwkP7BL4qvPyXJc7YUmCftiGLj
Mui2FTT4MhCpbyLOy0rcPeQ7qjSwu9MjzHnVsU0PUqHvlP/H6PLnXW3uZJy2cGGU
y2emMgzBMI+fSWZq2Jrqbjesf2usW/8MDvedrX/XptZCy8QZn2nh+0dhdKH/Amwj
BTqLrQwZ7gV6GphrpwvZtSQbyMZAp0kj4mPDwaWrt6Aa7u38tRiQL38dFOqlyxb1
kNPMjfm3WcDHgLwKaxXq4lzlKjxMz372uLkqND8VsH0UFhuDRVR2C2lQnazUwKpM
U1cQNl0IAY93WCM7rmzR8O9loRfVx9GLhKaWb8NewkJkmBd5iqAluBM5a49t2nX/
xVlyMIr3wIWSvm/nJlQk5Wjt3bk3O6Qx+hSDEE/hMlfeZnT0jPUCvMPREcHU/+Y8
BEv1K/cauYi1rBsLwPJ+SQxsLELztb0zYKz8pOg+Z+8TBfhirSWKqNge1Ca/fxvZ
3jS/dh2GFn8ts+TgMU6oykk3zGUb3Co+1wCn/X2QfebmbALxN89YPM79wGzEZjHC
Jn4ZRo7XKyUV/nGfYmRgG+tai24/DYhjkVjLlq9djv6EVHfvc4l/4wfHqX/lpexE
9/uZM4AwPdLpbvjGxdy8XK/pOLBPml+iocJ9kEIc5z80yUipa6BKRQBUxry2qyea
uKt1BKnv2BlYt60MZcA2LgawSLRMGBznDSqbzyDkcRIGyo5rHTWg1IpumLolQzo2
+z4O5+avlkrZn+nKiORHFqve3iMbpnmXz8nA5k9fcfLjYQB6AwFmD43H0Z4DSBOW
Bnq/69aidDLyIsQDEkyh8qipPcf21dPaNEPiYvD1OK0P7RvjeupCAUTWsLxrhDJt
7kW0PR8VW1AnTZDD2oAWeudH+8taQ4NL564KHucc5BmWmik/KvA7d0psl7TezD3j
TiMMtD1ZTUVq0GZ3ed8xFvC9l9S7+4E16fysg4X2Zei6lX1dHazvVYMpCR7gKar7
qm023ukwRpqAmha3/ZqTqVszRKBR2XGL/px806YRpNV/fpo+Yyh/mR4HcktPf1mc
/RJSPPIbBz7zr+8BB0y75sNUX+sji2LCK2f1uG/5kSrDF0mJQj1nBVX55jYDbwZr
JTmzbM151hQz8vN8vbkxFDYYGzwheKelFJLgmvVO9QwrQKIYI5V93e2M74HYmRpp
uFeag243gF1v5d/PdcaAzGmspLfQR9vaahepkUNTkSX0ezCdpgCaD1XSsOTp1djX
Voy2hqJof1h1x/kAWaouXcXYgwmSDxVzGley/GiDpkupqxjA3GUghyoej738KCJs
LlA5fb8w/M5bK6gHg4VqIj67bi6W0w24GVJCdVoCs/u5QsTL1LD11AYQQKY3CcLp
lWJZ5chlT7miXla7wE0NeB2MZQi2/2cVxvshe+LO6cWaPRABipWoN5Fs2tQxWovv
MXmZPGDWtLNQHbB8+A/GxHjFyDro/l+1BYhtsWB3ekTfmIaiks6uKOLmEZwN+rrV
TkespF/9Da3Z3SGxuWnLLCSDZWK5BplpnSslNdRQDHvCJhoMQpN6sC3o04LMNT2q
W/TTZbccSegxNTtpouNMNrnHtf8L2jYFBp0rZ5dzwTUZP7HaV+FrrV07uoGdsKQv
6AhihPW5nF/IFe0YsXCgD2abk/ArIYBPC2eNmNr0XDCxKn9Sn4Tpu+HM5GLf8e9k
Ep1LKaRNs6srbVj4VhLG0AfuLBnbWtwWnvd+LtldhG3+SOI1xKfCYem0g14CGYd3
507anS73oei34maa8N3otJMRTjg4fSPvBiT6I9GSoH75LKyiyz4QqJL6mqLsSBGz
n2YDY5uarHseOovJiAWzIxXf4d51pjFK2nZnDfieY2QFrWc7yFYiVuB4qqR5salJ
zo/O1j7gAT2hdGfL/U6vN86ZDdMqAXQsn9Il37tYkDAFh8KMdxOmL/sNAhYta3YM
JhO7p8bFwzdjMNOqMOuDX3igvesWwax4vmQPrea/xhA9evrzXxMNSwI8Wg5WKUTh
7oALXL/zkuIW4zbj3t4GUi1mc9Jt5ASOAJ/XRcOXseUMHcZgty4qDIhvH+7NBmsK
hhIu/rdpSFgPulixuymvQkBgBGqg6ATDTAaNm1cky3lyq2fW1Oh4iKg9GC+eCEk+
bMgkbasgX1bzmXp5GyrW+MTUrnM3afDAahgwK6QvZmSR/qATKcnybYrn1vmtzdkZ
V7JeYtochU81SDx4MsJJG7GEzcm0a0JhwoKVY6Nlxfa805Dbsj76YgmTrFm4ITrW
NUFcShZ/rj9p9C4aAEusq0yyfMen8A2kvukhsVp5T+SXL7LmsL7implQlHrKuX3I
MY9SA0Fj1Zbcssxj1Mv7Yn6y74xCScgWW8vVHf0rUQ5kAMwbYfYj7OYU0xOtOBLz
1xcIKV48e3P/Sebjd3wOR/LeDf8jsCwiZDFkbrCiDrWFt2hk0M/jGkQPADK4AlMl
imTj1cdRuBwa2jwAu4V1qxYHB4bPpfXJ9uOvH8y5iGM2x1ByX2UGcLLBvYOHZ+ul
gam4/TpS0jdhCpKSSW6AxPEY6m6udcQQpI4x7VycRsd4PlLB05kmK6/kqRAo4QnH
iLYTe2qqL1TJRXRRLlr2EHPAPJJTA6b2cTlMtBMlUr/x/GD7NrNvqd5DFlatsb9d
4xVpNgK/FsIhzOFP6u/94G9dhJpPEbcNb3FgpM/rTZyg/8gZA9INIGw9/5IjTsRT
Oq6nXYrR1VKw+X/Q/5sByzRMACQGl1l9oq7uf0QScQH+V/NBuYhoMj0XR8NGbjQM
fGJY7EJluIdgdo1vXz8j5CNJ5ND3OHLRw6+w4wu6cH+QmIyOsisIsSyNnTyRDrZt
WqsO2FM5HVBfbqUeNtEP3IIHKLw66vfvjPfDBEaRA2omhQpJy2sEVpzZvPlKQzOX
X9T72ZXNslVHl1qVWx2/NH76zidWt6kQ05myyIvE94G3eEDpk9274v0hfF92D98b
WGCj2NcoFYY/hmTzNPCDs2LLuzPCWTGyweGmh1qFTR5hbFzP7SViQLyo+fMSPfXH
CXzuCqoTgvBvoO6QYQIvfN4eLV++ZsbTLC1k3PvA2No1lA1KipUDnQWI8qHoarVa
zJu+P2XObimlmQQAWFgjK2JxKfKBaT21soDCjjcT+aNHTwMjGcg9aTtoZXBlRt5L
kTFP8Y7Q2W1rbe8qZKFHN9iN/VzHwmwcE6lAc4j6IHuzFjdNsVMsAWIg0Ca2aEci
jH8MS/OQCD3ohelMWaLSSmWk+jjkQ63RoDPJRBZ7bpKmqb1kqvv9aIYsSRGXhEa8
VWK9f/HdBbCYHV8QqFm7yUFjzsvTTY/Sa/H1NXuHbN2ZgFCY6dP4NPdwDAKfEiGP
pK4s8z/2eib9twWoRS1EO+TP8V3CDm10S6d8j6lK2caMUJwK1nyzydrm3WPLXabQ
2UE32uuaDX06aV+MZPSdjjFvwDr/FcqonG1rSVbPeCDri9R4qjU7dj040euApBpb
rnfetDJ3CBKtqw4i686AQ22Pf/uMsyo7nlIttulfhAS9lqLIKzTjlegPcsAML5+Y
eurClMFKpdrJuY5ROO3Necl1JtdOTEl+m5aUIcA4gKIO8pj7dRWsMSBDtOhYq38b
ajTCEg+QqAzUxktjGWAD5QeV5msrE3w83YDWEKyUBVD4wr2RezuF8hGrjEzZTamP
EYgFy0I73nTOpjCe2l9G1t2PYFGujO59+zJX7MXZFc1LVWA61sNSEDB25wCV9/o8
2ayTb7kt+5zkkKBcGbh8men00rqkoa/JWLu99KCFvWDAnPUDbimhc6ybgU2C0QMG
7jJtEgKsVlR9F1EnZtgneMKtz0yuJnKVzIawsi2J3njgUg5JNaYqjoZULUTnXlyX
cujW//xyFNZSN7eg0LpgW2dN3Hp5FJFX1YOFdFZet8GGE/KDdZ41PeyModUGbYHI
Ao6Bb8jZLflPOSEDac/7td/yjwcWG7BPAGyzrdP4Ybya5UlG1SnBqra2z46sy3Lt
E3v9LhtTFBieTiviTl5Zb78ySEviyYm5kYoslm2dTerQjsIienchvKA7LzapcQeD
CP3nnjzCMAT/TXQ48eU68hDoLn9buNTM0kvDJlVCa0qMbMhHrz2p8wMO1B8eahZT
FXHRIgMXEZNk91zET+Y5Sy7FaFoItpiRSObpWzOSowXpvknQqhNu4r9BNyWOeXDX
LeTQOu4o8c3DbJBILwzB6Lc+YAxz/oB0isUVmTBhQ4Ar5QNGd7Hw20yPDOGt4S84
PL+BMaWszP9SqmK3PBiKbG08zz1PcDBGZSyXYt5O1algse8Jexo+bRlmf1SwDFV3
VAKEpO9PaIDYIr+jl7bv3UH9RicU9/6bzwAQtzDgV+mIqQv1rFx1+uKXs6kQo+gV
EPC8YxdfM8qAkEyOQBOJ9Mng5iMfF8cJXVFBe/vKzLxQ0eHVTlTrraxYKj9g8uQ3
zgHzz4DP5MXrLEbxYynE23djeeRSWVds5PAJIyIVZBv6FcnJ/8JYBxJutemOkWzT
IsIdEJktNHh3/Ddtc4ftzWNGVdvhOYJj+uiJjJcqtRQKAoX4ibI0tkPfUwtGNbhz
Im/agHJy1I8xzOe0L0T+QVQ59HE94YBHaNXXS1TDUktQV9ZxxMNexMzRpnx9JdFg
r1xMFuSnTM8mh9TMdSLFbDX2iqoMFKrjC+L5bXAb/KHeKWpn8QUsuhAfXJ/Nlr7u
qMsakQ1bncIyNNncRVNo6ulcBr837J6qMsFzWndAB7r0T3sxWiqc/nqJEjIMOk/i
YvjzfYj1OLozALoCqAj+r8DgxIDYj2TJmAYef4ESuULyV8e28U3Sskf0uF6Rqytz
qYrQPXVz4uNiWrxyyyNYno6d73ZXPvyH2G0QMAK4heMZoenpN8g2+G1h1y+2l+TM
1/RU6gxPIyKQpcIjxPFxP38hp9c7KD1MCmWbUneirn3qMyF7RVkwok1Ygys6SgBk
pd0VKgwDx80mWDIXSYoFMAMRkGJXKWl7WNC7id9LC9m8bCeIxIQI4m4YblRsM/Zf
FhQv/qrdDNWER+Bqs5BAOUzg79R3XoRGcpcXqJ5nw8S6L11PS+6ivtQ20yeltJ4+
3J2/g7Qr8D8dF7iLg7MnxjvgefWPUnUiWRZ/d11+YWvfHduOjtoPUvvOjn/EaXJR
dKXjZg5NKW3WnFN+D1qmm2gpUFgSrYy15lWFKcwQDYFcQrIyk960qFUuNUL8XQdM
LyW5j+Doh9y0eatAijM5tYUwp3aDnPeu0/dooLepeSy4+9uAXc0nz22lugFpXerb
tBOuSk7BSEFYUF85p48VRhExXS+cfaWPHiyQae5sdIMpd8GZkyUeuPxbWnKBvz07
6DaP/jDEWPE2FfEO/HJXEz9Dy8cfevpcqsrx4I3yc66SH9P5LOBWKVFgn3oguSPQ
LGWn2ytZsJB+8SjM9tuJcWLRuyA5ATW5kgH1GuqFEcgPlyEWJZmBJ0zbdklp4nV7
a4hK/FgKluMdA5+1eoBpaP+Jzsi62Jpne2g9A8v8XsC3A3SEwiqX+bvUNO5hNqgd
IU2isY1HPsl6JjUHAJIYqFG3Bfn1a20CWbrVy2dijwBsDs9HBlTddYws3lA+saES
rcJHdCZtMvvK+XLiYHMQJUfNnYgLxxdi5zc29EWSjddfQGrsxXScw2JaOjVGO1IO
8kpSuINYrjm+w0D0ZvkuhwD8mvv6UCJF5MaySfs9RsscqUSvNqZ77sqYfA3GzNX8
m3gAXt/rCHFbktwHo5BnZ5PkpvGSxrmGXBSXwUZlRJWuDIM6sBYaond1h/HPxyXi
KRhZ+3zgwQAOBWs88oT6PDJuhzb1EQsWKn9Ct2vMBKpN0vReykQ6Tu3sOhEMaEqw
Z3Vg4AdwdmsOlnZqJSvGY+QUVcW827zeUf+705sJcoA/5lCfGCL7dn+F7HBi8eIs
w+PD9BOiD5XvSDX83CeI4OMdaqCYrXnGfGjhwS3USaQD6YwkJS0p7o52ZRX716C+
rmvrydypiJRVu+OQG21JRHiQG3ICyjy0XZyT7+XBmZ6Wx9gOSwncSFXiSobytDUX
aAN6z7aS4b+n8FTpQXgPQOKI8n0w0XOCO4KWIXPLg/+puauCua3kyRa+FSItmjQU
MCkYlRiIqlS6Fu1tVuwHFPP+oK+TKoBvvO7IHoVkcRuf4vWKAOevuM2f/oVglgZf
88NCG4ecHRiELNX3gSpHN13JqMGFnuigbJvBBFvVRhcU7kav7l+YD8KGKr/wgEkj
7c9+zSEDBv9HlyAUE+zzgsn8fcSEpUc3353Lkrq1VBQSZS+OHxQLdFkos4HvSsIU
pdEt4V/CFysU3BviAm8fSKkSFsXMs5sTWt6aMOy7BnwsuukGQuORxtaYdAQjbrJo
6p3ixFbipjeVJTWHmnVlCPL3kUeQIxWqd1ei3b2D2DADedO1htsBOrJEPW5gDqzP
qrc+3BI5kF5zEg9fOIh0M90SrLW/QQTHdRzf6cafIffrIQOxOodC8HC4sqfcKLaP
f3OCu0m5yPB+qynQujB/l3102NTxRxhvjkLVM0+gJJ9HpQhAPIDiKWHfYKqkpaUt
3K6uII1tErC7QxR5ba5tfEbY12EzhWYhzsglTqQYDWnIcUk3o8vJBGZJ5kcMkHVz
d5piHFQlt4QEnKc+UecHxtcS2wP/0uXaC36KtC8zolfI/ddeP3BT1d8rYTXBBhKJ
qGsv3pDvhmyITl2tS8ECo0uspzyrCRNg2EayKs/l8FG43dsoF65+U3EwzDJDSj7n
ukTqbfXWQ6O3CoK6pH9nAAD4zoBdHgV+ByS9ySo0fbqAqQaX61wKH9Ceyg9jhbus
ltBcC9ag06ar9+A65QINGjH8yrlrVZMRfqEjJLFbBZrW1BqQbA1P7fV49dFZRD7y
DRGje9pgiaHuKftlWeQdUkGSVYl7PCgeFpGYurmY3pPX/4h2HEU9P+tK+Gk8wZr7
Y68tEYUE97pKT4LCMdeFK2AUPPLMpWad6/0/XcfssULpKPD+lh5kTAYDkZAXzkV1
ToPESmpuwhLUcrD+ATXS5g6tc7e2S1qL2J6aePF1QHn3n35Na2NSoM/3Awvo28AT
L5bCxSmiQiYO6x4NCTZcUo3REb29378tMxkw4GYvzrYS7YKhDUg5N4IeC7Nfla0v
saH/CjkyRDpenOP7itjzRaRAFrco4MdQAwqWMgZlZzJ/lJ5W141PbByl0pJJtV9R
ls+Q+A9E5IyJr5QtmiAUodRd3wWbOq4boYG+t2qg8OLyrOcob9DXa/7zQdR8XAld
707JhrLwIV4Qig0z1SkoGyUu3gBqNXg2NJsAdbUgXv98KZauKCBBX6w047Psgy2j
MCa/HF5qHatB0sdhMUkHO4Ao6tTaGrwD2s/uqaRN9othNd0gRcqdEfeYygEdM4py
8TGv7Bptvpwh0gddGDo1B9H94UW4PBBsGw2uhedxlRqbvf36QISuL1EgeU46wWPZ
h1EMGidfWJc5rqzPOnLfdQAbiZmF0UOxZKdBwQrJhhABHl1y6UAs+hLiVNQ7ojcb
j82RfNjp7SM6xvxrLIC+juBgWWg74o3mogUCbqFFf4/Kek3HBV/mumqnymJgip1l
WMftjA/TxMntDdfL9099iF+RgBAlwPyZVLwSrP+Ec/suDVPd6BafZ2tWLLY64Q9R
xlTmuRmoJAmzUzCrPkwki6xxGlO9JJPgNowh5QwScWL+PBgito5bT3dcUPTE8Uej
jE6snIOTegvdUTsLucROaYT6LeTLFpySZihLGMDFImGm5QjaicBBjzIzVoBaA4fj
j8d5FAFM6MN2o8FH0Nk3Ze649T3G48TXJELpuHydcwevY0C/LXv5Ppj4WGK0udjE
nSGUrnrNyO2w5ROHAsZdSD0L8KoWM6Ij/DW5fEzDi4v/ra4m70szdCvZP2LltZO4
fNuoH1WI3OPvBjkPoXx46PkrGFDvmqCnmtT6csT3hOhmxHsA5GrZSmjvlZHyzW1X
1Tf8eJGU1ia6UqE/8FsjgeDQSbFw6VCrY46JoqYWjsaI+/YUO/k5GD7qFCv/PZin
A1NfAsGdJk8S1QcbipLPmpMO3+vlkdayBVPY7ygLM9LiVfPwuhT+P/UQmjX7Zbsi
0jFRK1DTImqLpnlnj0/VHQaz8FJ9w9y0qd8tPegJduiNEuF3XKlUmbGz5MzRbeVl
FQ+v7N9sBckK0/1jxMPo7I21Nb7Twz7kZQN+l8o0zGsKOpvetI/c9iubae3/w0t1
LjhJfl3KjAAdGIa0XGAKR/7goMY505Lf+SXQadfiwtXm5sY+RzLq7+YrM0t/QXjs
9zkl/gH4uJ5JiRbX4t7omFOi2FOBa8fwlG38zdg58K9gKLyeyBKtFnjTPxRua0Bk
X9i4xjLaekuWdee7LWy25zkh1VyZPz5yTDqBADBA//rJueSlc5SCr0R7kDHtP5CM
EItxbWByfEiyl9Npp468tMO4Zcg/XkYTslQZap43szdH0Ea5rb4IQvpa7g33/zgH
g4VIOqa0xBbngXL80TWvKk9E3i+1lEU7yYIRPImgeRFciS1a3zEQGKRbobrdB6oe
zJvvcdBn84DkS6WCAT7u5AJzeN+NlZLeX3ICgHo19h/W9OlrPqpddZ5KGRwPv6sn
oaeS9fC09feOZxH393J718l7bSulypl574QrRI/KBkpZwCNx1SdSaYBpzqItt3oB
A6yoxxDA4XbJyoN1LGyWq3tuLy59sLgzw3C/GvUDzrc+78svyEqTS6kGP6mQebGW
ed3BH6s59AWvrAzvwnZBN2I17173MIoDPfrq9InnPokU759D5PzcSZ8UTh7tMRm/
5HXZoIC8hT6XEjkEqkkXmzrhcCNU21LI7C/pkZIrZ8RR3OPgqdYnkVuw/wOta5Ez
Z/A/+KPzZEfA6CNs9Xe4OycJwURwnG09eFE8l6pDtd/X9KERCj93ZB7GlRxltWvr
C/KCFP8SIPUv+nLHAU03Vrjg74wuC6McTT9W4tKhcHph83gGzr3ZS4kDum3H+/AC
SO0V7kC7MV47R00wj9xvSW14/X3Jh9U1MoDKKDmGD2jI5ewbRiL0Ig3akmMT7WVY
LWQQ92L6LI0dlmqWGDrQWZ9oBU4IQcCpXsP29q1JDS9S/KL8wGKAZOYdcodqWl1C
pFwhV+ST8hfGGKfW4crzdyFHDAPoYQk+APgsWuqSlrQ/sU1WgCG4SkHaciCdWYbE
hQtdYymOjEN6qcufRicd7u6KSopu4Y6SwuLn3yAySjy+io6EYDirOLKMR8qrflro
tcOLKALpQVFyXP8zUoqEJGb1ZJ+sSc3GHVAyDKOCsY3tCT82K1Bxk0GNMP7nNddy
6F+HQ3U4is45oMUPT1VKoUieuNyQdRHiKxbCtYpTw8wNVY4/EwyqGrlkngfGUlPv
rlawzKNPsTdH5lyaBknF0IGriiUdpbtV+i90Eqopi5zVV9bdIm3+R/0ftDO1XlNP
HQPPysmNEjVXgi4XONtWa7BzT7qUw1W0McwPayH5rB3pY5mLyxzDTY+llgQpnfS1
WH9T9vqPeVW63sssWSh2XqulMDnAHCZhQODQtEY+pruHbOfEkL8SoRGV7AEdhU1J
QXlazYvrxWlPTnQVT5/m+gH48nsHMPApxAI80UbfBB0h2rTFbdqbDtEIR9TY0NX1
TSM/huzvyGxFGLZQfGRYpasoW0agYUXiFIrGx4+SfxshcQ3A6gY8Rwn5UhlbN3ws
d0IXXNCydPZl+jeIO55b7iJ0eThNiXbjRNZW2MayDdI+yTYppbPVe/GvspEDmrLa
MQVyXTodMQYjgOwb8sRIM/VhjOOnFTjDFDTV3ZFk868ZPBLt0FALHaQjPOas4Weq
VUDK4BNq8Ej0sUAiSHpHT5a4s3USP90B3rXTcKygZEPeFQHmE4CEgal5x33EKTht
uo8L8+ovaGAKiGhnNDnS0hE3hdqG2xf04t6MVXOp8wnPjdVbCmeXlefbuEegmTsm
37F+d/urHVeu7mlOTQLJOibEyoh8BwQM4EOajLzjDLlX2VWYfvBM+DkIH/tW2VHr
0jjt2otKHNGLyTGQPWPKLX9AmrIa8hXYEJXFQkJFT0ccvgnEC3iQblkjIjO0k5ib
1XQxfL6LXLX1YnauB/JjIPBt0mHKkKJHSY1u6SdXqlyC/G//C1cDsQFnyDiffp18
8Zjlg54YzgMpJJeDo11Rx9I33/vewFbH5juuZVpkuNZRNg1DkZeIEuIlw1XIRfK/
fG7jjYN10YXMfFsl+KOntUTtgprkWU4u+PzjhXp7watt+3DlygoIybNgRbABGeov
ktL+c2wUZq/LSFvZYACG0ZntfJ5uvEyDawnHJqHO/sgmqTDxUzhv10Oa3zgt5avo
ZTbtrjMKdo1Q8XvkpW76p/cZahkNyf6n00CEPqGOO9Xg3mghPz2wHcLITRI6jdYt
h4XE4WSBY3vmV7pv9d1/gf5/yHZofn1QxZopO2SUX30bYaa6o39cBT6PelSw4Ho0
B0OlDhMEm+ULCfb5Ow4Y7qyhZTolE7LlGmANORFka98S84sKU0wfrH0xrtGR20T0
sxWSyafP+mAZDMrdBPlYpkz31/4n7JOM9BMB7Hg3jQGKJJQV+v+ngJRHB6ji7LS4
ln3W1eOhwCWpXDtHuLbw99U/UAq30VvRAc/5WJF0Z1chgccb9U4YX5tF/BDa0gRm
/cTW90Umza4ocpMleUO4NEq6mWcdPGQ2NHVwXGSScZwJPNQuMqFGoPkTXHDJIRuJ
okXLhoyIi2/wzoA7H19Of455XtrUJif15HfvChuZk6x04FOgouGe4ACW3RfB2Coj
Zv7Yb45joYgkEH3puOlrT7bu0KL3uaj26Q4hCsfMBrYnsgMuozBhEvFipA8+phWK
wrwPSx/9bpSJBOzrFMMUejjTVskPm2QO3f4S9Ez8uYoE6bF+WmBAU1jKm8oB06N8
LVdx9OPSTVS3p+uMoRNKh6nwTMWPN6zKV/WqoVhGUdiWdBt7z3jjIa4Ylr1yB2K4
r/BXChBXTnD7+ebULsJgiSiRWpR38eQPP6kvEnfwfzfg9tdTAygEiWX8jZ92nO94
eR5AST/6U/P5Na68OsbZDrZHPqf/evFDWLIEW9sgugZaAGuT3KY/CWc41/ZPhkb1
TMt/AB0fC2A9cobXPCrJtiWb4USq2NCn2VwYjeqP8Iaqw08m/DauViCSKOa52mnt
CxGQI2LGmXEmW8wn4D6hZS49+DsC3Lk1dZey4yjNPxBURFKGE7VTEhs6Mq31aS15
+RE17D8ixHAXbbpIRe2jQaxfxPUZmXoaLiYKmwRqjAlN3Kx3uc+/fnrRfBSgeLRY
hSAKWBevb6YQ7XSPBpYUhGzB2Ra79WTptTVgy3WqnckQy7fxABzHcgAG2P7ImQFf
4lT8Nr917H8gQ2LrSBTfWEz1+wpu0IBd4oRgslrCk+PxZqnH7fkIC0AIqTkYxLoY
mOXNnxaa4IQEJ1ZiTr4u6zAUybN223CcZH6l5nFqwMylDZTi5N8doA7P+7L+pRpY
coFapxBQCarsDY5htoMgWHeV9jKWcrWLuk0FKzVEzq08fHhiR056SynJkS2udhLZ
D4WoYl5WKmTY2uab9C/r4X96g8vxBKpl0FBOdZAppJFc5an0ErHVv0ZyxmLe1gL2
BZjqYk9mTJi9SLbcugyVJhy7KBw0QuX231Yz4/zkKeGkfp59J6Maris1JxVoqXyr
4mhl28jARB+57qI4Rh6qtDlr92svUe56IeU0O1fT7N8c35LSBVBPwwMDMD5T2SHm
QI2jb1/cgOxk+KF7rpPjxhCoNO/f8IKFwib2ARd8gisa2/tbMyrUvBX2fkKA+FSJ
HuXnnAjo+ylZ5ZZXR/+yFQ0SqaVhDwtmwFzXuXdxyrU47+YdWaQ6UeIXDEeUGZQi
ybC0yDX3ewx037UBkflUCxJWIaUshZHcN/VaJ18Ey++nsI1m7UuIjD+upo/vuwq/
j7LjXiZ2ffldQcHf+8sPeUTm6/G0JCF+v5ylHGUNlo8DkpXdXxnSgOC3YXN5Mck1
f1tVebAvzk8WfoeMRHyMD9ODyNtOrNLrbcGMWxYYj4wCSx55c4UteOEpdiB42/kc
h2DAnbY3wxK8qXp2iTiX+nEqOOZLXLkCrIvv2ko6zoWIxwyssnhmSHG3tg9JTJVz
JO8dv28z2Dp2RtO3uyESe0Z8wNFBSzaCei3ywCgOZ/+On97CiuL46j+3/2z7KGZi
3QK0tyQRbRbe/IX6HXBNGpkz0AOgv4HIaGwh1wg9gX91AdjZ7u2WKaMjPLlmHWiZ
HYsgKITWPwC+s62BiccjmjKNg61j00Yxl1ISUFrPbVh5ekcRIBb7p4wBrvQFaaJd
9PmiVs+Vq0FdVs6MaEp6zA79Bcr4yYq2BV754RJthKDoIyGg0YYAvKbCAcc1sxsN
NxVXu3Lr8c3ne+es6D99vSani7h6BAH1d0DeuSX/oz9DfPpw0Oa8kuxfSCyTvMn1
7wQet4Ou9xNSpxufJXBF3pHeQvCwQgNtr+SKjqglrV4oB3yHZ0DqeSbMIYi6HC8l
+cM0jAiByrFkjsYbSqGX6zIqsknDr5RZpfx5HrODsSHyhJSr2edfo2sK2zO3w1ni
hAH1lxLIOnzFcvl0PLZCo8QbKFSBzdG7VId7JJFG99yf+h7HKDE0AObcgYiHuwG6
+22qOqBW+YySTnSM6ca3R6a76e0fELUzTlwXBIVhdy/+ZQmIMH9ffn5EUpnL9W5v
eetXWoJfP26eFW48uZj3jbSvEQrAutvUJlf4xfCaBUMMmcWj6jgwMgFOc1kliPiq
bSiEHh6avDExc6gcJP29lsgQlKg3FdMK7+Cpa6EJnjnpTInz39cHem0/KlB25ahn
koaRrxRI5X8cpVG9VocGGls8HMXXL6SZmaiy5qSENYQhLHEo3U9XyyxrnW1Wb4Zq
H742mr/bRErrIPIaO2WHn0vaau/Vv3N/6PKqK+H8ocSCyWi0XEEWGPviYuwAGf1a
tCbpBysDFPLecpou+FNEDanLQNUzhLZ0atyMJ3G+T1JcHBVaSl6Fv5HwVZWMIAry
QQNSwALppG/AMJ7RwLy1i4Pz/ZKHAcUP8p+Uuwjmb11aGw6uLW/0fWjUIzcrfyU2
nxoQPREl+okEXvifoEo1yuI92Z62qLDJuVMn4sGIsi/sz4TYIuHoyumfRs9WzqzH
oIZCixKKsVkv54K9r8lVThvDqWrUccu3HT67fEHgliydt9bes7Wxl27vAzUqNv1e
/GmxjDjijUKyxg664SeA5xYhCgU4lAgFcTnT7pcbsqJ9VpBVzCEU2HvL9jf7eZOw
+fBweHJYzdzdblrywh5ig6UAGm+90ZK7a1xPWC3bGNWW5hmM6jyV513W3m+pnuGV
GivzeZzwQ8UDkCIhihP+bTeDiZhQG0g5adKRuiQstvcqKNu+ccp1ZbRdHpoM30Pr
Vmsqn0SAb46grmXeAuYNrdTQIBKjtMi5EcL+YN6J/n8n69ug3iiY/rkWjmh5o/cY
TniEosYXiHEQqip8zGtSaPGTo/rMLpw+seOF0MNtukx8C1YEI1oVPBQoXP4jNqOk
eTzAzVZxWZucTttxrwhtkO+lC+yNsYJ6efCINsxDUXuDOFZZJ0I4+VUL4DD/vOR2
KGOrBtQt9BXLaahfSzOXn2/KtHq67koWUpbD96NvGbY2YH++z6AJwJ+YBqFYx1+Y
NbIUqafpGDBhWf0nObyxVDQVUhkxC3aG6FXPtclg+nk9Y716oX9hE7I/tlRe4Pwb
GFDjOUScQyWmM7f/NBgTmUsmq4pkITRMJtl2DklcGOkfGHVSWaRMpIInIcY/zxx5
h2O9V/fOtYsJruQhW1lGD0+VO1fw/Ea4gD4gSUtaBmWmTIHeWltfWF59E5zzDuqQ
FJ0ZbiAVgLaSFJk/8oUXcyuIXo6eWxiNGMsVoceKbycOwrTGWfSPOpYfwCB4irfU
JNmkdUzHDguYoTebRnRp8+yE5d2c0SPcNgjbhaAi9WVLrXSgTIOxAP21wPu1q8Nm
+sdb/EVK460UEd0nXuRKa0C3DYqdRpOOeWBcls+LqXKYWcbEHaYAojfFqZdFZnXp
A8jtjAS/emioe6+nHT5POx+bk4uy6VTm+epwecRX7BpSVWtF2XMdIAqF5FZlrvz1
wRGspNslbgYMRUSHRBTta/3JUelZpGHkJszRwbEWedIonKvDdDAvthT7uEIGsdF3
SSGDlojl4nMijgWTw62g0UQof3BjpXV1gsT3AvzyEuEMQh6njOanAJK6y2u5xlcm
jUdsQ9GFoU13rUPfMK9J3/vrIryxeBVIwWMWBOOwg8xRxz7vAORUn/F1JsH0KkhJ
My/EAUfyJGkQQBg5f87siA66LwPlnqwXWBzo1P3sPo/ENfC9PRMRJKBshASkOPUL
Yqum/YsoKc60ED7OqDnV3G+9/JmqVFcip3PYl7uS5lzz4yGZNK/ac86H31jlPWuq
r3TV7Oqyu1oJQCrJqJ4YQ405rnp3z7th95Yu5o3AAVPSR2SHjWn4L1ncLs6rM0nZ
AMnLJSMqrnrIzPZQae6N0xJV6V05oZJwkhDo1baP0gRAZDcY8gViPPLPB4/zbgBX
kwme67o7LXri/IMCITquddTvHo7DISsy/L0owbUOvxWo4ab7xKWqeb9roJAtisu3
6SDPp+i0+m/Gysv7dMW4zov6O5FUN3A+uV/lKKYHNYSA0bnUPXZHmaiG8asLyWz9
1e5AyvUHVJG2poAEamA79nnspyMtgHtf3AmzZ8IhGMh8UcifnwYQxoyaXKGf75F9
5YXD8tVBSWdvnZI/yLs9VzdQikcr6w47T/RzRt7DM1jkJYgi6SiMjcbNLfyD2X2X
XbhkYPCu+7IEp3U6G+HXK4UlhJbvvpha9s66lepb2C2YP5kT8G8yg/3Y5c8tK0/J
hOUa6+9gtLmok9ZDHBhslilvfjVTlb7R4eJszT3yQatfdByTCycz7pyqRhHqzZIt
IuXq+3h2CbpyZPqwGtIkZM2DzKY0aa8PLwC2zIO0uAio4707pQMlp/bLFoil1VcI
2JE7CBGpXIfSqpnbUhEp678M/gm9DUnhyEXnJoOvPd+uNNvfntOY7vNymXKdSrw1
SUYykNnqvZBAP0+eqzqiSfsSPqhA9P/6vm2bOZigfzZy8vpzePs17n9VFWf3Bz+a
dXSRSXK9N23Noj5vreiSKLVM8vwKBIUjp/kVyNlV3O1Eb5njhm4j2UO3OOlvAGHs
wVfGfh6DpF3KoHm6tadQmeZztjvc1x/NyoVr/qwAEYaZd/9GPiTZMfYjaGXTGOd2
o5hackVajuj17VRuNxc9l9+rFw6neJLPXx0X9ZCXWNIqYy3my/TcWfkB5I3uHN6i
+kJCsUB4xB8gWljCeVJ9+GHaJ2fkYijQMnOADRh8OrlxXUdcoVfuN4DFh9OY2WXo
TsNdRgYhl3znusVru9tCWweczSTE8a28OjvwKDgxQGWMcQeja14nyG3RDLzk3gq9
PGDuurqU7LARP/ZTlByfBj/moCUJkElsTHRfFBEvPeKMB4RPNBNA2Er2A3aN/ITr
YkqklsXL5R43k0e075ADlnipQZFP5fcRm8Unwc2Ik2KC3kYwizJQyCfkR82Gl0Mh
CbUz9FTuhKvTeao/o4JByTK14n9v8oEjrqz5bAmNt5BcGDxSTK8W91MoHHifhnax
DxP4bLeUgoOxPYGl8AbzMaxZsZ8b36BpX1UOg9861Z6eziyiOL7Z+H0mwTghJgQt
038VaVoFoXnN3bfof2DXzxOSjgc6ock/oMK8aHDLv+cvmGF0eIW74DFu0oD3vxEl
NuC4H8u5vb4Etg+2ySu0Uf5BoMkm2fsJtYv724VRrakBPW0WjTFDzqTDJETybWrd
yZu/a6/BKbncify/I0NzPLwX9biB6MQgSR1smlLrhcN9vnbtlb9/El2lOCaH4vJO
EvMbmrGE05XdavvqMwaQ8gxLQ/UEV89ttFIkpxCx3TwEkQxPjm20PMc2cIhDWgoR
Rxnxe+xd4b4F4cvvjrCxwwul0TQ03Ntb2cguIfwX5Xe8r9ZojNxjoJehKGQIU1Sb
1oY7kS3OIP2tj4ClguyhrXQWB1EP4q3+9e5hyzMpYkWHdZToSgE7QhPctzr/eSGw
xe6S/8gan9WzD05oE5+XMi/cy+UX5zZ9J+PF+Wqj7gpm1Rz5adOdbP/tz/D29+cd
bUpclT5G/OAIifCIb6vabrBdej+Ugsq0kQzRCYP1+D1IX/lALaHFG9n45NcvQTa1
KVztltDJnufP+TRqYfqEvvTEk60gyomDz05of2ek0KjxYFrINTtoeIqWtmlQ8STZ
IWma0TXLMAcKk3nHnVSfZV+2V9KhFG9lAZkIRz90m4TAR8xijxgVHVYr1Cc+3gds
KyEC/xJRHBT3aKO2DTboGg42OlYYVCqgZYUlvYU+ea1fIc0GOSLFQ1yre1prjpwE
O2V8Ud/09n939AminDqNbSM574eTJhkiDD7eQPvpuQxup/23FbDnS85k22mcoVsk
fe0CX7eSO42iZFb5J+j/ze6m1MK7HjzQ/d4qYW/pd2Zae5vjq+eu3Gxy0MtgmpO2
XrhtOKiT9WnOPckG9JwN4hRaeucnBYdmmltpLOPhkv9m7JBxc1/lHsqrXwJZgk8y
SQNpT43ahSRr2mL2CuRJS4C3O6ZsU1JTn7HASTbrLo8HbA052gbYOzyKtc+/dIko
hYJXdLgqU0Iz6U47I5RPL2hhme9VBuIfMY3ptWqeNz7t1csI80JjZcuKUNcyTH4f
0N4B/im7Og2ere+16eFpXuq1xuTowwSb7VXCTD6hgYnxW4ISmVAydVJObhWNw3Yk
iVDLD+FeEfR32Doq/5D16bbNCK74kToZbe7Kcjt1RhhhE75L3DmRY+llrMylb/vY
/ovO+jr4SBiw6f6QVUNZq8Ru2rcziMvkezu/TtnN4XHOOpHuYrBqa+0ozs/ehy33
JDnRbuwBUJyUF9Y4NubkrAhU7sa2oXVmB9LLyUni09gQRHHtCwgrkowRYv1E4rpM
CpofNpd8+IqDYH+8OmUUwihs9xgHf4XK/EwAP8YxKHzySFhLcd6vgaE3Dpwj9o+w
60A7JMfsxA9oJCQ9nNlSe7/L2LKvLprYjXbXrSin7G3iLTYdf42AQc/HW2r6pc4m
e9hqOwBWGvCHSGGOEIlWa9nLf457zQ39cl9/1ZjJd8LXMf1s2dtfxDKQpB1JUqON
MqsbddQxDsHr0zYa2PD8vAu5SuB1tN2/RMHa/XIeRNRUGg0OyWeL3oOpkbqBf+Qy
BU7+0+bTTtHCtoTk8KES4TdcrBy34vTC68dliQiFKMuYGLmcixEkHxVLhcfcCG+x
cCs3dHcTC/19gIjnIHQlGRGwIXsuX0Eab5GpPaPpvxpStI3MQqcL1FL1C4bkrvo3
0Ya9eHcWBCwvTAZFiIX0k7Ip5OX2ezcCf5hi++S9TD+QPLyiPnDF7iSlShSHsGf5
PmHEY+CkKsdelvw/C2XAPKuaip4ZALSzQQoxKg4gDtRiABS0siRSb3dCQ00Maufb
KogzVBExA2YA+vKJ3z8vC/zSP19ZSXDgWolxukP7l8vtztbQCayhn9SWZixecKUg
SRH53UaQGpQFgqQlnDwvpZ11RJ4eXn2Kp61xggvF9uqvu/nlJ2pG2JqWhXIM4QYM
7bxlujcwpIyOUhJeHCpGJOucPhPlBa1Zh4AsegMh9BBGdbKzJss1onHklYeGnJpt
1kra4a48adCW4fHTtPPKqRExdPkGdSh2VXGnKLqtfThfyAw2Cg7zHscHQE/V1KFF
sDl0y8LO7GHK2ccfeKpcAiTeqvMCnGmrkW9UCT9NGa1+Vgo1hFPp2VdB5oNAJ7Wh
265vShlkVXez+tWQJmpna4uEYpsDedOMMsI9cC0KcRCLcL0WuXUs1o9XuSmBq2fk
Gwfqldonw5y5a/80yRqDaMNTt9MKN/0hMjfpgNuyOMniqsbD600iBSZQYiwNcmAg
f9Te04FSVmV2pXnxd+Ja7Xo8KDP1Rx+PM7dcqptewZimGGBvrmwCjS8i/1Dw2jKq
nLt2TxTaHipJWvm32ERP6JYDTNcxInaVpMYbYMenTb8Ul9g5XYFOifpfzhHLEVcu
q1KrjfREpw7nUjT8nssRrpgzjcaOlTMIZCrROPh9Id6NGzMNzfINd8OWYHDiq4zN
c9fgSALikIGADoorZVMNbf0xZvA7vCo0lcrH0FLqs4t8e3tJ1YRPHiqIR+BzAPJn
u5rjKTaelp1gbGvkQTDVsIX/tOqnplcfTrFsBIpHv1T4jT0cVcX7jE0IOheD+32S
iJnEOwpY/ZrAHs6GLuKV4UuLSlV0OzIKm8U6LmnAPDrNwXn9eDuCLOlf9Ye1cUGU
y97sXHlErohMNQfpT9PTv+dCD5tWFik45sg/1zrYpHWjwqpn4k+5L7mm/1GAIlOZ
Z+pLuhuHn4JxRkZflRz7R/ePTEesDGY3k6dah+nDQbGKjdLYmMt8GwgrfJUy5j2k
7iO+X29wojZ7aAis7QJnrCJAoiaoka3lnn/nny4mWkWLj7mP3bpp7sR2MmCopZ/4
TeG1Zm+Bl9k3bQ71Ww1X5Zc7nUQT/W2pdx9JRzMTJZD0TgZlyTNwcz4l7HgM72ys
ei2sBdXDob3b+VV76y18UpS1sxTyqHNNHS4kiWdf0Fv39ocpbJZVQC98YITCavXq
FAg3cxxKCPxxO8aVQb6pEskc3a109rA9fI7z57iwuusR0dJD3YORk9gUQn/qg/Xj
m0N6rP4wfkySZ0D7pCBosMYai/3OxyX8LD0D88KhKEmeat/zAdhnxcAVnLS+ZOtq
+lZLr8AucykOcrKcHwRBun8wo6OVzSFOGVY3ataJ+Df1GytTbdB5IA8L4v6nCM0/
zIjrOV/ZeQUzTLJfJReodIvsraeFTlIbW2YvBlwWd8PT37LGUAnRCo2bCdqDRNSu
6dMDMrknzqrj282GBRFHOfcITuM5qpdlMYsXYtujbA0P10o5Movls6o77HPFfekX
VLQuEETtOg3/+oMl5Qaf/MMQqjvPjUkvHrXjRApjTlsA/Txc2faWjP4eN3jz1q1a
H2wTwVN7NJbA+PGg2VpRpdo4ePXOIuhNLjh+KvfCA1BaQv6DMNAACfOUsqqo+nE4
hAvnODcdVPVGi1Wr6hbx+y/6j/1MiK8sCnlcOsAeOzAxMaDgrnihGxci4VobxUXi
T9nernXV3vVF5b+TVq3Pj5eihO370vQ447MiCodRirKK+3fIryhx3a53kXwbvDfg
zQUZ7zXCx9tIKsDj4jBEcOlQng+qTiU0ptoCJfyS3w+Sk01uXf8sN4Wy43lu+5wT
IRx8RdbpqVGCLTkOQboTTNsxnr0mYizm9Y+OYKVnpt1txuSjTw1frW1tHnF9HCy7
H4QWbj4uHJNINvVxYhms0H5bZKnAJ5CE5pRNNbSNjlrrRpQZzTm84cfprsRi1lKS
G/TTE/PKuowGCH++Iifn1UyvBhf18Xx2Pb5IqL5Cyf8vxmcmgsbfmLnFcoPd7K/p
88vda1JgUd9t+gWn/7/iIj1iGh1P59CxHuIIlH4Gtqd4uF3XZ491aq3OQ4Ov1Xev
vJ3IaRQ1ZMF/mAsEyMRzQWPlERrr0D9UMuWmB4iUk50XnCkMRolF4g9npqzkr6Gb
LPZVmOE2pDmSIpmOIAijtqTlco0V4XDLiLxdE14Ri9+bCnzZTJXzLXyImDWGjknZ
CdCJDjhq7QwoEE6VCKIO789MftFqHpxh/Hs1Fao3m/S+N0YxFXaAAEmgyhO7ZRfN
vf2Ttjg74f3OxtbJY5OOPKFVW5WkyuCspIetYispYd9lj4wDH59YuhNRuLz/0JV7
f023FuiDV37pVvRw8JQ6wZuU5SyrFD919NEw6gVTgosCjFG+YmR5/DE4GbBvyuNL
SZy89FYx1VWCfbx2BMXgpxY4cANUpP264HkSy0Z3LrzJJLLEnsUakSqi8FREVf7U
hnrzMmIddEQYFZAs5G62NHX7VIYvKS9EnjLUikUFxIInnNpjc8bPSzqY47IRi5LD
DKrIPE5uTWhmGcp+/Cyb28FDWVH4Ubb+/cQE3tdO2RLJIDIKGMqZ3Wb/6loZ03Ln
ZvdgaSSZULhaqBNDeEa6m5S2PpEIJPCLNSZQywqxksYh39areCHeMtxh6qMYK6mh
XIcdt5ngPbwGy14HA8m+EQz9ieG7fQolUkIwV6grPbFPDD17t0FMeQo3Ctefa1fj
jLtvxCm12jVqtR8s22y1Bk+rAot2Zn2tOjvCahLJ2lMa29d/lbYW0opPnAgaHVFI
Qg1UPrG9XQ/v/bWXNzGuhzn1xuYSKrIs2mZ6L8bRHNBDG2MbNwhbjnECojHqpjAv
7yPcZax3hJuyya3Dk+3YLWcVcw6BumWIdDImra41v6RbFzBsHR7jgKE6ltp6OFEN
Cfs93uGwecHYKHnOFEaPmLPYj8yvyqGP1ksM5dvTZhLd3yzV4+X2+NcQx5Ri6r/+
2Bf3829lh1/msWibyOyOnsBB0pNOCqDFW0QJzg7dZN4etX44LNdgSH9a0FvmoiyH
BwWPf+6sKXbgOagGvklSrc7aKlApfblmLeNMjShyE5hEy/3Dy5HQYBAvBzW9bC5R
UwEjwEOAVqwd5y0L1DTStz3RPBgcKGZVI8cXRuwQrOrIGZHt9S0oRmGlsx/I9ZS+
+m230cyb4oLyjcZ75gfS79DDr1k+9gs/YCCNIFONAf9A90+o037PqREM5dxrgEm4
njaqmO4y/C62DidpaPpmRLytW1OkUKV2YXdZ7bXmaoJXkWck3JnNX+77OOLY/4tu
UW9lFFy6/fJ3WovuhmfOFZWzobJG99ZqmtuQQ4UinGMlClmTp4XkksTQM0t2wWGD
wbn86lEIGndLBNz3wOyHzhQA2655d+yCz+sd01XpposyeFJpILLCB9m8oB1AB101
0JKlRKsJTzjlOGIbplJgTUcxHEucYu89MZ262swivWOr7HnLNvh5PYEhHWQIqooT
Upa0TmUSv4vGsYr+M7sYngFGZ46/bCFx2ywnwWNvKprXMzAF/CEdnkhfRaRT0ryA
qxU0y7J0RRSmNdGCnrcm9Ptk19bqb+Oqo7EmpdELznJuoe0n0nh6VHT6ke8gGGH6
uh8fsVtzDpkXQN9jVuYOVaXjxWpaz6hEkTDwkDVKUafBBDWG80DNe6exc8H5svf0
Oia5fpeW7kzJjLV7NGf08jyrtvWUFc6D9nEHk4kCbFvgUiMUHAN9gThspvJzRbyL
5Ue2O+rttdfQ0HKnwSyd8qJMbKItzuXGjhGwSSSNvZ19+Ga2TB3jnihwNo+h2xV9
wKEFWuFtlc42IiorTBabeQOE/JNurEN3VW8bOGiLqXbeZlhtda/Kwp5z5Z6Gf/0y
t4Vgy0rR2oskFbFEe0awSRJIAw9/smAC3QzEYWoCjNUnMTAxy8kGMWHCypeOeT+I
4rIhlaPa+wkPB3HHILMOOETSIaz9ImW0zfgpjlGP6VyPtcgJDPBSx/gMulEI0mvK
eP8ZI76BrXRxstcHxAl+GLpMmySgx9VuB7Ql0Yi4W5abSzCJmsdbS3b+baP1B1Mf
Lig/iAzh4QsxJnUw54J8vInO2msGjO5uQIkif53Z8oh0HtbP9jnoPxxBu8E+wHeW
QxM7SIIzYdgfA4oOmP2A987Du3Gnq1W8PrC3XOOBoecQnSArg6ESNE37O7cZp7+w
pUcAJBWZOWhm4JjuMNHTC7+W3Gz4tot7zhv8rPqCQ7c3DguQ9Cl5GhDJdhjN+sIp
KP40SorYYXRgoFpWi8Y33P6E/wx9ihREvQ98k/3GGe6+jhwrnLQS9riPwwge4JXR
KXo8fhlEtwZIWPPjN9kqxwpdFN/f1a44wDzBNYP/W/F7RsdDh2w/IGzPlASBdTY2
TkUYOq0f5WBUFrYCdeZiXLWCdk861Xcr+Von8kiX+nU4PcrhYm9n0v7pGRguIsdc
C2XkWQaqGLejodP+RE/eyORnB8O1rV8LtA2xNsz6s0nM8opaU5Tl+DzSRuzK57o1
ESPkBRbeNPT8uXZvJuGqrme5ZwQss2HNH7XXENZ8ZJQTA2Yk2IiJcjzNjQ0OvFDA
7wlO6cgVLg7ER5nxcLC6soDuzc4hZ+O2NubMvr9Zx414WW8o65dlQcRPbwnmflNA
ueVh1Yg2ACF8vgY/dxtLLDPLipjt1IsAY8s8JgooOuOz7lpKdrHOgZnkVfKV1gC0
iGc7h/+ZdIYfTZZNRA+ZnsvHJMVaZg0fri5WiDzIqmZ77tfn6ZGm+h1nHDTOpRX4
7WFvQG95mU9rVy97Ka/OUPgRICOIk+fPdZhqcKS9yVvZups5OmacQzWfQ+ezkMxX
Eov1lNzPSCDBXhl+0lSzbuSJ6o+URqJEl2NTwuCrH2lRD1kEzgzEC6iKpj+oIJHS
6q2BIx2Xn0lS/OP3bK52EhXEFzisiDsDqBwOKdAu/ITm2eEPyjnHBotoFa0xGdqm
FTVJlGLaIY6snNokvWSLSgPgnXPwjjzpYO6zDLrwv+MIjngfLdzb4fGnX7X4waoJ
WkO25LCIZxqAvDEnOsmkyLx+jtlHhUliIyXN7ZrsatiNoFYuDxwrqHFcYnhYsXJ4
ZxRHmqlfNZglFOybMuySFXwnm/MKPLO8uA/NkkOay1/9lPL1I1CIzfdboiIKNMpw
b6HIyrp39NMHkGiK51BaH62TxVRIHgWD4KxqsQSOsxv43IM00xXQBojXI8WjcLP6
wB7ss1Jm9mC07c8A6hzSpbq5oYsHC2CNRwCtZCubtrCHvRQoflKWjYlaZNR11gv0
IfsugsZn6xaHDlveCphHLjBy+cirv6SAX3OEzHUNWH5vYbQGEftqhVxs0rIBDjCK
/9AN4T1ybXzv7X3DmgBxaQBbgY3BpnVdA/odiqbyPa6Wm8JVvoA+zO0VmxGefsLq
a8XyBziLz/OIcXYbsgjk5cZOrDiXGIhlaTpUoLE0Z6QU1V/p8Onn6Gj8D10ti8Zf
/50kbBO8MC+gdhbJ3BOFn4n5Gv+U+pTOlxV1SBjSujLCBltsxjR79IWTAEgbg5DM
D2zoC8sN8/99mVjstjuPbzIyvD3cm8OUeACWhLqdtQ/qRNd2tW1OeWOaE/UNwF/3
wzA3X8V+Rvlv8dn9b979OLa5/Bi1USquUUbI5AI+Nifer94ngAxdTtwe1KFebzFK
mCBHgN4mfP5X6ObvS+GdoSPTg6wnKwW207YS+LCqmFpOSxtMw39oEqz6IKKe4iT0
sAmV6sJ8KMeqHAXI8zCX/at38bJ9Uv47k81FriNMPc+5GXhoUZiyzS+DlNidefXt
YnLWrlws+4RFoAAw/R72OFCkZiOw5dZHRK/cbAPMh4VWD/goGbT+yJg47h7dJJAi
MKpGo9a+0sIz3Dd+BW59IRKf7fwEZlqnYBa2EFxhpaijowpl1Gv9/4JtR7e90tAX
RhTRS3+VFvq6exiAEho9AJeBCdOtySEHjJejltToYQ5IlaWZTgmHrkjFPj9wb9J6
IIVcaZZmGKC24m3TkV0LeePn9IiKWqNQg6qpb3I/WIXG5GqckistfPi+3KxreNCP
I1yxE54m88ns0xo+oWW8UbCPXgYe+3aSvt1SUFqiM96MamqkKIKcpurUYfHLIfvX
JBwbD1JIBRq6aZqjLQxht/+YjT50qGNa7ZyGSkE5eDqsjlQ+MaQujaxhQwJHJFmg
91SA+1CpByoTF5yOLh9n0VEsFzpL83//aTgsz5sRo5uE5vYrVgJgelbM1rFyaJ8V
D/jlYj/DCudVicv/9th5coHfGm4eG1KDI4BZnKq3d+RHM+WSYCgIzFWiEIxQKG+B
p2tnL5bwma4mrdJgTDFfNOraaFoXzoRqmQ0l9lYKbdxNc952c7il30zCNREt5xWq
PBsEkI8PQYuWJJwYdjBh0VjE+O0de6lRdPEyBrgVzDtyf9Hhm47UwQg7YAsiN+Ub
tfWCojC20lQ/7LDEZie/N8Um+e1J11IvkYrGHVDq1SuBak+j9fwWVtmfOn5ZOryv
e2SNVfNsA3FOkaX8tkfkRJRG6ymjL5MDESpuPo0Egtvb65KScC6KHP6R/2Pncex4
MuS0PMI1NSuRT6B2p9w6pUxOZVHIoQdvKr9C9ibYOwt92751rdw+U8xClG7j11nR
xAksIhDSmjM0sMR0NSxoG8kpbhaKI28GtLY7FmqCdOHguAttQh494jl1kAkR37yM
Zo50W01j6BbcGiNU9qmJn+v+ahHsCkT+dLea+3iO+KUypjRtEOia9+xZGiZwaYts
Yzi/XI4y91RaZNOTkZaRbxxGovN9uIpaGN17+NZCn5HNZQbG6JsoqUTEOphcxr2H
FZDdOxQ1kYiaJafM0KFB/W8UQbhRsDptzebu5U4MuY25PZQYwd2n2UvmUl2otraT
FLg9/Cu2yzbCt3c+6kbVLZFO4MZUOC6YH3Ldkxkms3B3mZRimvlphqFhbjT2Hg1H
SMoLRpXdJokOOZRbLC7gChulUaO7hqOuTXYYc60z7QhsAhKBuyaIXc9wOiwEBY88
10nCPZbF9FmOkaRLgw6Yoe2F+xwFHDfHZpn5HSRL1sXns+a7bSLOfKjyAOmsmYhF
p0oq0AjaSrYxvMoG7klOvjTZFmG6CDWLX0I9vBkMuVH283QHGEIA5+zTeGlbDjFp
kwfwPrgvBb79woNADkEl9m0Q9bkRXYP8NgtGWiP2sK8ltEQOQoQ6UzijkJN4hHLF
NCkLA8ldHmom/t9IGi9J8gu4zIGUzp5coeY/b8AAdoOCgA8r8DY3KQrmZci/k2AX
SVUtGF4EHcEdc6cvlwmQmySo9BSrYPFt+xjk/PjTsNg08rItcBnScTjMSbnP4CHP
D3JsbIHjT6kuq/Bwy0Y56DSzBul3HsxadB4oIvDC4WmgunmSJhrvl9wPnLIHNBXu
ZIs1c9qwR/mBC5mXhDmpSPvCU+94Wr215V94vCb2OIh01BV4sQcYR67VmvJ1V5di
zlGcdPLENXyeXHfHk9hnNLVXlCi0f7mAtx/fnQMwb4LaYW08AltsyHpQmLAwaBga
Hi49nK0mtMeZ3pjGTe4ofAnMvYcHxrLVK4hWUS9XFtdkq5Ddfb3bAIpKPCWymqPq
Bq7mQCT/3vTr+N/6+05oTNBvcDzwSufUm+kmKyRw2YjYcbRwhvfPHlaNa/Nt6E/J
6Kpxw2Qh6GUBuHnffxCpIjQh159jGItgQXA7nemYEY72f+VFG9J73mQzgckqLxRg
6KobvTYv/APMSIx4SUd24b+nNnsFNHDDde9dsS8+uzgsu030Mf7kS4QhuT59RQ9t
q7+gs/U7eMrjBEb7S2ic4kvRGLf9tGQ9+el0VKdMQyW1mHdOsG77xEYWrWGzG/HV
QqY0VAjhbgVIYNHh9eY9c1thxh8Mh9KMF1ztd1SUxH0Cle+IJnRhZ8auPxvYh9jC
sred1fRD6aRzp5JY8NUBOV+gLy5YuVGyDpBNcRaXKbM93CdzDhchU6fsVJUdeFSv
7Xoo611Jk8UC0vnC6WHEE3JLxSB3W6yL3vSmbOKCSn4CTh+LPul6j/TP5VebZPoe
9arKwNXzXkUA566Lqhpm2AcXAXYaS1ugm+AEXBBoNH9ZYraxG1O5f4mpxglS+d/C
vtS8oRrFXEd+Jfb4WApN2zRF2XEawUpYdpixUBIk4p3kjtYpaOz17nSo4QoxfG5z
jh4xEnOmo/FluXiaKZh/H15UAjBPr2NbE/cb76Q12ermDkPuW28cjJ4XUBXD649x
/JCT6hFXgbaM2/fD4MgXwp1NlwJwc6PGY2dhvOLz+QzB7rXkNxBSPtUri8a6XUmw
z6MQClXBqk/6pH2cadRXmYmGrng/x3CEbdxoQ4NT2mVHY4ji8xYe379XqKniSn8Y
t3GP6EW10polGTwsxrPg6bSayBNewMN+rCf9WgpRC0dyBxPfknnz7rg75gpOCPPK
Y7Go3cpqYJ9YfjHVngScSbSiVv+W77lWgDEyaIdvGe6e0UyBeOHtfxx8gRgnGpDo
5WFLfi+EZwCzdPEeRxq3g9Xq/vwmy652xrwTTYmFD56K8RH9XWOzSH5BtWFD2b4t
8X5tx+nNS7tjgs4a4UrZr1gzSuVTwgrDkaCvkKa9g4f8zpLbWT6gaypL+/oLsAoc
EhsBruZ8g2/y07nhqIh6qBRxGHuu9MlQCN7WBDXh4EKrcaRDtfEXQCdWPNbWX04x
UEWTCmpMe9/nYDymktYa8GwFv4edeHyBdMKDNcTOLpTukMg0BZLbEbs8TDjcoaUn
eFnYIgghQ9BzxkevxgKez4jRHr9uHT+Tk4c9jCWqRDJVcqN2jMT/K1HT2Wv25IKV
GpwR6cIuABYybhE4XZtNCFI9FU2ELvWwhau4x9SvZy3zExm46carV9+NmcR+WlBP
LdHjlTnoR1h+5qFjuSZeOZnp9dvuUfRmWhafh5Mxfq/az7Zg2HBYuvkNuk1DCPIP
oHtp0AZ182QRuzg087tuqlgtWXuDmgjqX0xsQtj9Hju/rsfwfI16U12jvSdy8Sqi
Ew+hmcTf2u+duxa87pOJi+W/q+vRISbxKAPjCPWfeLc2m6mhK/kVySHSDwvy0Djn
KyK5BacsGBFub0pMw8rL+oLwyvwuRZFx1lbr41bzmSVWcZc6Jzo/Cf63UnyN23tf
l8X9RpdOR+ER6fk8ko2oXZv87AMx1gxa8jq2JR2yyo4xSDx+8DYJ+vrr69v3lAYe
7Fp7jcWFng3hTus2cio1JXwS3FO5tQxVMj3rGaibIsAzpuW1CtaHZCsvC4ICI+kL
Og2xDAI7Bu8p/M+DNahNFBBn9hRMKt1VT1Wgie2jriW2yfTr1i2ewG39UJoJVJmr
vxIKc9u4VbMPqJpVnwAFfGSY7lHIs9lQu+bbCguBkY3shWh1JBD8iMGKTTrWwzFT
YYzVTxwEsGE2h4C/mWLeTmf027DIpQqi5IDQISuZ+9125yTPShcNl9/T2nwx/BFL
l057ww/3QApPszQcPWpPOfRqHOATXC32BlnGTAao7f3JgkOF3XG0Rpf8SVMMIJli
31KBHpb1lQ/x9wFretgmwUgOq71ZMZYS4qNbyb1V4ZUrZzPDP5VBuBFsJfpAkhyK
jyjBIU7xWswX0rRGFxTBuiy3Y9bYQmuP9om5uyR93b43BeC8AFqS5xUsNPsw5Tr8
OnyPq1537oCBbsO2dT9Imf5GJ23fnfANAHc/W1oKe87pt1PlyB9TdP+lq3mJIDiB
N66iWjce54GE7yfTCKnfRGqKTXTf8K9HHbMw7h9J68UZXBnJ5juj+ntN+fOiWrJF
Q2zG2dSkJU81NBZwYuDiFpFlFl9kEVVnwKapTOhrx4ZuZSB+12xStYzRWsvKhhHs
NcREh8x6nBZP3zdiakGt8tZIgZd7io+jIjeeell5nJtucNhzKRssBnSR8MF3/mfu
GCfU4zY/t3az0hxfE5gxMYq8AJDonHHegytpejX4LnpljzJ1RhGtNEPPdexIRTyf
9ATSvLi+794VCxxpztYzPCNo60FVxMJF8jhgfjVfSgJB/VB7IRRPtAKy0pwJSlWm
O+ltCGd4erR1lFlQYUk5xX2gFBdhKgCNpUFBJzeRQTO8xflIJ5Cd13IOk/QUGlF/
9NtgaqSgwALOewnvU1iEVYJemHjPiomh5MYVMHaGdT9+wAx0wN7dslRjrBsIUsKt
51LajoR05AWkpjoThx+SbgyaPz+l+UR3E/nX5Qcn+KYcRPwTMBV2cpkIaq0HExqs
G/ckr8DJ2gldtlZbjLfmjcFa0OU/fGi9JeINWNJeamZnn62Ftsyf7vceWfFE+oFI
ap+WdFE3mvHDcdm6TxDcPZjld7H2ogcREDlKRSyo8z7df8VIJzV7LZGNCwP/fosk
ah9VlErHoTIhtlW4XuuJECgm5UA7tGZAIsjYf1bJvQZbWJjSbj6gUOr73x/VauQe
rPlFBXzd+QMwjKIY23YaxJHCEYydTuXvT+sJu0AaiMwWP0h2lqPPe9TM+ZRGhdfr
8a38+oivtMfIvaBB+i9slJmy/4lHOSI87g7ouujPYpNwgmeQUMM5l3T5VC/GE+wY
MlQdD0oMUV2YiPgeVcsF4+QlCiBQx228ErFFY26JvUucIuPxWtC+F9mgPD22Ag50
lcY/TiR3ezJ1yZ2ou6sFYadjQXwuca0niYu48svmhlNRIOsiVurOcXlN7TDxf215
MtaU9NS3AzZWQbUvY4xxLocCysY1ZbYvXwSmh+h7NrAszqWP98GhmmB2c+j6ZrS1
0tEuyV60J+DS9NaHjaQmiwM2j5OfaRIT/xF1EEUj1vHY1PdUmmpyrRujnMD/pmhP
tME2EwzPZZFs/oTpUxdNIFv5/o+GRgrAxflAK1rhic1Kp41yo+WIZ+bcXoHD4Clf
14sNH+rQHdM1vrPJTRxI/bzpzTUn9tP0X1v1iG62JkZRNPzOuhxYUjaUxbBiZzaK
1IYHFRd8T3L3Cnapz7T3Of/QluMtFz/nkhITG1jKpkEKqtXQoh4QwvLrfZNn+ozQ
OdJhrU/qiR1aABT+WxzlTal0nySahPu3VI3m4GFaoaXDpAF9e4Kc49MidADaO7X6
4jWGdPFWzBlUYjJHLOjULG0c3yc1ZgL328QZb8BFVD9joUGMYzgbEOtfyjek+WLF
dOO/4nr1aCg4toaKspRXMd70RORX89XCmu7sLGYTmlSZ6X4Z/nTGqVWr8IQyuZL6
GViVDzYwHNGExWxqiaqR93kWPg/FaIPyc16nBuOlQzVX+nl4Q5HKGEZvRSsdpTzB
zKUlQpk/hSsZHQ68ytydKXA8zbx8Aq/c8YustSNTpvRLhO6VAS5zmu2kro1GBpOQ
X3p1wVrOrOUyg0vpI1k0NfqATGB+aLlxZf8N7vlEUKimY3fBDihEc+9/BWJlkmYp
jJsV+UliOtl9U7vK9K5r4kj2GCChzkXFIz4JjX39bKc2qHX7SsBU0Vs/daMSc4Wv
rbKOR4jMsY6QGJWe52Nj0FnUqnQc4XATy3j0+648HnqSeyK45WgsmxnwosrgP2bL
JTzB63DAIFK1Kr2G+uA41yqjDYgoNS5THPRG9h3tv8MhnHhxnLi5qju+A5Cuzu4B
XpP31hrOLe/GHXYCPRTXlDhNdrCowYaN4Uoa/TJkoM1tGT30hY0OqxevxnNI3Uvr
7GNN57B46XAKWuijcGLQ5WyeQytx6BKEL9Hs4tBvRMSm6BOFm/fGd6ZConqzKgcP
FdSFst1qYvk10U0GqhECMl4ZBwUzlZ+ig3w918RqKrBvm7UrwemvrdIgOD7J62YQ
92icGbToROMUlw7LJ5QEhHjxyks0R+fx1AXHqGkBPOjtkBph3opeZeUCcYnbFKb4
+esv+MLB1Wqd4/IU+7PuMaAow7fWxcLlN6PpfOQBNhFp+C/QY2aHVj1C/tdMDdIp
BEHOHaJIYCBhmw5o3bvml54Xx+hk4dQRqynUdQEjjQ30TWk+FlIC1nlNEPnR0zlr
gsOI7GxB9/C6NQMVElfWx0q3LDTKQRx7g/t1Q5Y0/c10dSySAffFuE8NSwxqu075
anVnffVOBeLNIbasd3BbRMCXoyMTxik7Ch9jbTyQdvw+i1QRyeHx4Keit0QztlTA
zUxMz3inVqC17IgYLJXeV6XJZsq14ZkoN2Q0oaXRqBcJ8dmEiljds7dpsrR2ZbEN
zVI0KI83SUPDL5fvt9ZnBUmYxR5cM5bbTXJ0oCJutfG97mJePQV9Zh8PjlAdTAMl
AqAYA6i1Qkefd1hQUJdTCs3D4GUHVeC4J1zGkJVrevorJjZQSTDCcNRNIrgBAKid
m+a2j93sTciZXQqkTLFYk4EGMCvJYjZcYNyag3rFdOHDnPW2JBc7iMXSQyD+8dZO
L4Bm0tEE7JFHw3u9ReON/pVlTm8kU6n5OT6lS8QNKY7WJaQIqtnLIGCcMIsvppyG
hLSI90ieDKF8zKfAo+o2flb9bazFAQM5/4CxXBxWPBx6Q5pGhHMFe6+KPWyYQtb0
JcZsFZd3nJZHHMgskl4J+/OnUeaJ+PXxEc+51qEnVYzGEvSsy1hwHZWqGCnS6tNZ
/RnOFNt3Isb41aAd+HWCCb3fQgaC71gL6r975YVryh+XDt0bCACunJHh5yoC2NWb
N3qKsfX8mLfnUs4kGHqtvzJCt5qvWHboInllR037JSP/aD8sCUBeKRPq/9hQvIC7
oLB+NlFuwjwCZ3SXAfWU3kKfRnG5/jeZfdCvAcwqKsbwB0G6q8hE0Byt1RXn5gKD
13tZHFs6QolH5IxU1EQZkfvS3Yk67mW60YrxJxYvHokMzgAf/US368vHdfwXQ6JX
tPUPdzBTNxg9Zyqa2QZRbOYJlrjJaXp6iGxxQPeDrJ0mBJBdQCapByqRJuC9ZeLR
9D3YP6ZK8QTNBRd8T88+6RCt8lsuUI87LGZox9EeuzKCMF3r+6MGEss+NYPbOHLt
91B9kd6Ie2l+8e1Zfd3I47HOVeBPHlbFlrHh50nnkB72xuodEciSSdrHLuQPgONI
PrHy0mvOdLAMMz0GA86GjaOfRxOX5TOl2GVFfEwLxBXcANPJ5E3WZg82FsJ3cyvw
K28xh65g0uy8pN7o74SA7ZW736ZS29Fj1PR250yARL9Vl/A/mCIEnCmmMXeImO3p
bGZZTz+6T9BuF9UYQeyANZ71Mpq+g/Ke2rREdncjJWWit+9XFeP/JYzoy2LPXyDN
qQdl75fuBGmuZpQnNPD0jHzIXV9Kp4TIkZtgJ8orqkVLNJEra7WkiK5spPRGWYOs
VoP/uyCa64VqacP+Au6kz4CSXetuyt/hBrJ2suvqmcjGT86g1ASI4uFK3MJ5jhIr
AeYGe+uUYUuFH1y+zTecak/cHkLIrZbYeKvT8JzAh3cFboDb8f6kfLb73iclUikK
YUoGLK4G8TFZNk1PZDaFWSGqEh8HcIZvA+UbQIqUGBGxlLqaIjhBn68pJNp5z/9O
yf0RwUWLD94xXiHI50YlPkRqoxCZdAgYWoMMWYYc9iwgMMYaVvWX4EyXvEOEDNmQ
isoZjJYfpQRiZp9aQJKmyUeGtgrM1VBXgALVN+ANCAKXeAYHBT9wtUkUSafNpZuJ
DDiaKHYpOPomVKQ0jZFEt/6Fp0oPG7/9Sfci1s7UfgWfpYaAejTev4emuGQUHov5
/VYttjuxb+U3XMYMWHw1FITSpFx+vKbV4coSmW7aaDXNLsOZ2G8k7q08ZQnNOGzU
eo08mxdkqgekvCHSk6D+kq2dg2wSyCtAajA1liwBj5l+7maXjtaIFwTMOW/emz41
ZoRm4Cg1YsgGYaqoKg7tDjae6D7kEDMKNvOsjZlBxoeJuN+YAjr5iuC2GWWg5RxK
/qkCKGdMac3oRFDi4WLCZmtEm5ELYKdxQVeHM2eWBha5kb68H3ewjbmOJw0NycUN
FkntCU5tCdozO9mtCx+1iCOeL6uWtSjI7J2CpG7cKfOcE6wPfl6eurXk459z8zI8
5MziOzwthU1JC0lXeCSIX5xnyPsx2EvyTRn5der1PAhJGqrTiDbYyq2dyToUR3Fv
vDiP6Zd2Db54nf5ly6xK9X64c0ozLJvfXmYoxq6E4Z4gIs5N04rN+TTPAc//4sVT
tajQ2XBwBgYTffX4lq9nropNe9Ds/ff7C5BRgwR4s826gHE82L6/O7KTdZ/8ZrTh
QFMUwfRJQdfsyUrrUoejSvMoTrm1z4Kyzo6jBQ32Z2g5zFgAuKVGOUZzw/88W2HM
SxIaN94KAxyeuRsLZjkSsQzLWte8BUbMy0s2tCCHrxaIc0B4NQciLCXBh0oV7sC3
RUOvoK5SNjk2wMoVGYVN+nokC6chFZv3v1JUsWPtxrKiu+JalvTdmEYyIB/jCvR/
qWaHU5T1GjjjFC7jyCAa3clhqzJaYX/9+2n2MKxeNl6pOc7wvkF0HEEeYF2tgfaI
+vvsOXMIMConRP9R8GnuNUBF7zkZ3VSOxruHmDWLNHc9cD1Ncmhh4+B2AicXrCbg
k5r6gyeVCif7Q3CaArpw5kpcL3j4KbjKrRpE3p4m2cbD3c0hVTP3OxO7zDkZn8Gc
6R3JWeBaso018QVl7lGn252Wpfgfx0W5K2otQrcegXct84SHZ1MyzmOKb86CPo6w
EPx24GLF7mwOqGuZ5ng9RmmX2lbg+n/SQp4n5NSz9nnByAcu6gNWllW2/CVMlOty
ueWhXSXXV/bjDKW3H62oC5ooj6ztJG6ulyRe5fq+HEvI2uL09Sic33rwRsS4IWLJ
uLEZ0TZpS80pfKm/O2/iV+me+HiXId50WYie3XkxFumbjIDg9ITD8aETrJbjTRSi
l6IAx9dRKsK4EJCn2Z1wmGKlsPhxcbkgYM232NpLumdBobJUsPmVpUYkXBlpq18L
sy/7j+KxBbkJ/up1ERAB6QOxJpgMUPGcnav3PvxvACyJfuMmGuQ/LkiFBpvIf31I
m9eBYxoJuMvAyvAC6Dgo7KFMvpOvwptwOJvwz8QqvZkE1Cyua/7hZ6yHW9UjmVsj
ETVXdKq//Hr5unzqcsNOhqmxNJ/dLD+jKDaf2IsLPIEb5wrkK0tofgDH5OH4F7PS
OAybTz5JLkicAcUDBIvdsWy9CJvQgDD9MJK6gPMDem2KFfCzmrQ2iNQyODK6gCDx
dtS1m445Z7No9hNxLAmUts7p9T+zmsa6jMoQkOdMYoTTN6QdmKSEGs6RLVCfMTf0
EJtiGVG4AZyQI2PdPJ80xKo8ZKkK/he+6PrIyCziX6FE7LuSXVUcqOKYH91QHwMW
qV5d75CdD1+YsPnXgPfizxS/B7Av12p0NL3UGfH+8C+6NjdnNzsMYOIr/IO3I0A6
5Nq7MPoYJzj4gsTh4f0FNleCFTz5bKXq7m+z/qeA0FrrwPyQR1Gn3FKD3mJ5H0Cd
kZbi4KSZlqLvOFrxJLzWitSHbXe9et9+I4lMpDYfeUPi1pFiC6haLVbqoER8StTo
7hyfHw0nb2CSiOIUjZte9JgjajgFIa8YhrQAGwFVM61yvLnx0l04q/u76G0wYjC4
taFXSm5DqiX5RDfuKJKCbALlNIq+jpyXOdpKrYtPnDOwtPKaFUxcg9+imqZCI1jY
u8AIUwjkDtr5R6yjiJBRSVXv7q+Vjfr2uHTgA94r57k0gc2bseDjdl+cbW3ZPMHJ
QuXaDuh8Ha8VHzmLcQTOjL9/vprjEhaGuMbhuxtUSEeKjI5Miyx5kfz9iivKVXJn
M5XthBLbk9qIVQF3SOMnTmPAsFaTiTxqm05sqq2DbERCZzIA7KJqyzqwjkt4Zz1H
fOryD1EcCwqUpL+qHZrPZNLufngZvnUHDo++qfZYoQ7Ge7/fmK7fUUpeggXK+2pC
3pgWscTolaamNf3KEDBWxXbvvZKiGXWjeBgwvr8pvewiQyNANJQh9Sw021yO6ADl
BNGacIwXD63qMlhUIzI7YRdVAFztL7/bsgq6GAbA9EmvlFNSetF1//WiTIw0Q8I0
jfUk41F46Np8CZPW0KgiU7bsOmgu8TsH0hFNamh2uKz1aT4HiTvn7a/LZGNOE8sj
K/PVfEtnC+NqcsTHZhm5EUg7dGuZwtu4EzwXgsJs5kYLodevbPRvhZvAvxeJqmVQ
+iQo/xnsgG/j576Tuus2cx4I5VQdeyRC0aFocmYtN7SPtPyCyC6502TuzT1BkD2X
8uZEBXm0Jd0holan/Yb8uH9rfGygbZDvZzykHIg06/t4GR9To7S/tcVuTxJzfMrb
nFN/bA0PPqST+a53tETZvE/0o7HRDyAzyGHhZusEOVE4fumDrhfwTFjmoOq7vj4z
MHeXTzGJOQLrr+BS/TDwSpYb9nGxQQQyx7fFK5hsXiOFcHaJuZpJDBQRPZc7Px/B
XNy0i4HB1bpkG3VfN4ZkRVU+DyU1MjzliQb70ee0iaiSqXznUW4DdNV6gcPPGgMs
asvAA2TFgUuyzgyee+bqiO/vSAueejDlP//DZQJ5T6HzGtidWJ6KOu/Wxtsc0yzX
MkK2rFdGGzlB9Sp4IEYULt7ZMGQplGoP5GagUm4yz1GP9B6MYv+HW4I388J0R9M1
K/h6KRfbVRHv1U0XIsw9+LlMMuUz/DuU+p8IohDOn1aTmMw7lUnRmdrW/BtbKtEJ
hBBS4lFFvMJKAsdM5DH1RXHbXdgFr0kcGJi3WKBkdrrcdb/3WKcud8P1BdQPoJ24
M+J+zl2Ijn3TemZGzT4TqwmNBfE5MkYLxUYY3UJ51VMRaV0eVP2DdCi0BF0Dhkhk
LbQZwGiThn6vaqo9KYou/CDc+0kGbdUOkhTN8nqppRmnoOXvqUENnBy/Y0DnMiDS
SEAdBj9M9LxoDQEMwCPUbjsRtwz/+uVxfO07JMeJhwm4EGJL2JJsEkMB0JceRDNV
Khk0AenyR/HsCdvw+usQ8MxrkxUYrdtqgM/O+4Is1oj2JEFYbqogIzUMvc/pj4GS
BTjUo6UdiN9hu2io1nMgai/ZjaO6rkvAtgIxqUDHmriU136Yvp0Iy8nSn2czQ890
l6CwvYGz/mflXG5wG8cejjFXLJoFYCOAldy846PCCUSxyaOHlOFF7yjaci7KqDD7
6Go4xxRYPEOfvdEfRINDRD+QMSm1IJERNzyq5uVpzf1tJpLmFcKFP7pmpp2867Bu
gZR0ZqOW2ENBt+Pym0IvJOKhP77yW8fvB0ZEDePQ6n74R0zJPj0RS/wvIXVRd12x
Cb3Zhjl6hVfAFi4AX/pKs4czHPEiuxG32vi92lAKjVps3mYJwDP1WPX/bLyDnOGf
vHpBw8ETHZHjYDn81pD0KVjB4ykNIpfGJHnA2L0F2jvkusP13ccxAwswQmYdf7QB
UQRer/cv/mK1H4GmmIRWx5HP42OHVjznbvFfRsPp8Pj9jxucbuCJSj05ojk7yGVb
Omcxp+Kbx7AYDaGj2IoUsZ+DqbhFI60Glq+lJoa8fYCNcI1t7dsN9vjkhoW8sZGT
QXvUVbpivKPw14Fanlc62wSwKIY7c8moqvwRCnDr/nBT0tl/A8uVv+W5AQCWBu0b
okf7ZCWleKPQ9QS+i/jYqI8FnfTCXy0e7i6TRwTosJ1TYOWQRuzjj9qgYAmECabO
8yXnN3gB7P0Mi7VcP4Fwp7O/6KKUmGetiC0CP3kBjmtBe12iNN69ZyWy0RY2DGM3
FKxAzQ58mfAHVcyeJykCfSdiUm9dvn5QwJfdefRRlU3wA8zc31RNchkPhzTmbo+3
+PBMGoSClXT1mqtwDERdLv3yYNXN8q6ufTx+XWAJFzT9qonFAEDlaFKvBTT+2CtK
eJm8u8aAgmFdtVkPosJnVcU0fWKMrNDE3KQT/baSGSYPmPFuQkNwXeyG1E57bdfc
gr0xDR6kdhKgRZfOudN8Fv1FSlfrr9K5maas7zv3Ci4NDbMcDyxSclKFy+YHEEpN
VCVi9L0wbmXnXcp+WxZWh/xkCIuphPsGKJHJRXwh0MDKA+addc609EkB6h4FM4wg
wWpwBK6dxD+rku3D8dR3tqBPnqv7uAe8PZjSlLQLQe3gD+iEwKBMTQBi5EcIjk/X
27GyZ2J5+7vY5qWedxqrp0sCJCAqEudjuDFBSOm2tVjOEM4SkMHeAvjatz8Updpb
Us/w5365b4tnddasgYXYwFq6MAE0IybQ7yzrDYt2V7TaKzJ2wkXsRzG+14nkrIn5
K3c8C9LjHkHKy9E/tKGR+6VybrdZBeoqAEmUy7X7fng1anBuO5dnsFkCjCpmNOC3
eCOzeIX7Z5hD/a0ZP7Xgse3KYgrUTyz9nEuDkOboogyiJ9CA1cUXq+XSEmCTvY8u
SbapY/T7iQnpC26yGzlB9Rc6JEhOs9CiebkSDSy2gVYLAY9OEBk3LOymdriykuot
h6NZRXMqz7Xl3hkkkZ+i/lhkfgHawd1aDF/HsZUT2ALGIZgjgpiGs+cq+hmYxrq5
3fIyWxe5dKP1WCD6/leNNjSFEukVQgqMgAG7B7ZiMAPVjQrK4jORT3MhBkqd2u/J
9qCLbtWhX9djFWNS4UUJ0uLc/xeZRCanKWfCamYP5NRoKwCF7SPFHy/zHl2m//e/
JAEtuvaa44rBfqIEvw1gnSNuRBzfGw7ZKuWlS66SNJ17FJ+I3Jrpdy9JP1fG4hSV
L3UiGHDWMdaH0k+8NCoAKDNJcTVb0L8IpXsdJ0LTRDGrjA4T007AeDdU+UB5DQHp
AC2qxc3AllCHUCmIP0eHTwK/3o1xqa8b2pLYt5UIOiLgq3PBBEfJANK4iWOXEmgE
ZRt/523evdhMCyE4hQVhzssXG2LJGRp51IxK1RmrOo6gUDIBUQyxaIoYeAA6Wawa
PEM+RsJD5rRPspKtw7/t5edx3ZtiNvPaKii7QXxVPqdgPUrUkru+kEXQwVLLUXDt
j6YD643q9mx5HBG0qYbpohdE4EHV9uKxULxEQwyBob/XzXOAyD7ycsZhBZz2MyTz
a4zxBUhAiwwp2loy8LIVmZaQBm82T/kmoWbPpkXPEi2IYeapeuzZYK4szUPfvDeC
DfwaDxStlm+5uFkLQA4HwXjsnHaK5HrbHTQUAGKMQ5B9bfL2167HReqEnb7dnKRJ
UhX8/JgONdUpphI1CncddeevJW7bcYINjWTGYAW+nmvkE1EgsuPX1Re7DVLudk+t
XW4p5honGlEAA02Q2Yeu9eALwtopj2kzAE+arypfkYgAK8GbTfr/yk27xK3eSkZ7
ji3fUD8TsmLOZ0lH8rEIQXsUJ8YPeNAYEe861BGC4Q8l6KNBiqDiB6DrmeZwcpmQ
koAzyUsHRVuahFhQKudIfq3uBhje2K4Fs2iUK2ngpLiU+WV7ZJmLtdmu7whvlDdV
vayzFGXZeVqt7NnknNhx76y+eRuqm0hQ26d5SSR45Zy6bSJt/HggXu8i6afbeXyP
e7CEFlTk4Omv/JLJV4EhvE+/ralZqpPPB1Ju9pQ94QhV4HuaDi8dz0XxMFmvVnWP
Dib5roEVjSpyC9lVIu6DXzJo2V2jxp18E3FSSmC4h8uJT+xhsqxj17aeXDJKWEO1
sGomnafr0bSciJo9PWrgqri3xlNKDSLuZ5xqMPtuR4lWREtAE6RJOQoArhGieV3C
SckEa1yK6YZm0YVsquX4MXMw802/O6/tnpylh2630BZMJBw4bacyudk3/NmfVAQM
gfhrFPwf8GiFJp6NeCr89e97yFmP7BenDOhr1NgidhbE+zvASRGdynd08+HKsoRS
xT8P1fbK/RYI6wotaAU0C9wPf79w/ZYPlP7+KptVdgvlvJRvUNgJY9hHySkoEWjd
52hFWjfW6pTR6A86D7ACup+APhWYGFptNEXZuvI3KB60BqjBzUD3D+k44S0SJYht
T69MSLhTHz7dcGrN+T1xIIya7GqP/D+4dKe6gZVLhYa5S6Z9Fn7j5tZ0mD3BcpK0
Ib8RamPzGPr4tfMb7T6UQiUU3fe1X9HF9LisM4NPERrmZt/7AXmq3OJuV+Fwr/8S
6cMKvAOVupqGde47IE8JuxmhiZCar18DKA9mSFzBXge+IshQG+/efJ5aMxHzjFQY
hJvWrcmILy4UCTyMQlq1ltzuPe0P8dQx0F+h0VCxQoy4fjmOrA/TRufFoN1i5Ls+
tiMvuWZ5itQ0X5+713Zfjiq5xCszBQd6lSGDlDJkPHfQQnvR7Y2TjVvs767sJdWM
xG2GvOlpCSpoeZqzzQaj+tUYFPUeFqW2Tu0I5cs9yXGv/E1HOsenb06YuBhlfOx1
r+dsrfmo81H25/oVEw03hIj+uPDDXHh2hGPDEzWyV38zu0KKigzZqX4s+CjVbHjH
HsbWO+GNErWswvCRkhiRasxA0nJa2MnufwcF2NSLVtl2ZbqCBI6P76ohR0fxnXNi
0Wf6VruAVQzaUADWY4IjlQ7QkveDN9mWadS+eg4SQ6PT/YvwVIt+PHOw/Xk2APvx
zUy1OhzJzyNTidEYHrJ7xmU+awre+L3ACj6RaMcewwk/wet94fmDUNe9nMB5kLSH
Jn2iaNPoNBCxSqrsFPvrgOCDMM7BDk3nL+Gk1ETT6B/mUN2xyhsxbiKkITfxbIgQ
qcsOPcCeU36vZGDmY3NHUnzhqcgytVBQ4anBD9Bf5ec+uYrN7AFjw7aoGvq5zC29
/45lWILlQhZTY/2rzKW3OgrZhDSSJXYi1mDODQVy2N0xiQP0u54k3wgYsFpASfK1
j8l0D0pI6Hfluv2GnghxSWGdwOZKUZO3zn6Dn2VOBZdkEQZcKMmzZ3/VyJYRrtZm
6/Tz6kpLQ/zZIyOHJagfHeFKXBFeO/SgWmyAFwru83lDPKXd2Klea4HIXhCaVkUo
eTGS9yHxcQnnZJWt5RpW2sqIBEMf3fdnNjpvowxJUjv1nKM0GSIcSO+Gl2ua8rs9
GrvO3cjQDAlPo9cpKJJrlgzJsfGSMmsR8iu0gaBi1WKpiVyAkekzXIx3N+VFzfIX
9WAgLYZsGUVYEcIzZlsEh30LQvRLKxrzFlWTtG+pVrppbJCaTM9bbGAzo9TkA+jt
ISh3wwCUKLvSF0NL7wy3SXmSE9m2EUW+tMHwx7bKh+Itk67rhUto5R1ieAA5q1kz
FsNDz1pRJoVDP3FhC2Hwm/GT/Sj2x1Td+jYZvvXta24NZHJ0VwaNhBW9XiaJ1SZ7
IUn4tloljpyivXQhXPu30KMlRnR2TqDf/S/ZJ0sEiGg5NdiSKby8mByU4VJxzCfB
gh81Qc3s7haxyIk0izi7sCOnbPAX5K/VeASjzILLiX7pHG6D14/ctOWjGU29kOXE
EFkjNOLwxAOXAvyNyey0NY/dQ7fj3L5k6+n8Zm+MP2wMj5ygw5U0W2P3yAO0UAG1
zl7Qk55foNNagUX7iVBNcxAtAVpozjIvqeM5gii8HWO/McdvGC0BUxYFmdwq8Fsx
mSOQfKSLdGH8xXekL5oGvEQfu1prWp/w9Le3IQbiGjkiipmfpokRdwl8C9sHyETS
5WBVXfwKgtUfXsr/qmnBBslDFMiy8qKC8O0e0t8YYNeNhdF62zYhRv4MlHsys04i
xyB84QoKDrDITVxzty3AAqnf/8RtKqMcY4OcpO4NiVleHIqwg88O2hOe08uxkBlU
lgZHNDpEszuzqL2M9IRr3bXYZVRlPAJ+PgmTjloeeYsgOzZ5+uzwi8fMVP6T2jth
AU7cOqEb/Ir0+dRcKKWYFJTVGYD7Kfu2mI7HBM59J7TgTvkdQi6xqX3v9OAcovdf
2H6E8kKBcCRPvHImJn2hC9CdM1C34yrpTdOwu7E+KSroVrCKp72VMjKi/EEWS+JQ
10aI75M4f3y/xmZObQ30q/VCp1/NF29VbIjCWS+sLClXE1U7LYSWrzsi/k48rnXa
OGhsX5lEbH2wKElsfnVj6ZXtds4yLhbv15O+NN1C6V4OAw/PlN+6xhUEQ+gZ99Ju
BTR1lKf6NJsyqWeDMqQj7QJpNJi2kprz+q4gI7TKKz/biY/+Thb1Oox9kTNYuu0v
+0ddTqdEHkOmbluxEzcg/Y9JGRLdo2QA00DNWs3GJIAQKZkMSOLYTuh826EoiyVc
ANHMXpPKnp10P9PxDSIxguUW0WEMfu7AbA9cAzGMgvlzP+y1NOiRYtpisGY74Qv4
6AD/t22ZY5uqe+Z4JJbrPQrM9iuz023BdfxzMTwknyvqqFvImxCl5WOLoeEv6aLt
nRdYKD6zMaQE4HzESdk+JSE9ROIP9J/sR3GmY1xd8N+/N3c4AYqeVR9mBKJF6I+T
kQvxPrPF3s6kwanWj1cGUwVZkhryOGt+z+GuNcL2MVe1nji8RQXj1H+EAEmo2gey
FyUpCvrmfQTjbl6iyOHjifHUuJriDQrXbUkBZe0VCYb2oJVMuzeMkYTJRMQshTMz
We+DWdzl735ZyStFKpcuR7NvrIAoPVMuWgJHVTJevtg8XZq+75auK9D3ny7D3BST
jDvha4I8GYdCiBln8S1GVAAnV6yDdfpSgAr2N8tGQ3/cjwsjCoynULoB7yVMcmdz
JBhZFQhKfc7RvwUZPq3fTYmiuRVCFp7XLuZsRuz2keq4Obt2Mul8reQuMtVdQb4e
wl5AFFmP6/PX9qwUA7vRxyDR78st/xYtK1sT1QFWi+0BzI05LeCNS9+to/Vg3Qox
SBId2Ni8FpeoFciqdb/ICqPnD3D3XDNmOpPGMuauJma9WS1/YyCKWsqnvAVm6Vhq
kfCdS3b3DXWktniD6eUhQU3RTaRYFzrFUVxd5GFWkiaCU6Hw2+EV0ox9/H8M3qLx
qOFzroZQegy3ZaH3WHtrtCnY3c3qe24bAeXHxzrk1tLfAU1QT2JN5JIMwZVeCk55
t4KlZGPCBhNDOXX/6tkQqz4cDRYlyPDwH8FTsu8jN8FJeMq2kaDz0cVJ7U99QMYQ
3lXfGsvVRRL4pRn8s2DDz4gQ5SsrT1ezKhoUbCosXsnVOt/IxgShdmFtZqivf5UG
OblTOf2gchY3BwURzv66cpJJ3ds1TCHMi0zIcp0U5azdUecfMFQJRvtXHdM9qSm+
Dsqngmel6W/aFlDb0QEnybC7JqKpMrnUi+l38z1hVDfMVHSWNR9pDrZiy2ltOe4q
/0/ZcbbLVQD/wwcZ4pXn25CZyC7J8c9LcdGoWl+i1ppP89drK7BHfbiouaMx5qEv
5z3cdTcUy0bGNTJi60sNsRGgS7yxUKHd3p9ibdjgBJUrh2F6dhZKgaTFRbupPs4Q
r6sIl68VYZywjmHnmyKyKIpF3K2D2IF/xu3L5coH8Jp782JRqWlp1v8Pwb9UhUFX
kabt7PL3UiBzBofC290qB+j/Ye7xcXWLv4qP7RK0hSc54rhGytTQMRAMrOkSMgiI
5UgKzn31NitFhwYE0Qu2/RbAQS0wPCTBZR5YgLO7D7yVI//ow48IAlS0Z49DSkx1
8T+Wn41GdeyM4J9sL6Oawhnwqx5ad1eZ6XzusnU+kH+UuQmr5pID5XN/W6JJOlpw
YJdWW25W6jhP6YowOavzdoM0yc6Veci9wNXbshqSX1f/5I72LzsspqZ0zIYw8X5y
lFefZaov+pCC0Sr2Q2JzpSYEsTTI3rIuk2cdy6Ysd3eulhVvi1BLpnOGjQIYkvH3
P7QCigFHRHV5VRwAmJ2JTIJf36EvwNJaPCuIxcORiftt5MmvutJwqOAllljzMt5v
Y2mJEzgmjyBR5v3iGsvnu5YWspaF7QNB0rMZ5t+zVQDZgEaEGJRu0P2+7YidICG5
d/OKNkKedQ8YzH+Ms54FRqKzF7aZiOf01kdQAYsHtNnbT7zrFYEqsVDKbzBN/Ypd
FOStHOf/SSLLHNpA+9PRzqz0+cwzQD6Vb2F9QTRsUngx1qdyedJHBwKe3/bOjMMY
LpsuKYyv7mTc3zoTelY6Mdm3jcuMvbueTQLTqSBB7XeGhYh4EOGsujbHMmtEVkiX
cQkLUPj1RWXfAGliq96J3wxP8C+OrYkZrHRUInf1lApgrwiyylf395GofkIfaESw
1JlB31DdJYomHTJVd9AdLtvuCrJad3orTigJd368wADCcByVBzhfMaMw32fkn952
XO4Z/K9wFVw8cSy891C+yIZSgI94J3GMtlbCt48Gjy1VuehmqekZ+n2oxV4e5lMh
QPESxlcCwvDKGXKmas5k88/7bWi3wT2xN8Qt68fr/tohVzxSFCfpw5Cqz5cUuQoC
KTu4/3h9UFDTN00iCSCYMoJ3EsB8Z2UuRLdB+/8kV6PTIbI4gtFid1j6D7BOLBcf
qu/ZOPRCEnbtNcv4PQxAvcFsNljxLgPZzvhlp3EDkbidRqhhIwI7Zz+EXAcgj5yZ
pZmhBtCISxKS+8LiysOgFo0j1VOTlScTobmWRfDjdsNZTMjnl2JIww5dQQhwKpeP
KAfGSnhNXOrYlVzRLYdmYRdnVv334QWBKCrkq8ylYS75zIEHiAPudN7gIkVoCiws
D8hMGEAeaDKGMYUDT+Wr6RbxNdz3Wq+XykKmGtNPHfX2FHwkPIDiiyctZoq8RfIV
KjWPezrHiehnhdqbOKOs8h3LUBCOVlu4tMsP1XGvQ+FNVyFyrPz/WddL47b30F19
VR39r7gpJXzTY5Vm4/WfAXUv+0NcJBYo1z10Psz/1oHmRK7ryWQQ5cWD6LxzQjWF
yTRNNkXIrAjf1cYQVjXLmb9EfKUYlCNRtKxspTggvTLgNPq2zSbOsZwWHKWjUeGj
J+7QZoPq3/TcdjlOsGUgpr6wJtZhVDZZ2l5++VPD9was1szF3vLAQVB0W+DesLrO
5DF6OoR4MQCRqZP1UHIytyeuMgDvPm819Vr4chNIpTqxqdMIhC8tImAFzmtWpgz1
NYCZtBg3kCVgpBECJR+yeKVjbqCL+Icyav5IqYzNrg1L1tWkW/ALiUd6f6IuTsuG
va+9TGr3K41SiWZbQCoxA2zp/zsgppdXhY9YOlidnyV/5tYH9bjJQEkWnbhDIMaw
kOXMJY7QRYvXWmAqT2VlMKa7le95btcgFl2bJj4lalXO2KnBulm0NQ8c9vmieAx9
zNOv7tW1U/mbT/4cSkt6/cnHymsvtId4GTulEpwqObsyc6lceVRPk8BlLk+H6mWv
LXRFjwwiObzxqEqpxyhg6uG68RZ8QtcDZo5EV6s5fWdL3LN/hDG5WFMGqW/QJlda
WespAt41KXUfJdIsEPOtkR55UDtDSksjn7scOdKR29QdczxcIGflUzn7O28ysAFj
CXVbMb5oXhMt5B9dbxUHzfumspafBRFYt6MK32VJgXl61MJNSQzb6naTbsItnxv4
+awAkoewE2RS9AVxZIsg4UJW2cWiF+dGrjDQ8WXqZXH0bEMqeqzrZlM/LJFEA0bZ
JkUnYKMhQBm+jELt/dXHbuytVEZTiQUKGhoRulwLoIH7YphO0wZsf7+aylqejWsj
YWKW4Mj7dMK2KnemMg1bmctAN0WeqxtEPfGXGIHi+trEovG5O31Elbv2CRnKqLTp
InPx8b7hutE2lJD6ALsnlf+VSztkZx5YQ4JFdaIZuwQBAn0ZoKx6myzq8/wGCk7q
IFkOEDj58G5IQRKDD3fe2coLLruUwLLv3RSdo9R2uq6y7YJzx2r6SlQEZlDRBzaW
12vzSLP0FBjpU/65qwYH6yEo3ukyT5qY+V9Lgqwes4Chj8XJlnNVt0fErBA3a2pd
ZWM4n47meF0nj3s3MkiMg7HwMih/lBo/29Aq5mBxLdF/dpA5xpH1+77iqwvF5TYi
5VKOlJLhCaG8HU70Tv0I39vI6RN1V8SrV2BKkmaecTj8c4RpUVtLVXTyzy0eeOCh
oaX/3f23FdM4OpcIFrjHn/dXH3BBRK2+Fn46TCC4N755yWbwOWyf7sjXvu5VXIOs
JtC4d+Sgbjk1Uir40PPuLj5Ti3bNwsJWDBEVvEAjZh/fHXIOzqM/t1lHTppxm5qa
r4JL7C7zESKPaJFT8fQkOOXKMiZxqxIiVU1bb8NO7t+I0YmgYDt5WTsJesqGbTT1
vcscW0zrweWSQo8KbcTc2SQlMYwWW0Pm7X/tysVcDF23DeBkVKOdOZ/GsMrPbrQ2
vpeNyljFeVo/2d8wk55d0zA21msfn4PDsfvBn8AY1AWdeCjmjoTwKZmTtt7sOzxY
3ByD0P5+/Z0zF/6mItEAf52eBRW5/x7RVA2kGbOVSNhWp7hL40QDTNsWnE+TmDd+
F9SNuK7zl+T7ijPtaH/kElBVUOp1UnO9rvEle6BH4bLTNmowPekDd+bb/uYXBJuI
zYTD2pWKHHuJjmRt2QBQY2aUYCpuRlPlUbO1jjVy34ttJ6rnHkfKPWuR5CG1cOwD
ysWhEEwD1p0l/7IuUkQ2ZLggDmGB2eFfI7mgO/TVnWcu4/4v02q9c8Bnql9z+Ebe
1Ixheb0qP6PyEqGZeIt6ou2F2NdCrBNDp7vv3UbkIEF/mHNivJhtjfn/WSXu4D8V
qHRHvqfreWeIDLzByyBKkpogiTJDEktSK/EYLQn6gaB5YnxlmRG8Cb6YlbK5nTnR
naWzImboJrbNGcRmLQZDUDgmMDtXR7P6uFJ9JLwvq19+epbvPtOsxwpcxG/rrs9c
QQaLyZKR2gal4V7r2Vg/mGnVo60BoagsxyxzvgUnCIH7QRWFa6PQ0Lbo2rbFvdKa
QgFtQf0ZYE5EnljlIxhUQh1kcuxMlzjnXlgednepNShu02IQKsz5yyMnIhdx+yrq
PXmzez/MOkf3ngp/ayjusdbpEg1HNmM9amiwl97ZWoVssgzD6aEHgxiCN5l3JYL7
JoA4/FnGv1PUU6a2+2RQRNTWUPoVUPFiLOfENhHV63SmKW7A1pYZxPNNsFvSqH53
xQu2n/hcLkdoyi1HH+y1x3neGPePgWCpHJSmJ00Yvza9c3sZJn8vbQ4a6zYNSaO3
xI5aWlv1DjJRzYWzhMrDmAUP8x/3T/Ooc0IU3UJWghhmFQT5NhFNjTOK+NCSM3r+
QxkcrgPIN8XohYvZO4cwLXxninj0h1TMqRP0cBEcmLzS8VXs6+5eDtir18dkOvnw
JNglcJvgL9Ts69KPUf1WjRvav+4Llqfxuuf3qIFvY5iewXRhYrdfGjz8mFB5+e8D
XPDZgYHi1V1AjwIxlj8iNY1C9xPboTDHBNaDFCbUykW6d/FcKIE1/tL0jpI/qAqZ
6yMPTlE4CKInGC96s7O6iwL9AebxHaDu+V9uF0/oG0SlGjhcbNJsH/j25WzZv2mI
uebWW4+BZNqx1yFfQaMSPb8gkTL36C96NnQOK9OQ6lb+zfRkHjHfhlarNGE9nqDA
jdXE+7bIVRVbLXYKQgYjF46nYJh8Vm3/lpwAdc9M2DZ7z/Oi+BaIB/thaYD7TlB2
C6J4Osf+P7lHJGciq7pB8w/VGD1xCi2ByJVmv0FIlJo4yXrD70fbmwcpVQRKGY54
aefG7k3LCq7d2N2AZmvSqtCIVU3/Fdz6okwQ+Si+3l0vyQKdsPR+V9fUyXInnDka
lqhKRP+tRv26ls5u2wleslJnzmXbJsrt5QdMYropEZmtkiKQ3fzXa8MJky8KXh4L
Jgu4HmsjnuHjnEPeozDyyLPM/4Jgov4xUJIQ1FpHtb26qVXpjo013yV94yxD9gww
7Lj7SRac6bqG6I1BslIceH/SU0YoE+w+FuKfhasKKBSiZdyKNYEvLjW8D3OF2XEA
3/vqSZkqjjuNBlWO8O5qWFp/acMD3MHH23mq/g1ZIGqDs2K4fFM7gmlmMKOUwts1
/6MWDauQ1l99tozvODUCeLTXvUYc//FX0nBCjlbKPXq8Zj/TbhCrUk4aPp5KcJqM
gtKPE0nxAUDlK3f74qaM3UGpXPRvsEmX4eUrUqCL7kQPcjaDQAs26gE+HA9Db+qN
RcLeGkrFZMvv36bp/8MMC9mAi7gXMo7erie8edPqIb4C1NgpD3PSZpFw2DPP2PMI
ZbUMdVZGPw22HQ8cfFD5ij38XgOi5sqqzAualbf24Z189VOMk7+U/PMcadcMb1kK
U/gh/xeWeWF6vsW9mEAuAH0Q+KsUnCdIL3vlPmvJBk0cAdfWWX38tvs4fVFDZupP
bnV6XuPtD5+IroGJ8XBasT7MXBJqk5FD37luM3wzvZ39mWaZMFVbMzuarRMAkpgN
2hBcjfNRQsoreGhEJUnMYLx7SpqLv04/lIeTZqqXguVdDbG1yhyHoka0yCKnmVyW
YKX2sxEQX9Q8zNtkXLfkSWEte0nKrkJ4fehR5H/XPTD3EXHo4xOFY3aU5IBwnXCj
A6Nw03IjespxX/fIW6ArMFhSrqGlMD/Es7r3ktOqLo2R82ef3cQwHNkjHtcbxn1z
wwNHgYiQcAhc+lCHH2br+Gf7R04eCrJbReRdOVlhjSb6aZ8e6shXhOv6fIF+gOxx
RDhbGpe+Rwx+pAm5ZrMDqOlNRw2CSEO5ZRCUJTb9pbSInzVqHi9+nyUSL1L7xHGc
wXAEOEYGqUfPPSDXe6Tng47CyBsNgrerphhPVUedFLiiL/ZW83XfidFZpyMoPHZT
ZyemjgVWIilPd8hXOX1dC70Va6e/Y16qxAdwjDOhbaYXeLA6f275YRwWlYT1fke8
tsjhIXtKwVO0uDMimzP+y5yL5NFzQs6OWSK3iecWrbZWhq2ra7k/PqfelupAOXvn
V4gyWxq9ooLbZvVqZimQYy15XOE5QDo7OA5TqTxKH2i0JSbU7uNZIQSJa/J4WuNw
HwGKbfDnAkVe1Ci98RoCa/0LM6aSmk5ki+wFJzLi9mWRmXFVwBQC9a6w77mu6J7u
n07DmAjd9qNhNPfawe5PqddDyMuDZknyBqBAmc27i9nF+gQoZ1igZabKVjLsQ7AQ
8Jo0fqkmw6F6p6Hq56CjtHPzptyFqN2IKo42+/7+T5av5IaA9P2NWQ1whxIS75U8
jFVDBhoDuXIQ4BOYw/eciWot0cPSZ3gtoeYiZ8pOiSS4mXLCYL14SBzQPNhNz16N
19f/q4HVtXOjMR0IWLQEMLIYfGCLAcL/hKMFjhwtY5E/txcgadLP2SwCAdYjzdL1
WFsPWBiPxDMNNoiIGurePy4u5pz2UA2vIXDgGMGEBtp84cuaVbZXA8O4aaufyA6u
H90vSFG87bMHq+QrA7Ft64xxrE6oY3R5C66ln5XeoLFMizVtopsudJN6tXKlq6yl
XnGQyIk08Gjb5z4xjQUBGxKsipCrin7r9L11W52rUDkld/Aw/iNYfxSUPMw6FuIj
cGyAa8RBQsNnBHyWo54Lk19SMeDBXy3MlPlZIG6T/ou+CYs1oR6e752ky4g5fPmd
MHuYXVvGrslNwu8QVgzDbjGi0Ot3oWbVmZ2nR8pH5GO9fxKROy+mXuYVemCbIR0l
Mu9TAMoixNtEZ7J+XlT9IfKt3rSKs1igbXLhTm8IAGTpZF1jDnmNhDoN6wPtq9Uf
TaJo1Pv8T4OrCyhZMdNQIWRT9xs34JTA2JvGFMx0bT/gvWXkIV/7NohDCAR7OctO
+/8va9Y6+zrPAcxfdQmnCCw4kkM9NmSKOXeBStalL0GfX83ghzXg/GVqlP8GdrUE
/5x42y/r4G/wpxqBtJTVhi7gjIheTtMJvfo+zsFb2F4cWDY76D8+kjZtVt7kOW/V
Ygyq0SpbbYIr0tRGYsrKoa/wrNBHG7IKVj9Smmhrfvbtaw3vy6t2Pf2o7zJ3fh+f
aNTZ/WpCR8mZsSnzbBExTksc759atTwKFjGRBJpQsOT7BsSrISA5kLzwpSgwOXYo
dhCSbnHHy0kYAI1SVp0RSx17YSfoHvE3T8lolTNL5wu32A7mc2tCz4oAsjMxH/im
xwmYGmkPA+thY3JrwlJ4YoUes2NeHWaiWGB/goRFgDvPPKlYUXi7CldRr9E1YZ8I
Cwm3bDjWxwsC4flizPlviH6LDB352uRu0G+I3VmS1nibW9hKOeIjcJC38MrM+/na
uGb6AfLQwqGeQH2aje7BEbiTXGmsJEd4OV1ofu1vFOQV3y/0iFNsEH2lM2nWuD5q
oSoFcEMbjx+59AFjXk7UYOXy/RVV5+VOwtP7MflMvIqOesZNsxtZWQ37A248bg6H
bg/Ruw5KKdJkBMhQbtpcnisBGIRQi8K9AxFgABopvaluRYxdi8u20Z59zrkkbZjc
RK/ODE03/cw81ImjCYny2/Bq61dfxY9FoI5HwZPNw0sTFJpe3yjNBnkmcV02fgbB
5p2lm6DtUoaqH9EyjoPerBoeFFcSR0BmTzoB8V+5TTwRKudZX/p8ZGIwHpjk6oxH
/syXAW22nGewukq1TSDu+89epdSsW8B0Q4fdVz2XkUY+G1qSEfKiAzPRK5z0fXP3
qMk3EHdH3VczEQ1CbahS9p7+lRJoDALX1ZWnd5Evh9GUKxyYJZNqxQwmlS+XatQX
S++UpWIem+RTLgxSVT557cpxFACbVwMvldco0gLQhr8ULTaS0OsZlzbINwlMXHb1
fzGZbxQUN2ZGoDSTIikVS8tvxoqnQvbindCDpueGoFTSUFMZ50bqEw1IrsRbWg6M
4mC5mbXdiKozV6yVmEV702T88eBoJTnN3bFoRoMbqNwo138IVUMLGuZ0osA8hNGq
Q9H9jkRN6Cp9gltUn0Q4gT14dzOZLAA9JYtObbwjoog6oNh44rCCjEIFOGJNh1Z+
xmgEj2ozAB/RCYPk55FrfWx198mvFqZNB94RyBvxPd+rV8zdJtXDzTUhNb9iajI+
Zi6SeWmxb7Dn9I0wLHYD7Zxj3fCmGeQVwuzOzT87LFm6PToWgl7JCcf5Z+JcXeW6
uaJJM0b/UMS9YVjp7QV6d3uDCgnDPgyKROryaNteYWOuERExOk+oWHCO/NDn0OXs
HkMUkjl/JIzkvmma0GMYqG2WF0LxsE0GRwbU3PzF7Vagt4zCBZ6OrTCL4j41okbo
PvB+9ntkoo/YPVyjxkpQe4k87U+RzUpLLQWSMvDyiNsL1ODU5Ce0ZN2CFB79kYx8
zcEImaDvbIr/AwJaviOTEnRVz9kuA+1kaOWGU/0P+GCIDJsJgaaaebKM4fLiAFjo
tsfeJvtMfpCS2gg3ri4XbQ8pKdM2FjHIW2tgAJTFsF7vxu+MeyIZtKTOf3rMAyJP
XScgTrqEA2eaR1IZ9EK/0wsIZXba6ZC6rJoRi8MRgcz3fxYHQxTRHfhkKSUPKC06
YagrLUEuqvumsWytY7iU+WD7gZ7yq4Xy1DICgO1wyRMt8U/rsN18IsJokvRWjJF3
pZHkuT13MAbSEkeigy2k/2Oaq7zD5yackr5X8qfwIoXkIihYh8Ro0K6Qm5AXiLwt
cpXPEt4kzFXuoN+nTJopGvWXpkaATrhyNZegaldieus+6+QKLgwdL/hfsIBrRy57
XWluu6TytUjaAhbQE98K7bh/8RFhy4HejNBUOLpSUQyc9Dh9O3h8FBVltWlAcyd3
7pAmi0rJrkUSp/VDccp3FeBMhTsyA8qvZWw9SUmhg2je1NveRkPW1LkM+Tqfoazq
WwecpwiuBMwb/FlDy9Ho69OI4zUWBDbVRDlXPA1J7vT5fX+Byi1D9z2J2fPbCb/0
67o/2gQ3OFimilGavOJkLdraKaZEovdxEbItaPZUOAvbX2QcG6Tt/h30gNwYPSDT
wdnhzMoaVX7ftZp5WChQJjmajE/N1w7+eAT7sgphbnrlbKOsDprnZ9zuADOSyTiE
TqKSJjQFBqVVAv+ACprPq9bjnskVsQY1NOo6S7SxYnIccM9LUyj28Ot6EuSAkklh
7auiYJ7ih2zO6620ms7dYCQV8CPD7AWX0aFerOFjltkVmjVgVJG1JF3qbxUu6YzO
VC8prv0KM+pByP2FbAJiDnfhBmP3DyGTlCrmrg1sLlzQ/Z96bk4uV4Hx2aKnchDG
ZiJ85LMuKZYdw8rnyFKkG8i60baJEl1Ri34vNJY8M2U9gqU7/3MK5eo+7qj1Q9Xi
pdPyvfJzxJUksJg6ZD37z5TXqSg2z/ijNAhImiFN+wMH33jrS2JfcJlprpZyNFiB
Mg1/DGRFeql9gcyQkG3fLmqqrcByyynCRqOYK/Y4lWaLz+OVi/3fpsAUJjNTdw7s
fbyOxJ0J2Jtpy03isjm+Du6PMlPH4nYLsqv8/ghTGzVre0zCB+9+I7PmvDA08z2/
5KcEMUQILYSAO4ATSblXwIUwhqwPDaKUBW5iRfZPsjpcTHM00dW52NnigR73lPtR
posQ3ZjUyPX4wqSKGsNIqhSyBi8115mSvG8NErgULNwz2XYjP2mXww1DRchP25ua
6FHsLryu6Azxmt9wwjF63LzLq1/d+rSU/leJXUkTBlu3mGPtBwL4Q+UvypS3gKKK
V2G7KbHfElsi2eX3EvsGbR+Gbd0ngvBx9Dkm5U9236uuo5JrCmwPIgP2usAkayPf
7SNLXcpfVBzC307QK4c29mScokf1ITYsqhvSWhk3AG/E2JtwuvGXMBCdM5IBKIPF
vz4R0q3itzvBXpxtCDm8xk0N+tHrU2/4n4kpEKPccb66YT2b9hLCZv7GtB1o+Gyn
2kpGvWgdA3LCxmJ3UMth5JZwxQF1kLqzAd7QJfxl6bqmlwtqUCQ51zHd5cIEdQze
NFSuNuf/rvdkYAkQpkMuPo323YO1avYLo+NsMw+eXU54mw1b9eYOVqtlBS27ebSg
FKZxh45uwTahvWqtTtHv4HOwli9cTNGsd4Px4OStT5UZrHJyF48eDqN6I+zqO3hL
5xUNfmrm4gw1k/yAP0i8uOJTJQKcQhcYdRCdFfKf5S7lPPqmeAezjvGVW0n3PiGH
NkSglIY1+lcJLhmsG8LgtdyHGKo8ZiiRyaKw4xquivC/AvHfefm3zHD84qXuoz4w
Mu5IS2pkdu/WbyrgK+FqMAziPmIDIKrOytCRuAkg6rZjWcKPVdpzik4Zh9xJRrK/
H6EBywhcUHQ38NJcHcFAkOH6DVc1BakYdMuz1M4kmKbX2hcH4XLk6QkeVsmeIUQD
9NoktMC+ENSJc85VITfAlrvfqs7cLxUDkcPsC8Q5MWo78+L4jNLCU8508lhIMtHO
Yu1rXRVzhXWtaiAELefmvNOvAPsIFLXknl/IgbcnghG5KFtwkqfbqh/PqYXYTkY4
oG0ZVamjrDI/ddasUw8wHVCqnzjBkiz44jTFGC5TkYaWqbfGS7h834cI7H0b9ZAS
5DyKQelJzUyO8h0YKVBakIYpr47IV28stGwSX3xF94fJRs7p/T/i9G/h71rt+GmQ
xriR9YJkFWs3Xs2AlUuR6ByKvZA+BUx+AVobAgiztEFnJmimR5DprEaxUTTD4yBr
LAzsIxJcEh8Ofz8D+bxnMZ3td7R70KRWMwFzOIL6as3PGCswmRQLf7sPirdmDI3t
UEjMPhsEu91hHuOsvh8wA23mSncL+lgUWzKnya+eNdPfm1MLjRbEVgNtw1z4vOGo
SDn4+sVfYyo94jO4paQc9XT3Le4fUQJR8jeDilZJvmr5jzEcjVpguE5d4tyADehL
x9gO4q7WqvZPhiueuwIsEaHG8vEZx6pZGxBZytVk3G+ejztjG4aUgcXW3B2Y3tL7
APAVnRYGXAKlWM6wx3PnuPK5DhMmtqlaxKwbjmWrmg0hM2CZ5UTwii70elzL9UZQ
OYjFO5hAfU1x/+XfDadoa930z+HrwBbeik4XkoFDDmzImNJuig6MDCs8RLwYtIWd
znuLfC7eLs0q1gk5/SoPjpd4Il6RSsLrTxfNa/wJuivMr1dv2MMABb0y+h7HXATq
LJKfnINYD8qe5tgIjcc9AZAKCnqWiaD/+jqbwI/+DCTYbdFmV8NDKSPWXpLKxsMG
ZmVhJ0Qo/xCkhDYD+WVfAyQBgpQnDjKenrtG9hgPQ1KKR6qRDssgwcOa3/rRN6Sg
8ZeCBrKvNv9qfEvpMv98BzwolYyJqUUhDwmXG0Hsty97STvv90uhNr175wUrv/4X
MG8g++8K0IU7qHXicLDadLklAmizpH/TrltcngesP5q5+UawpdC7FGN8jxSZAvVN
jCR1g3N8p+CEpLJsRJFn8F6gN9K9iE0DTLifoGf2STLvGYnnLyliwp0nqYMVOH3/
lbZmSmpdpj8t/JmvfPuRbIFfyZwkHEYMPm7cEjHwJgJoKzSB4IfpkM0pYJ0sUMEF
LN0KFQIuThXPNOd9kCXBjikVQiTXjCuSnio2vqpFgyjQHgERTxbArKHjJ+qA/GR8
QABvZuqI76zQipsAD5PVkpInlUCDO6A9uR/A9qa5ujVuOBO7aV4kmenWQLN++0hl
MIMV+ycVfIlHA26xJ+I5Wn3CuGrEcV9sbog1dkYE7Zig+Cer5r3GfD7vvhZLDmyS
3IoM773xhNa9EqnfX2dtKZccn8wqIuWJ2Hvlpuf4plwkgDfohh57YDVM8dbz+sF/
EBort8IZYbSf4Zfo+8l4hWZtt4U9OuY3aeB/w55THivl2JXLTz4kQVUE0ZvfoSIP
VNQlwQT6uyKwNyBBRDzGjuR+3NYiAOvlCsGARZVNDdaAifIuYzb6S3jUuETFQbyM
lr9NdFxUhnSP1cDCJACdo2/mnGxcJ5JID30SQqcj1fPyn+pRizERMCQ8ib118CWQ
W+VTklm/Z2D6JCks92jF4TGPGFrXf6LvLwxh7WbZqW2NAXwwJL5a41wdoGWKgCJh
xVya2AI9+5vp1S1C6Mc2vxgHz89QZ9gD6LJLXrqH7ej4nSo7c0vXfy+1JO5cji7s
z+6OY6MtsIv8uCRKASwobycVQi/nk5ZWzEfyr/rAJZHqSMVDE0SyplL/fVFxPClI
WLfuguWWJiD8+1PEbM04//4a4a8DclpZdXDT/V2IoYTfGurmH3iIUPv5vbWDvFCv
nbmtHMLBvk5JplSJSaxN9UCB+CmrNRF3h0GdY648rv4L+b1TeNS+/VFinW9I4F2Z
XPiTRk9PmvoH6WSKezUojXZkEHeXbngXYHDIx0QcTp0+cZOG2TBaTsfdwLuPl1Bi
ohvINzfJJ2jpsKgmg6JFUZIUEOw25kZ8PY3PRBcioRBoKRqsQH5FaXEiM0g5HyMi
Po1herUJ+2Gl18wsgBERdg64Mu8cwyjK8RNnIE4DqfcDiwU902YFyLXgwBGT77rM
YLkRHrQj9eiplWwp9yBL6xloZkEw3LnuCIFZJNmJobeC/uee8cWD+RMLzG69R0vF
zDOpw/v0Fp/7RItOdfCjvOXzMMN+2/3yHSPxQOvaOeCy8PN0I7y0PYVYx6r4Sh2q
MhVP0BhyNsNz1RzTJuKtFBf+iU3be0HXPKBL5T2/U4Y3TZkDdKw1dYLDfh9SIhvo
7NzOOUGxfiBdj4znZ5V3dJ6EtHGJLvJZTftK2TgkKllzHda+4o51xkRHqrbbYCQ2
YcAjbZolgi7QhL7/wGtCVYMhU1KTHXLwCFR5HUDAt88DOmNu7Hoff7xSPm5TpQK2
27hExU8HcAk9ZwcyVsW77POmX3Syc9Q467seOmAi8iizHAA91BnmxbLwklLp24Am
ptFqgL1fFuTYJHKzfwRmlRGMIzd28kL6Cx/skVORlBcsvojHa33Cj0zvnueqJOlE
W/z7Kj/4KzE9SuoXYSSJNAmyzRkaIcJ9dtetrKF9Z7E9Ru5vHfuiu+hYHW4RWZoL
DZLY0yCxs7oSoSHLDpvV43OjShXnNN4LAvKzs03Ro7RZdOCLBEo+dJ6LoRnaQiWB
sW3LsYBWD/OvYCjD5V1ez86CCS1yBdB29l6ImwjkSRGToVdhIoSIJRf5u+O436pR
axoiD/ZFL4DverYD0Kj+o/BfZjpTcadQPiAjcOTx3XaFCs8veTvl2tSY8JKLobbp
vKhDjnEZoPumgE7k0+qwNY2/fIzx7c9Un50Z3q9RgbtoRNWYi9/q9fVln1Rv8/oA
NqpxJQ/KttxTYxYUUI02lDIYOPa081Onv0shxEO6iA2eOAah1FLUhw2os9n5xHLd
NQ+Ae9YqtGKWMwvziw8PTiBsaOfneZGIQNOc0D+ycBICZ61qWZzFGyObMigTrw7c
BkyV8uYjMY8XPQhI/LkSdh+ACUjYUNu834sxT97u1o2zPuxBWRN+8ueMCUeGsRnk
J8xu7sDgR0LJYFtF8oGUtpZ7TWfCr+sdQp9GPXWlmKk2vwY/bSMKj/C6Ebc8G98M
8jpP4/O/0ftiuXMSJJC9cOgp3x62V8l4uetcdXbUA53zy7T5aYhN8gJd/uETrvDs
NXy2FMvUSRT5HeJS4RJukI/pVsxNLm+8H68kJkj2WMCg5v2dpwJBC42AlW2dKvJz
PEd+SnGzWk+Isn8Oq6a5xeG+F3J4V6WIEyRArQLpZ5TfV39TdwBN1q5URBzaNQO4
8o8MgT8gkzQqGhlzapo7LkjKpXp5xDDmkQtqBa0r/Rd9B5pofhT8zpmKcUK9mNxw
/DEv2cd2uwIzHa1s9sOmmkYhuZa8iqqoTXrA4GDsEiHAw+JbGqHYwmLpsWzABXka
J1mvpSt0buPRVcvRKTPsHtO448BTG2IYuQ+I42J5TZALKdwhUMgxOiO5kkysdtPq
c62IYIkJxnT5BEgM93EZ4a07hpXPWry5uUKAn8Bygqb2unWc3vZmgA/+u8PRJJUG
Z0N+ZIQT/mzat3R/R4XT8MtR08M4ScvqoeiMKgLdIzo2SA/xCbWgm2GndpH6Y5+D
6PMyMg+aL6qzOE/nG8WkNi+cmsCkMmyMZ37vDGYDIL8dzDslhPozSHz0lkYg7C+e
Aoxli816JXhPGvQbM3s2VeKWlP7mzubw9D1zgi5PrQxGN3flw18WwW3vKh7Elaxn
WmRfCX0tqrDZ9EFM12xq3673GPnHQW2ELtKDFsZFV5vf7oxn28hYjFchm+ESVok8
RYBUjsTv1X4J7Wg2N8LfkqzeStqvzWQdfD8vMv9lKjn+dktAyNeVfxUg2jrithbf
rbZpaW5QxrvTdCoc31uysr7PSGW47rrh8WYZOZEsOzkPPQOby80tLYNAAfZuYcyU
LIaWjmWHCve0yv2m+YDkXQ7ohdOfU0xYhJlBE1B3MRub9LJXGCbjelPa4DrXEtsC
3cxomXmx1iy8uOwIDs9XWv9H9XbGUbsRQYh3pXQurPr0MMJUAp5l5tPS534glHZu
ZClB5CmFsJM+Ucg5w98kCH892Fh3Rqfj4m+BjD+9oDf05PK22XY5n1DvGVJa2Nmi
CjlW2yn3HgJrgg3MEgZdLVvJ+WrXsgZfGqTexiWU1uVIqpL+HRmxVQt9jIzXoY8W
PAkknHI69W6BinnRF/JgmhgUoUyS0M6RLlZqDa16jxFf3C4c41lHNAWEYwYyEjbO
zlJTtZYV6Rrr4qAw4SnY25/Ta+SlHhbzsS5lSs6YnFoDempuQAPw3FqGQ69X1y9D
Pbokc5Y+v05yABI0pOEfrPqqtWNTo+XOCjM9B+JHz+ZVqEw2ckHqvZrzkNZXjqx1
bpOjVbyP8/kh1NBkqvO7y0U1UunBmxv8jwtGjvHaSgCrrDRJ8/FQKql7ZzeFkGLi
SQUSTELf8HFzTlWylNzofV9sxBxDDEDcj3B8KaFgtUWS14bgpL3yaIpq6QkVIgNm
VUtkLoSsH1sVLeXzS4Ual2q9Xm9AiYfpnV8/chirfPYVc9kiwk55r2ltQlY+1TZs
QJZ6Ahwy+sG4Iv00JebRvEn/4r552OIub3YgmVFwSBjHrSsDmD9i57J32IiC2AYT
LhjdAJ+BlZMHqE5WTvx4GqBceEXTvf1u/DnHJ8otBC4qOzX9WMEe1jUTwcW1oxzb
bjdNKfdJza2X0pdTqxNAWXtFIDrKeB3/Fo+wIFSeiVR7x14eYs9RjfEIgX1yoLsv
60CRQXd2nkiOs241ynwJ99N/+bYayK1Am9jFPsfq94yXlERW5m2OIh3g8jQo5jrJ
RGydCOkX0SWF/TT8hN4U+GJYoxyxBKAhNnRyvvVv/Sz4qaHIYC1bMJM30qlwFmsf
fygLYuhcuVrpq4INUIQ4HYdXVjjgNaaPMZP2Q+N6RMZT1iYCxgUGeZGReC37eEP9
4wGpAFEUvxI0QZZkSbuzK1hXhAKNp9ZC5PJA1bmI9A5WUUVewtjqroUF5IWK1aNO
uJUiR10O/E2ucHuBCTn3IQxvPEcfo2EwukJifxHtiFqJ3xGZPcxy8dV7rrHCVK8Q
OofO1zHIPomRKBiE0zIOP2XFonqHRl/WKzn1pY8yGpBoerPM0LKZorcSPYJqT66I
UipRihhzwGPBs56C0NZcnrFC5deh7CriUyVWm4lmNU5Y3YHmtjWloOW5DHg/4Hpd
Fv8ukKYQ/gVRJbUMHe3ScgZp/Ex4yfmWQYDaqdSUovv+w5pVd/vTDkxeods+h/hX
fYyMFfTy5Fotk+pUpPw1/HEfh0DBKSm4R33oQ/zFNzA5M7efHsxeFUd2QptrmhJ3
/9du6jWbRhx5NgGBZyCCkdp09aMeXJxS/RM2gFXy6Sy/piG6/xDIJ5qqwjL9OJAk
wgrw9/AsEPYLuub7eTnGbNYPaRph6ur/drAooXAClN4KU7PyUGkf3pDvil3B6q2X
1QjBB4a2CKYhfCnT16RUwvqn6GkxVROu5kqlaKbINVuUvS2a5Gg2JmyfIVi8Zzoj
j9L0IfQnXBG5bwdZhMzOhCE0VDnOMdD8OZYwtRQNF8tOdw4K0Sz1dzM5Tv90WDrr
XeaJynLK4YlgfsRaXuuU9mt9AOqqqoaqKcTEYmFGlQAArY/3JkRXfcRqLBNj7mrE
g2o1AisOSy+jXG/zhFrcJeAnb7qvHGHn2HRERFVOPHCF00fe2dXUhJ+YMko13onR
MaY0qeb94FnXhLyve6kpCtsOnRpEOyjK0n3oIcXutS/+enQ9MFhB0AKTcx0694nJ
OyXjwfcORmNOPSiN13eGDAb1Ed4oQSv3SR9oG0MaGN7JBtl/bOJfdmbMHshYb71I
gjtV7VTIct/LazAi/AF3MuwLSbHLebj9AOuq+JPm4z+8+ohzfv+zSfkvujwMsfYH
hpSuz0VJB1jva8KeMCUgOI1AD/GaC8XmndOYkHf28J78Cl1vD0+pxy9xDFg7lsIo
yfw/NZCcrj+6SFsESx59SiF0wP+wpaT8SCblpaxK6va9NPKyP83klgGEDlZmwLd3
+KTrLpQyii3HP418v7//9mM/UYK3ET2pAhGXo8xZqsvW/8rR0d9sTzSdO4nZnuuH
z1s8e19HTrpo7+Rfl84oeEfmJMn911eD0vo/XaP/Lb2uWDCswqzeIyUEaGs4mU8V
psmCxk8lJda+EytURyyk/ByncEuI1CjgpEGVb7MlSHpdvCqiSSC51SGrI9PqCBDF
YMf5Q//u2ZqjyuJkinQzLp8q52o3Ovw3R6XCv1zhdUypejbWqGy7Cx/2ncvqRIeD
A1lQQ/TC5gjsSs+TYbyqNp2ug3ozZ+GwmRCaw9bY2hAnyrDdiYzYmKt3h+yFDzx1
UCdo8+2vcIWvt8WhUBmEhBfKW88dALr16ZCtj4fxEVdCsWgIsaMC0ui+mJ9M25uJ
GS5xEQmflh3zFVXtSxZ3dTwvBePULE2My0m/d0fHmAupmyexY9BjbnU3/wgG3Xcm
N8O/O6JXHQLIma47ss64fnzfBRuqh89rGvEql92DJiiKNo3CbKoEP6FXtz4TGKMs
eaTZU/7uBrkytOclyTfb+QpHlOoUMVn6Ytw2lqtyRBHaYszgVoVT4JIyjrNZRkOx
2ZMyB9fzT9IeRANqFgLkb+uNYsPWWIVb4gpFDFCxGGsrt1sbK4fjwNwxszaTtKHD
5cO4azsC+3WHQ2U/724is5fIPLsb22zojfF6qZ2pPcp2bspCXWEcfYM6SIWLM29M
aND+sh81ak5W+ua4qhkxR+TpI+u/Lx/oe7oaCuuzgcbiKGqFN5IHV0RuIXb+/O6B
XHhbar9eqfa2qvcO+zK12QxSf8qnD8YET3Liyc5dG5XA8yha8ojpcsdRAjnb3Wxw
3ZmdW9i2TUHboTWYqa0sBoesFIE29iREaXZ8HO6B3/eMtynia4fGr/j8Oth0KNXb
kmobfqAamDziATK+XK0Fhb9lthiRwahs96CFbhV9AUHaJzayPdIBnS1Z4FHkhoF4
cFwpB1dfwBiQ3MrDubj4r0Q7dXTerEZcigfhRgx9R0Uw6GcyidT2A3egnXJ+z+W/
tL/o7w7ynjgGsatoKtXEoPhjVCKk+TzGLm4Re3RnhWMRIpFaaz54TLq3lg86mo11
OzI2HJJGX0KQuOWSPw69CG5L2Sjh34DoxNQuXMdGvUBsShepV0aDp8LX8sp70VkV
HPy64XEtx1fyyc1SX1F/dE1fx6k7ObupqGlxX5jU8xLQwx7vV2tjwLQOHX2Lv3Z6
2w6brlNVgXmx9MTNuBKTA/UddArXovm8/fNbWpd0fRaI4r51espDIs+vKgiNGBEx
YvqycrUslB1HSSILKsKfo1MFLgtjkLBwcQaeIPMvbg8gUNAI8hf2/ZtJAaW+hR8B
Drt+psEXWvf4jiUdhgcGqMuWP8DlrMXdoPVjrJcd/FOr9K4vaUlkA7j3JIoLINP3
bGx4NYJ8UQX1wWkEsiXfT2zdDD4pZzmNa60AalTajfZnCgi12Fd0FNovvSVWkDcz
QKSzRX+hbq9VGWX46c9CA4vQxr4noAXmYqy994yYL3pwCSx44diOJSPbzgHNWWHe
+Tu493oSJn2hfgO9EBPV4cLp9BzhojJsnd5urLuc/08QDFxnSvfFFTgYLv40iSYR
d1wRzDKYbILI87Grk53ZGqd/0A3knX5IeXwMIAOcq/L3blfv8HUlfn2UeYNRJHdp
3GmpE9ySwoX1Ya0GlK6lginS6KS1cYy/ff4hoa57Mzq8NnoZZ5eVZEQVfvq3XJ9k
qJq7IVdWKSSsMsRM/70scaSiYcIJ5lj12lubDs9Gq6/0W3J1vhvLJtksGquM4keb
dWnzSOuWdIYviRs1nEC6SSFL77ESMVL9Eb1+2UwCGxCdZ25Kw/zvwWbcwiLVJhdx
QN4COANI32TllPXjhgoIr4uO2cPR4v67xjZUGdNPruDEor75xEP5U7guv7w6ahWE
jswRsgZtXsNuD7XPDz+ohj41Zdwy7PCxlGvDJ8mWdq2JoA0dY60zduGkgbgMr2ZV
B5X7jdiLXY7Jktf8QzymG+KLaRyvDwRN86o82QoO+2/uIfisgOCKL5vLfTlL9A5X
ooIT+lEpUnFeBg5E/7LhxlDO9qn511CPHdC4V3spdObUjcvP4TcqFI6joBRN5TNG
TDckwT3q+D7n5h/wvGNzX0tylZGBBR2I+lvfz18WreSM+3v8e0GTals1ZQl1M+vj
tpN5Qg1PBr+x1JXTcB0pdQg8UGd/8OVYxxl4vA2MuDW4+Em6Ifs8Wt2yIW1TRmCS
a8Ba/ucH4XfnU+XI5KPdwHQbAK57Rcid8bPr/remWHx5jVHu7Q1o/20CXben8ax9
7mTp1Or5c/FGMfMZIf4WV5nbeAu2Jp+jFGs8n1JEoy0pg0GV9G/emkFoCdtB4fMr
ggDX1ZMi6XZy1QmB88hqvqFYwWjGV5WDFtOqq1gk9aB68vjTr7TVnL2vI26GaAvb
UbGBKXmlxdkzwCLWnnFktPcF3Yuu82PYQonQWm3kwGS0xxnqj0mOKmBGAsUPBm8H
YYo/qNheTt9nWa2vKXEj4kYzTgU2S4/xDsvyHU/6QMusmFWVJtiPOQVjo8UUMlCR
oJe51BvRSsqsAW1kj0nD69V9/SGWuwI3CykZ8bXk5j2D3+Yal3eNFy7HB+vnoNSL
cUwjd4YbII7rSbrj6GMwxHijwOwfIcDMf86iw8IO0dG44iBsPDypPONVxqh8e/26
FPTymfKzat7wo0JZboeDJdBAVKWjys2h+Ov16G5V3z4oK7hfhYDGfZuTqj/sZv+U
s7CUqrRHw4GCksWF6qlh6Pr+I1a65hzInHMt+8zLiBkaAdlt7km0zMbjEIJXgN2G
Bof3btK7Q76s3O90q9BJxgqO3/qvQAgLDh4x9zB3EfK3ezfW8FPtI6h5ksX4g5ju
KrI6StExkaOPnVSwE1N3/1qyrHtN9JOewNE2LKQ1LiBFms+cFu7a/qkxLsi6xtKU
QMpQKT23eFAP2Wf2YnWya0oHnbAKv1vZpjrXfPyq+t+2Hx7x1eaqonxGYsTJnq8x
mAHx9HG13hyXVX3+N2w+mSl8cXRiig9u+zxLmoztb1b/kLiBZWtuiEJnY1SlKlh8
xnS7BWbQGE0dni+to+C/mCdw5tEw1WPaGuSqGy5/msqua5F3PAU51e3ySJUd/DJM
m5mQqNWo9qiqPKuLgGtuuLbNXpm8i1XSlxzKaGL214LukaeG4RBYAZkZMyjXZ80D
KgsBEZ5XKmuJrf4AOvjjBIje0OXhJUjwvoMBpfdB5m/FjqsmimceLabaUsUl95/y
WvElrsdygTe8nXzRimpdlmMYNSIbvXJtovpjEV7YkN5cUUwlNScIxFlAy7ZPNYtm
/lO77DGRNp1iV9C+n35L9r+XnMg6395UtDI4tcGrOS5C8pOST1T+ZvrqO6p5D9d8
XDevChbo/d3WQkIy/EjnklDV6eGast4tCWtdlsdIqzWR9Xe8hPdlfyT4RsMT576j
cm5bHLJ7eoxqsSSP1ASgQ9582sWMi+AP6dXE1Thx8tzesN8bz9RVGsx9dDuIFvg0
oDwqII0ynYflwPgf0MolpuFnthycbyNbwiB1juBaT/0E62md0Wh2p90Q3yHJuBqh
vCEkzt2EGD5nk141q24DHCU2kEoKhdOwLob2/y4G5vWXxpTSoqEheROom/1YGajw
v5I+ZXQdWb73gkhrm9xhN98EuY48ReQ4MtzrARKAuISJLZZ9+rcuNa9QcHlEe6td
tcTwZGWI/Ae4mhchws5sHoTZ985SCriHoKihoAMwj0umQeDMUFRSGzMq/xG+LjQO
cx1524Hsw8UqSDJXwxL3m2PTtYp3oEFoEewOteIPxxofgKFd/2e+iG1Qz4PIbaiy
YihjUV6M7Cc/V0MXcLH1KIQYAhAtjQCxS5RjFo5G2jgU4CyTe1vmFZQ9VEKMvDYs
yfv0jouKdMk8NEmkdA53ckNHNXnRY2MvK4T0wxmHdshG4aDYMsF3tqoy3PTrjr/8
Nbf36Gkmhfy920MiZN1pEAFCB0JGzSjXB9eMzyMKd37941S0vawvZZ+c40AD5GMM
+sqKgsAtGDNS5k6+5jQb/xTLa5Q16pf+EI7SsVsrwKuErrXhp8hv2Vn4OvghpzNx
Z393jCEdf7dUSwMxWYcdLo+wz83UGSxapL4GMAVgzGwvIa6DRawo+5/Xet9ZV+Jr
0WQdGEi49Bt8sGW8JsZbLrW/IOFhbI2rwDUys2oDjtZw6lqlm00ofvXsy5TRIgfv
FLBAzKx98rvlL9D+QR9iiqpWrjEiY9ibGxr7i2mtz082Wc2aaZyncSatLNCSCqXI
uJOuctFxAHUp9/a2eZ83NdYmiFO1o+Q7E3alXhSOdRpYR7lpk5eCjphDwt+2sqDc
GCY+yTUfAniNEudEhnS1+pv2MEVdKSWArpQRoAaowF+SJk/dFeDIW6CyPAZ7A66i
Yl8Bb5PPLgtU+sIsgYFlOqsawkv+Rl/KHTN4sO1rJFpX4WEV3IoREkQi/Dlr1WzG
0C+s/XuJhn/MgWI9emT6MZaZj7iHvuIgBp0gajHLXIlvGU8x1peRUts135hiIRPB
USGB3LHMMOatycbb+edxKvjapGp8nTBi14SUw3KQkGBbTb1UWzujEd8XOENqAVeN
AnAO6xQpJ2I4RYZbTm+SFwVnYjmE/UdcmYgVNW+b7WnowGiEcz9fqlRHvKSf288Z
z4BERjmRgOX4/N93dC8p8KsFXWW7Khxu+3t0C4Lu4w+gzIO7ZqI34JTiyWhF19Tt
jEQqnRJAONIiZJvDzqU0K5mE1ZkKrbZf1bCrCzW+3ylRqSL+XS3WaeCifL5jLTvH
FDbJ5GxDR1hldUkmw5ErsTh82I9lFJP3SQdT0KsgRNkXFCfPBuQv0ldEyb1WPG2P
OOSbvdhhiVLc2MezvQlwO8P6F2rCelFxkeGdF7WC0jy0yxiZaLwlKC845cOw2SEK
5dlPaOTEiB5KFQzcFACNe5pIS89vpYxDQv35p6LUFNOLQBhU7ZuwXFPyweZZ4WCT
4YKh6HrU3Zqq/wnqs0rcv9oO1w79HqOZbepS3gvP0PkIpg/1lm3n7IwwnLxeAbcl
mDNQBaoYiLFXQ/VZBZ5t8vZoyxKfYxV3GhFtSJzgC4jREoUTcZeGOmkx6gOs1ksr
HrxRw4QGpvjRa61CURhFT4UTrpUXQyevvV9byQlGbf5rta3JrZUgaVwZsVXk27/0
HjzyNKmudkn0uvQJTjCXO6BZINy4Ll7/sspyihTwixuKIfaIgudDPjRUmrpGVga3
aZuMIu+IhiMFuj8RFIZ16cqhDQrHZTwgH5dOQbK3Y6pojcp7OlOrSDrW2guZxAjw
laNA5yHf0e2K0hfJ31b+Czce4kiREdKoD4wfO+ucdhbQ9LiwDNoOClc+5GIrBSj0
tiCvYyNosHL7ep1t1jIzTrSns3qiR5Mdf7jrrWjSEiCOnESI62hlFVKJpZEZFXcU
jBLC4asAMkOIPgJcihnalKbwmFBipg9iSstvliM+nx02O/YhCUuGNBnsaVA1krBx
WHuMSuKDIaQL76I9t3jKaFbfetLSC27DfrSHCK7WQ5HiFq9egOQT3yJef7bvQ3dA
/FLo0Jq1gdTrq9NA6SN4+M2a6XnulhTbkXNkUaNxMmUCwzAOFgA3iwSteZpF9aWa
yxJl6mPAyScMeepUjEwrTWXE4Uo4SY0QU7dPoqlKYKiizoBLoVhJivz+nqb4IT0n
jsopC3cwT6ORdOsOc+IJ6ILTRkyJ3DaLHnIFeuBGFHALiYqIMREdpoES44M6SeAB
KldRCekOAZMlNWcLlxQuyDmElcw0p4cYi++cnVuYCKPXXXm+wsLjXFBPTdXvw0pI
nk46fhT56RKfKlk7zYdalHF4i/BUGz3I1Cn5iJ6r+p8mY0X3m7hJOT9C+eMxUiQr
H4upes857WeoamCvROfpnsPTvv/fpDIVJoeG9OTgE38X0bOAq4xXOAwg9Gt71ssa
SVE1mAhQtLGBDtCe8puozBMng9JEazon/6zrkWUrBNXDsTUQrKzp33gdj80TlHJv
IKF7iB+5Vk1yNM/3AW4PatxwL93YnNmSZAui4jisr/hfnRZMkd0qOBX7gtJyS+05
GoN9jWnXllMsrQqZ0JSjAC+V7kL2b8zQmR8/ZYuNb+ORNr/a8KvTNHiA56/VGnzi
uezQoQW8VuP8lmJnH++4TWeJhvbAS37BBRZfK8/MtKtFD0shxoPwfPDzegnEQPCL
W0z9+e4b7l6JBtjoRKM+MR2vXa6e8MD/ncA0HhVlNiOESthjoRTMiJU4cUrOzzdE
WmVatziLyswnYIOjIFEIv2gGeya501dTK2uNA3khRAx2X4yBg7NSoQnY8z3MWSNr
nr5nOev8maAvAFzlh847Fd5d9OhkCHK9/pF+e8+1TnB4NXI39jEIZDk5jHvQo2V7
tT5HzIGdRtIjm4sVrk8I8D3SJjIcT6IBKvxNBuo2g4TwF0Q5pN6r0q2BZ6bShCZa
Y0823AKp1GzaighWI0eP57OAHFqslfAOaHV17YHpxULDFTC//lc7kcqGqsLPaXJR
PWS7clBZFCig/ci89M3FfPE36beh3KTc1ArBSF0RDXxWcWR7RwXLVRi3aM1RYIDt
C+ccgffzlxQ6H8cpwWwEL7qny3PxOIteAnddlocyQlVj2jvQWmmnBdBDDaafmY37
IzZ+yYKYDXPFufGvMYBe0dCed4ymNjR1IS0i/6dBqHXsO5Po8mV0sqeZEwz6SvBh
8/aIl6u/q7kGPDdiD+AwgVCT3Vuv8FqvBYFIPcAVrMs1lQkCBIjKN1770NQZ/TRG
WASiEQlvohGE+CsKjJf5f9kOZ+dOi7B6nfeLfXYHP9PvTj7WYF0S7lk0AIYMasyt
rQ1BXVJiCdT873qWw2GXP4wnZlZPKtbM5QZQwygUsBvh8KBN8ig6UHnGnpq3Pcoq
KtxWwrHeqegUGRNrHw0Lr7aphPIaXTN9lEIQKkCsWJv3WOothk8WC9S+NpsGtBKV
REK2ozVLfvKAgaEAh6Hrtes/bwK0Jmh60v848yBDO4Fx+YAcutQoUqJcxg4S9j9Q
KtWidsHpSN7TYJx/IZMYe+F/rMLDl1NFYenlCydQBXZlenEm0X9cG/6n078qAp5F
ydNqgXiKfEjNYkkSTIpj0Kf6Jsjqa06TF4gpvckgf42iLuuH0Ss04LGiAsE6WWi6
F+rgbYkvTKYHzEFQ3M04oZCvqs4qJYI3ff/U8w1xiHk0sZCF9tbuMC73jUuZAXuB
YQooTKmtGjFjkCN0ioAyvf8a4sw7YTlme3IKrZZoiXwJInkV79PO9fAwTnR8N+M7
BiWfY58/RDf9nyFtQyHM8IwXXgJWssis/1xLtFgTtwN8IcrnmDuURkm97NCSCCrb
DRQrbC362Tghmt50w+/+v7ThgY4t07LB4aYdcXnXy8/dXpKH8yMPlkB0tWZCf4X+
JX0INTH5N5Gyej0Geaa1csbF1ZtgIJsAmM9tki3+9YBCOBpp8zirLIxzcbdjRvlu
pFppPhfMEOdfs5WIpwyiOXJLikmOgq9+EhE2LMint/+n7Q5M9hJ4Hgq+vwR4w6Gy
m+u3R38slFmiwXPWRCA8BfLoTz0vWwa3JB38yAoz5KrenxkJBMCYBSu50dB98sGr
fa5VpkfAelJYqGGK9z2OHn47/gJ6xN9WZCuWYFAjqgxkBoxIX02C6ERynkqMQhFv
825MUcHrNPuOMIgdc1cg6OhtIzHbJlWAio7p9MOqtuyE/78i1p+ve0pcHbPEpNPx
utEGAXgd8gNqX/s0I5HYG10dilrRrdrgCzzPCy+d7Hupbx+cSYHpS8utTsJ28Nk6
B8hGaZIqF8NC5NKkfqs6sjdF915ddxwlDbt6mt9UCXIvlIcLYbc0cGwQYddD7DEW
4rSMrcYc5V1xKQYFVrHnXQb/glwnKxxPEXVJiKJUcv86TytBuhm/ha7V6sP0Ouo8
bt54uxcTGcsO71zftR8yaxhZbqHXvOQAi4VY7KFvpDkwOotxUi8c4cYIJmBdOvx0
Z2eVnrgEUB/k0HoZueRFbZ4vNKeDWq/HmsIMoGjBMAQaVfw3Byj3lqI8XLRBywx1
WUpkpOJUnK2vaIR0WC91wF5TVf9fjOI+Q7t4hQyyAPGoIbNaYt+RtsB//vYW8rlb
kp1YzlzSxArVg/FRELtadCO4OAUjxRDdaXXnW4mM1SfcLEibr6j9veZ+2TzQXHWB
KFenW2UbKI4fqGRoQvpGGUBINdxotgALIdZ/02ja6pwb736j1vk1nubbCNUSpq/o
/Imqqy1+OSCpDjRp+dMmkG8/rbmU9GV/mu1oLxxUQH+vxlyBQe6+qq0fv+uTJxmk
a2VizZt8y3jQtlIu/M+OZoJra2PPiZFqGuzkDPAJVxNcNz76uAYvqay8sBlwepdG
qgSWLYaV0gxFMcRCz2Q2vOilgEG+xcmPXp2KhufhppvYf8cgaBiYCgmg06vOcAex
3HlKDIhVd6D+0M/wbqaxt5fAMqAzobxEGuzgfdj9q1G/a9xmzFZbMB4eLILLN0S4
j0cS5PYypbBM4flVgCGcYN19g+O13TCEYgo9pyzfNSzSjLZQm+EOekzEnS4rDUTU
WBoCezZT2oaW1WNVQNCGkaV0vHURbfwW9R1i+iREPxDc+1ukhPlKwJ1jjgHK+92O
QkigR0yzXfuGCt7lchQ4zkYNZ6zZUZn7SsexNSVXMutOnYcqaxEFvqtKBZGQ3iuD
WN9Ti0vtFOeyvzbKAlpfSzPOVbcKmEFTQJ90vgTC9SsAlDbVAPYdS/Oh+Fg9I+9l
BAbGWPL+661zGexLFVQohtuO+cyvCL42bffm3oAnP23b3hkrBY4LGDhNf4Sihw5Z
nNa5IXOe+Q5IuVzH3STJAdu9fCDHpKoNHg5sfGpSitoxQUuF1YxJnSBg3klqxt0R
vR6NA4nxAhef7cnREADAUVumD6BzOzw47SlomYsqPdHW6YVbwD3RmuRY4bpfWq9h
sYSbrH/Uko0YD54Q2vud4WSAInh0F/3D+AXMzp21NXK5HwNp9+gWCdkr2YZNfVeW
mT1jL38km5oTRV1vsBIhuRD8DijNL7aymFXggRLc+I4i38cHYbUGBxIkC0w4w53j
uCNzyJbpMPPLYB1d5VS9zq9toVptEG5GDZ3lKArmy9PjOH/YR/4zzzF2ZtgSmbQY
u84Wudpk14t8VeE+7akNDSnUAGB0tC1qw32cPfIaEmjVHzvDMZGrvoh0BuX0ptlk
JOgyAAvifXUA5vBts+NWPRD9XQSeFF95C9rnIF+Tjyxey5B17ua1TxpiWtFz68DH
AMXBUhlv2OMfn08KaHMf16BsM2XJhoJGAdGlyeFkdvvl+GNi1Zu7XQC4yHHEhC5A
FZdZKFijIxA3TU/38NjnkRNdanE/Jy3TJtNPqwfbIkXfcPQ08JnBCQab8E4Rzbzp
0xweEZ4aMgA35BY9MzXvwkv+bQErxFOyivHW6WpiZ4z0uVoN0gA7YcLnklRUZrqe
DJaxMTAN5Xdq4xTG/sXQ27pMW873vj6jw8983t7e7FP3u9y9dPxrbZhrcPobp7ov
bYCx1P3WBlsXTdid4pjSATqr636mICeynvprr1fFzTtCNsz8fa90eJ+d3RwYSeri
OHDRUkDS/UTTtobpkvgPb8TgmDGnaBr/aRQLEgBVNjo+yVKea4/Y0RerchqWmx/D
6Uat8RinNTb5DY3zwNf6fjj3wVvvsZpkHISpleQnxC0/pxo4qhKkC5iwXfWMw5Yl
0VUHVVHT24nyMfjwCsOHNO8quHPwIOm6aTd5plBI6ZPfxfcwWGBPXC9hEUg6TzIU
4RF3lAMvfnRMcjeJZT+cH1kKkCVApGxp8SbM6Z/3PgFxvJoUyzt/5qhIyA81s8Iq
/FMXFnb/yCcZxtKpLYNTaA1lAqKPaF/WW9rdARVt0KXlOmdAXAmkc68WaYBkDrG4
NdLkX9YlV3A1kKRYk0WF1b5QXp6yFa0ZydaUx9m1woo2u/NpoJ9C3/KqS6AWgBiO
kjRBSEatVIzHPiuyDs1E4RZUAwPLNSkZIQZZkRJpi3MxRVVOrgcG4cUyZm/v+FVn
XisruCx5DxnmCkKNMONgSCDDmkB7cZcXpI203f/aGpXI+NgWtdc2pcv082+DSdD1
gt/t7kMaCZiLJaCqWzZN4GFviWL5tgamGxJemVUmiTOTpiR2GyypcwX0cTiEeNZK
v/BRzyeeUKhN+OcqgbULKRho9D1XWckfH7yrJxF89MoK8geYwGzmnwHEeIbNVjWo
jF7Z1qsDSwR6kNbs/08+3u41VLV+lCqsDx6NmdXd07PhAzyzDAxHCX/orjjwd2rG
LQS3GbQqc5YRxrT1/HzWef/A/GDva9zUCMruETilK3FAb+IREmMqDzeAFA8e/1VB
2aZ7XTgY6huOPz7WkTOd++eqkImmj5qMasX26ADezK89vrhp0RtVa/l99CDmAHhw
pndfgo5xVo1AzfU/MQ6IESaqIaEXQenchg5Q82e6lmtXFrYBI1K16jhtIxmAzmVm
rcAIb3VW576RzqWHN3QOy4YF350dGmMxq0aom1Z6fLhntGoijNi8BGv4yOjBCR96
aGLYZ0JtP1urQpjjDyTYBD0ppmUKA9XODkdIrtFBKAu/rhTL7fPcJstMrDIGVsIs
I6fq4N3iV36t8oRex6dfrdsx3UQPn3vU3kAwS5LppbdrNT3PvfDlaeLZ9pA0IxAM
ddydOvOYrV7QyzS0coXgsZ7hjyqUsMzjpT8iZ5LCCHHbZXP9ssKQ08jNVk9M27xQ
YT5YiPJ0CLeLHnYcTSwxjd7Piwm6WRpaly17l67zk9MMeyh0uUey9jkZJgNGX6SK
gQVDyQqHWSlkaHZv7B5WuA+s4x+X8EQV73lx/1wbXRcPBcTHF7UVd7G3Fxbz/O/4
V6JWHIvWQeedJvaosdPb4f8K/Pmlln/VlQcBZHSGxkUSyM7v8LzgvMALoofpEMCk
7F7koEYXfvlB8sOGcqn+bs4A3sZ7v3TEdwy+nATQApF4/1CVntOgiEqnkYjw/01F
Deh2f9iyEHExqTQzu6zpgHSXz3qJnMx8xb4AT9w7lWmNuyXvkFb9RL5ZCJSvBkWW
LPiHJq2CMvXS1aw9wry4hNxRIO/nO4bkePtKFc+esWYLQoqvr9Qz2+6asEMX/RU/
PPLmOKeInp8IJ8GmOX7veZ8dLceqnvoRzxQ8Emnz3k/JVuttYDlPsEv7MtBBA/yX
UOXUewnHhLDcA4LpAuZnfZTQ3joMX08tLhFS8wtMBVvS9xRRPZOaPH2cuZNGSXY7
uxYcnB5+Q5EmDYj2z7xfyOCrK+ASnh1fI5Sn08WBe1nCH94XWvRXyE988YtT+7wK
xjTYA+a8gG1IZ4Sjukb2Ex+RtmlKORyUxatoND8ZRHZ9kuQ/nPrY00p+6snhJkzH
nsQlTZmp/VqcvLeY3WkGN66PzNaDfax4D5rsZ6vTQTEddccU+LxfVCqckTur5K+y
bnnNoXS5/qVJUiAxoJZI7pAEk3kKUhDgFjZ9lLtnRZbceWaaqkIFSANkzQAvpykU
wxuLJEoPnd9SiECfQ9iy76kcbx3eDxDi8U0daGyFNvwB5+enqJv3qsavCR5b51Rc
YGj5+Qfc8LH4wFXiEiogqOgh54Ev6CEz1UCtuoXNEp/PRFvUqWm7MLSSuxoXtV+F
xQGFXCtx9NOHFJnfSjk+mH6lXqj1ZOD9XVltW6RvUEsVlHnC59wVGgRYzjM4bdNH
0fL4GCKsjsv0+ZY1AOXGkl8DDv3hUyQPCmBQ8YGxBqjRLGaqkceBj82r8SIUXS8Y
6wEEkn2C/QIwZT0qyhP+lfhcsrvtfnB5/W/pf8FcWnHf9pG0PCA/YsuxjGFnhsYY
bT4sWM2D364qfw+Oxb+fLZJHmOGjZtaRRl88mWBF3YsRCBck/ObLTFFnAHgJht8v
9eTAh27s88YY/RRR1QwHhqHZOUIBz4kddXn5s6bW/j9ur6QFuO2UpEiGW/mM6nOq
rxv/ranAIMtOKgVX3Tuj66vY4y3djSSCfzGCkV+Sv9NIe6fa6HMvGb5LXuz/3vYx
wRrwLdBXgJHfydRsPgVcV0ZJ39JRhRja4wOAmVNf0cNyHs1BvpZcsigSgw4CGi9J
5H4NA+PQM7u2YGG5t+AkZZy2kBwoH7ScHaSJOLjm0+G3bFVtp6tZfNxYjnmsok7z
McmfI8cA9RT4pR5bE2fxdu9xTBi3fMGB2oXHkSET2bM+5FoqLN9j1CnHodm1/P/w
iOsmh2zSe01j1CCxxbyNi//gFsqHCyyP4/HJHdMujWs4K8fOXxfzysHuFHoqZvKK
RYHfqinnUvL7fxxxpWrCn/bEqC0CdPCy9i9m/TDImk3jbTcDEL3n37FnMq4zqk2y
VkiWHG7oYIp7bfmRbfjVT4RV+h35kSbAGke4RQAvX7ytkyD2VqZc0iEor7nosu8L
Pc95EA7IWbGVtY/Q7UpQhPU3PqXWw+hNxcImfQK5nc7snp0hynbFPk4vG0DbHMm4
sp9mKh/Tf/xg4QzvOq/l7OL0ynKcQE91iJW43Ma+RZHxVKauQ2Jy5rjvxAiUxOfF
d6lfkc5DRSY/+Bjkq2qm6aBE44e8tG6RxUoffzD0TuNaKGJv57XDRE2ALzfko6X7
ycAhSqS5w99CP5AdWLqsWPumOVwuspKzTiy6EQlZ9x9fFDY3INb4y0k26ibDv7Nf
wgXuI4WtltAaJItYEZcAwQFLze65Tnn43GaTMnxcCGuRpwYgtU2UhDTksNtBog/7
Ss6Wil70f3BlIyc+XKa4M+X61P+zIDts0mg6OilD/Z+xdvBxuD3lbjo6a0cnnGcp
lR8o7Yxtzw3+ay31kkRVuRRCH6JuUuZn3s5ORQCNGhOHv222EMKJuGJA9BX/yJV5
D/O3uKcX+EqhdmrIg/XMcliqggOP1PlQO9KKIUEKkIDrlCxJOdKkKC+dynVHb3/H
pslTMSN9ewZ3ds2FViK/U0iecwB6LPVfghWGc6bFTpkm/Bl7xNUtdvZzJGOCLWPU
Nt4S1WlwjwbkM9xclkEbAdxWQqzb91tOoFYmA1D3M2wevKdhY2tHxOkmMtjMltEa
tJLaE8DboaPVPAga2vWfG4Lq88bvJDY4ZU2OJBNsI3UAHa8yeXEvXnwoTGAufeO8
dXIltXfA0ABQkYku32dUvJ7MJc2quQCARFSDzpidO21uk7B8Idia8Q93U3YJPrQe
FUDv2SsxAvjWJDhl/BUpUoWU1x5zgVPVOL17dF78KFUrIT76TFwpXk6MhHS0snVW
Bpapt4jj8U80FHK/nHY901hLokd8CM59nH2IU0VgzWUvkXKpcLCgt+AHGJxk/rei
qFG9+ExRK87HCMNCg/fALczlZF75SSlSdN9Lkqrpyz8o7V8FkIlq86bx9KV0sN5V
hAA3IBSkWrxlOd3tTMruOiqnR1WP56xiF6Y5igOThdK1MQy5Xtj5W0lDZZoOC4t8
so1qcGetIKTBJ26Dq1uMJ8oTIY2UInqUidJHaJO0RlYFxr2LEk8Udx1EsdG/o8yS
2S5g9tqJgobsh11prAjprOR8qB7b0T9awgxO+oj26uMGyvB+MaFbefJTTi8mMz+X
yO1znWZZIsclMfR3QBh6Ridfq1++1fwPwxfqQEE40jtbejK7gTBmb9eHHAnQo74X
N2THgRm/zU7unQ7p/MbWAU7I3/SywqbnKrcM5SlwURSaYtT5kNmN4aoXYePGZdRa
JISRffNVYLVaA5vY/axmyct4cezFBAVRo1CsVXLgyTWsb96YtI9G+dkGMYesFtH1
vcmQtRVH4yD+HqaG8gjGQ8BXBRwdee6mLTeT5/dIQZba08tgOOL9kbyRGcV7S63p
EwutzUXbg0nWEBZU3eO1/hiDkaxLFe7y+uEgNDBds8KeGicphxrbbdHLI6tQAxcK
r+wtWDM8Hk97/2wW+IIOwOYvl1fThCrZJeCBcQoabZ7heP0RZnV6J0uIg4sOAPGW
zLI3Wfr5ZeD5wYWF2CKtJSngJTHJKAkTCy/hQN4dq7PNLKqn6f/jQs5G54ljVl9x
ynr4uCrp4YRNNXAhDG7J32P9DMJRC/kr8e1S+ElIpgUnGhAKwUfxC1FHACI+NAdE
BLvvSzzyI8jrz1JJqMmc+tbXYi9LCLTPX0Pn5qy9x4RMrisv5c9yW1QUJC4Euqm3
w1ug9PtcCrBqkzKV+rCDxEeBIjpHci1PktUQ6RL9RUowqcZA1ZViY2wyQYqF94L7
kaMEmrHfZ0jdA6q9mHJNHdBvHqGkJmjNaSdwk7w5oCiecMHtg0FIwHI9S2RrQEdw
j+ryhaaLBHZo1utHZV6gQVwhamZq9xY11n20uD7O4IoLKry+dkIE49RW+SR4LXDI
jBjeuCL2Wj/rEx++VYOtZ/PNeYwlZUgwKTMSa5x7/m0h3iLOPe7MacBYn3vq1PKp
wYzRa4iRcfZgsf137YNnI57AXd7C5sBgTh1W3R9bY9Cir6NlHugHheFomybQ4rf8
hpsCXa3O4Y2bBlHUgI8KO7CSOfcgbtG3pvYpqY4YKGhZAUCBfiFQDCd0CGER06sk
TQrl3uL3iwEwoImOFXIZEVeHjQVnLbDu9jdUJqzLZutfVFoOSYM5T8TO58YPoWa3
XrCRUC6PbH051FNDkktTguqOPXOmgk2olqnMEps0Ypnd6B62qg0JPjEq4osMt/bJ
V8fmix2BTn5234CSGf/6KEVgEN582Rcldrh3ofhr8So2lhD6rwO0j4d1fa2YUNJc
23iyoDqkNKWvFFID7RuQKPL0nca5qkogfveOAUtu1vuqDIDBcf5PKT2PGpTbDwiE
Pa5rBV9x/khtBDTUAfu3PFsBfs3gHeCkjc1KWiTaJNkyW3qmups3OfcKJ1VLPltg
ckwhpXLFBdPNBRksa1qRPj1F75gRmc2Un3a5cLxiFh2MA/nej+ZSHqxSIMUzd4iS
XYDApasUWjMBUkWGSR91eHRieAKpBQOthD2Omda3XwXLWepaQ2IQrGebZzxPA6N7
2a7qYieDQJ4JvymWb6UlHcK+sB9cxxUVv48q3h/MBktdG105pCZZXx+ExBxfH+8v
H9iwkt0aCxJ8KX91XECCy4ydFS9gW9sTSB0fs8QkUPEn8UcccwWQz2bObm6OhjZ9
CJvSiSRdnZxyS7T47EMfD/hh4zavzPyqF8Pnt6cUUFGbDOeQyKcRrmwhJpxRhBrP
xLTTyKcvju78KG5HEXmGlKD46GNqtoEND48zE1207G+ZYrZNHDOGN3nk8jzyJ+Ti
Lg3H32EXybRJJ+78euz+WxoXtq0T24c5+dG+iaGu89o51Dqj4tNbwQUbNlQCr0Wa
skvwu8nyZVEbtcHW2Z4dGtrRpwaOS5t3QCRUCJDUN7d69662Q1VCbjsuVd+HDq6y
6lwQNwVm4U5ZS1Qg7TZhnbgJ0ErRWZmHfUjblW+kNgUAQWM5H+GA327V65WJ/Eyz
ZKCFZYAaFzu2iyPbfpMVZ6sfHXX1A9b4yuPrcS07ow8ffxCNLWce1YFQlV5+vKwo
bhZ9WhnQGlEicmspFJr15UES1FnGQuM9kOaAW9JpeLs7dc/CiPND0M604OPKy0sH
fY22QyjmdqJqdDSGFZWD6+xMfA92+J8BCYqRl9IhCrcvnjvjvcZSjiCUZocLom5/
223JhScoEc2UqjpMvBcwnXDkRrxwnNeTp+8dGICnfwJNfrZEqzv9GNatPoHcIRfO
TezVHddVxmTOtLPaiZrZYEEXI/if1/aFuz4LZMtlIFq8LC3DE8SrbrfjUU3cz2HV
Izim9EeI6DZZYsiWgFTRz563GhILwmSvQ1N19Jpk3FPMoaaN1fUzNw/aAnCBCfRs
4rupfG9BhiX2IOAWrGu/Xcuw0IATDIZVR8YtLoIqQwh0tWYcM/NHQ0OUvskEBi95
3YlCvH5xtvWkzNUDjuTVl6fb6DWWVoH1q2xYxgeioV/WPebXRLLdZ9AtZ3WY3F8L
rIzrW3KBrym90UndjFZuiVcxxI7bvEVwPbJY4trtz5IDc2RYoR83I35bkQEpwJtp
mic/S/Qw287DQ5DrSAs2LEqbBpL5W/xc2XlyYo5uSG6IB90VDk2GPC5YtbJuT2ag
IJkWnxjur91PRKL8DxAjcXjOVOZJPiE91VZLw56ofBTAiAJK518u1fC2W+VDrSNq
G1xcR1ArVXSirYUz0vqm6N3iBjP+3DZTi8pnt8BJms3KTLnw8eWk6pKGqukjGrFs
nvUF7IUfx8Erh3QwZwV1BZ4WRZ9Hks4FEFsftmXGFqrLxlFySSixuAZTNSfyxdGM
TlqAczVCbSTIn1nkGBkK+EeDn0q8qqXeghwcOHrggfFMhbX09X9c6q5NLGO4vLlz
0wRCIjDGarUah02UkqIr0TYmrDgpEBA3522OmEhymAO/xgH8wpd2872V5/QwkyK9
EgFvalWIor8lzQCF1xveSWZyyG1SCn+9dyUJ49+eKdZeEpVYue+zd7wQlT5IW7q/
96vH6+fcV0X6HJTdMgc2qYWd6gXlWHBh0K4l9QSFBvHy490oC3yMu7LphHAPrCF+
TByJv0pilpbpiSMG9TgeHvG/a/nnuJUad+NrxpLf+Ke8ep49wTQiSTGN38EPbpz2
erLSnB+gPmePjZEn9vc5inYyL012V/TeZNc9timZnspBuNjmFrllC/Hl+DC6Taf9
fVcz92yQUv9bfkTIvew0U1MdSS4k+kwPyJW0n1pIwjSG1uOmFfyP4p3uG7WjwQWb
uZw5u/ONQMD8WnfXr8mzJVJNPnSRcaaUWQObyjG1b0Z7/hHxUvGEk/L8GWHN+AXO
lkWuIwfb3fCncsKM6H5NsRN/9QOoXxJ0rhXAraXPWwMkrXGYEZbYd4bJD84q/Gl0
VcuWcnOTQmTxh3WGfUYc6dy7GdJvltRANou8/eTjb6ProSYhlsqA+B8SC2COoKSx
2GSzk38kQm9DXKNrnWS3CuSTPHxyYmBs6lRN4O0ZXHlRfQrT2XH7PhqDqLrw8bnO
xTRRzRqGxIqpZUsJ/UzkdGNtTXELUj1ET9YjYgH/o2K62CodoLrPp3rIW7gVcEJo
9J/E522eDeECqxkOaYiNOmaGFpfHlUgOW1554oP4kWlfsCnGEqnTI08gG6UVLepQ
rQl/51Xd28tTDvj3p4LlRzoCkl3t+QmnhYovI+v9sUPcbuCMB2HrZ/NoQHDRFxCG
ahKBxxYOuGW8Q9MhIlxnDsaKx0TRd7Bx5Ijm6Rf8jxmkxfBLrTJ2OPoXXflCU6T1
N6b+1QaRIEjBzRjwgAgA5l/GNxn8cGwFuTGmLd9opmunZB5AodTLbB+TjCXs9Qvd
IxrdK9929QZd1+uHhvqTZeYEeTZ3pVZnut8fXQ3FfYwKFRzDiBtpZYmsN5Tw0PB9
V1OGxXVpp4dZTieGeXEx310IQgb0ugCVvvArdNYlcKZVGYLkIZjoWZtM3m0r1hSI
b3nEVUusmgi97dtc4YuCUj862XgsQUa0rCTjCAbeJYkZkCGfMVetYzoZs3KdDinT
rM6poBTeow562GeKQlLPsY9TkvKo5uwvOXv28zeWnZ3UZozK8nvLZz2R3fAkABTe
1QVJdU5i4pGk87PcLpQvtC5fNSf/R21RLjt7vPcFr96+URLcj5dgy+9LHWznJooW
5uskr5nKXNe+7nWWHv1cSiAFz0SotG90Oi4hBuc3dBU5lEIzEYMoJqfcyoVLVZs/
NATxK5M0ASQdMnhbwEhULZhKZ/rG1aEr6NWyRK9hB6lAuDTBh+68qfcsu32rRrbU
luQDlr9Q5lN6iwxCkW3ezhlsmVZnn9IUWQgJsAzX33SwzZz2rM+kbiIVU7AfMnfd
78vTWrKLS2+B5dAE81wIPn8DnLVXD/hVtHwlLSvdcxj6SH2OFYw7eri1AakELFL0
+MvuUNCTtLS8nYarmCnKO7GG0X8txIqFG6J3NcXVtvt3bmiZGMhptXZAzDcjR3Zn
Kz+qmoGiMkb1dWEDj8s93Of2r49TBvPawc9ep4yIXbvjjE5qBEL76EZ1Q3UcDdYk
EipPxaP79XQZ4x6GzidH75n3lMqe2LPkvFe1qsgVNyvT1WxbekhehE0I08xG3RKQ
t1uxGV+JAxjtVSGaJ4nd107Y+IP5R8vEVG7mmyPAzXKMUPknB7fYtRyru/yyUo5g
gobDHAyMN+jLOn/xjVSux/ZpBBcHx09EpdMzOuQV8Yp1u/kJjsMv3363udhf0nlg
z+y0ms32yAeNuOcP8VK4oPJbxhzJG8DCi8wfzA3Rw00+bvThU1cPLPQAr+dqrUSM
fVMZL1PK41A7451WqojtS521D4sH32Raq+7y4ybrjZGCZ8Yr5M983qFXBKJ4Nzin
ryjOX93doNQzJKNaTjgBBqmo/2a/8JRNiLx2F6UE3Bljvb/bRb9L9mKJKQb/f+Wv
UzXmRvrsifRrYS/ggh047df0QsjE1oCdC7EvIIvh4ycO6NLqK5CbcC9PIwKB34b6
N0TTRdzHB1TyIg29ITar9Ow0Gsot0LjE8AvEel3kz+AKJ1O+okjB/YMR3jETw4dy
dmrKR69XByHV8utDBR3i1wYo+dAlwojQGW14khrtj07eGGZX7dz/WtLueA9KQ+cJ
rnJk1UbMgoJA3iCoQVER2rPJuKZPmXqu1aD14w7ZhGW1shTA79RcBYIkrcM5ioc4
JN70YopiQF40IP1TfFTxCRC0mkzwp/F17wyv7y9DbJXZYh50YkUkw74hm95LlJNu
gcpEJyOQkZBM4scHTIiuGxQhlpPkI1ah8hd1jDVyMz+OmWJsUNunXmIIOgyPcFwP
qqeq1JBGZ8vJb7TOCr0LfzIDa87KQ1+ttT4JEVuMwJEIFom8wGP0+JvPpJPu05lp
jHU6Hzu4ZH1gDeDKLN+QsfzDplkldMqxGjCuQWofyWCh9460raeKCM4yNJ98EaY4
pTZChRJBqMlY//DmXjOnwpWww97xT3UA3LynFqHNqqODzqUVBemwWqe7kc0iO08V
7JToWj7mzKRlGJyDK/ondhPgGgP8argsF8bg2m/kNQfC1ZSbtNe0CYB36Y3tZfjg
yzwweB/gj9kvkfmvkGCTeuEH2orCRdPIPDmfpBkqRJzfcEBTOszXACzScJnSzoGj
wZ3qfLfowWWWnpYSf+uiWjTtJjp02G6LDjgkVSVeYCwu1CG/3DKrApNFad0zcnWN
P8pTi7/AmdsqwKFZs7llx7FDt6K35+g9KIDMAqZrEG+gnR3aEw+a249b4Cg2x24C
BPzRAVRDc1BF9f/kETi0UydeO3wAmU2w2QZ0COncN05uIlaXzKjvQoGG1ZB+/G8r
gJZnaNngwtAYxb81psEu28NscEsV+cb2JAGYDgGJrFSB8UA2qAHc/1XAo3CPRHSG
RpsIT6Op3zo+q4z4G7qHhHSuLTQ8UbPXS/boKU2H6JTCl0gWNc24UkvQ3VZZIWuO
uibftmidl8n147L2et2EQ8qRAzfwsVsNXFxlI6KhytLOnMuLCWrseROBkRb1O4dq
mtXl49gFK3xdhVS25Xu2m9l/j5+RbzblIbJJWlbMbpnPfUha/eT7Rqj0xqQTuzI5
4oymYptlkxXtXQ+c6hmSGP9uGYb6HmTXBStD42nmWL8/l76UNFT1oLdPT8TCFwPm
ClyajtuR4TC63W7i+isxfZs6Z2lt40Kxwws1R3I13RkqMDtSabKM61ImW5I2Whkw
Y2ZREyv/V5QDKdFO0LYkwnPRNKoW0hkaadiLniWU5e3jMgcj8PgWRtdnFp38AWQs
mNLoCtRAi5FHtMwPPlvST4lvw482XiQ0ysGYVejulpApjJZYnNdS5VONdsEVkAtZ
44brFkfmoKkYM/Tpg95laX2BH2b5xFlQ0tgcpoGQMuybYED6awYNn7n7jF5TwBPM
VHInWNFJ+3EMHTF4Uz28R4rLXlmcSHlvFVwZaF9zIxbgQukS0XGq1f5cF1y5zq5H
c1OOotPgszqLPBLZIzZS1H5fhhuyMaFPgFpuE7o8dkJak8bYfT8+G191D767Nzl5
JQpYOm/v1ykaCVaPMWYCJJzQOiYEJS2H82NLEj9ugVmuiTodoEmF99qHLw/0w48X
q4zYnTK8HGbd2ukY8fO22dNSCzDcwie+/7yo+INCgc92if+i1mR0SSJqpytToVXK
XQ1x5h9ccn9dRJ4moBuvPCQMIvV5kro0tlsBe5TiF/LSSnzY1HoRwpqxxxm3MSkI
tm4QlY/D5Hh71nKJV6T7qAYswApdeQp26K1EqYk34lPQ3oyYhAW3/FT+9ehPz7nt
Pzi8LFzFi9AW0DsvO/OUExmLb4UV0dqL0PWVxNm8M8kojY2D1CBilHiruBcX8PXy
gLEGnGDYca+MBWqKc9CDa8U4MhWJg+34M/BFJPpZUDXPJxzYxeqlWdPctlX9AtLV
mJL9Is63V6HXNNU3Dz3PoL5hpyBd4YYtlSSTyWzREsL45jplvW2bxUD3NAp0q6xd
71zm7mckmtThZ6vUGgA+balyXm6ihQ+O1Ag+nDhwLlQzS5K3CwxTISR3Y3/5UCH7
dQv01fSuOjsrGuYEaQrEW6Qk+p2u4SNtuMPhMsWxQOsA/3SMMjKJvObbj16Fy9XA
GUHjZQiR9gAW3rhpINae5wVGjq238lVlMlzWLOeDiPU9V/Om8PDsdTcRhtT3Q37k
Ri7rAcczTUkA9AdacbEYHfWwnA6yYuclxXGZEePsV1vM1JgAUb2HkBXuhBV/amWs
786ns/B5Z6/zGM+WUyBt6evyzpUo3sFkofr+JhRKZC7ehTqI2VKk8FBojztf0Efs
CFxtcxaxjtF+DuqFVTNRGmFNni1meWzb4fNh5Djl4akJLNLGI18X5sO3mWkLjuN4
TUl4suQ9fc2X1VL57UoBgxZASZTRe5333hV8MxUH2ZHwTdxHDxWO4cGD4oGl0Isg
bC2INEwu3m+igCW6oyBZxSnWDPXEPnq+XbsCutJdPZT4cJG/BrtI1hJU0sZYvCJk
5mt5+3byerPvKLXNFj2k6fEFqMAEzq0OXOdjuK+D3F0UQ1m7IETDd/EHAzBMrwpi
J2qv5nVij7Vqr6bMDvzL8CykzBGYXWaxBYmT5j/nufliycM7OtWuThGI0c7m9xFv
oJMjALMa8bOVSWKTcdx7JLmvLtsN5xLlIdNT7VbGFRotsTlHKphWFxV9CNtiAIhv
PWHWa0eiaYh4TKurfmQN0MRxA2jI8JIgEHUZjdwHMyNpGMQhvNCkFf6YB5m3eEol
3fM1eax5oySLzJbephUizBt1H1TORoD57+aFEX0Ahg+bSipf+rWuqbn/kKxKGTtF
fXLBryKdfb+CnNsinujZwJOQJ54WT8ponW02ocvxUb9JDbCOIeA2a6mX361GohHY
d8/OYBD27+NfIoa7g31I7Pq5bypCNoWiGvGuvFq84hDUECVDfcXrnDgsSkfMU0gd
0K6LGlb4L5pn9M9JeEmLn5YpQYHHt5hl6+6XF1O+PFCEUQculLypej1RAGJTPdWU
pi8OqyGX4ELOaOd3m21864RLHGBWLQD0or5VoqI448RkTvZdvRvdrWi5cN2chsPP
yd2Rk9qoxOll/ifV+crSENJXLVca1lwPoDne746ga59MwJU+OW5w7DEIcwsF8LBo
pjxSoFgI30weB5z/w8I15o+iJQ2TqkTTottJncd/Dz6QyLKJVWdLCGXuI3d1k7kc
+uaDujNMFvWX72gTKEa4pXcqBtlRTSK4WiFN+gGzRRlr4K2WKG7eHyIfdZ7KRMq/
nJ/Q2nf1Olp5eMIH1MnIrtu1UeCErNDUPDOmPV20X3sqRphxTzalfA1aL1ps758C
cN1O5ARybfse64LTnd0Ge/omXqOU3ec0e5uzb+exl+AuJtt+7saXRljcynf8tV8w
SQwMuA0sTuALKGCEzQKFEtRgqx8bcpBT3NHY/ZQ8FNogrgrIV3PxSe7YwV1kj+KC
VqPLTUNuO8g7PP9klIgNrjAY+xWyTYLejEQVSK+3CqZqNNmCtZdcDQ2FBcJBgY3W
RCJJBcdxXocQ3ZLzvlONIyuMaaeocM7w7zTiSjcIMTRURRPuxtgrtaAhAwsnQv8B
p0i/RjUScM+y+WyJUGmsxG4iB5UBK7I0cRAGrSDkoItvoTAB4ntfvq3tXXiPJxyY
1TdTOMPe0N9sS2+W7sROwfVYB8oiWZmjhx8ntGoPNIzI9gyzjZ5pfae4pbXbk1KI
/b4lz4kZAeIWW0quAJkZDfgTRmVOkggQuWwcti5dmLICgk5CGjsmtPQPp5FO8jF5
8yK+QkNNxzkNDB2BA/AD81kX32qJ9PS8Q0C4ME0iMTlLXfg6Y0nLid4KTQtIqV30
V2q6AhGUhDtK7ZQ0Eyaqwq8qR35qB2GosrK5Z//acqPUkNepLC78brcXsl2ExJ2+
zG+YH43NEQCDnheQAMOt9WpdUfmibwrqnBqygaO7azOes6KV0uahMbFzvrPzhg+z
+3GA9k0RD7S/ZwTeLaNTsVA6WdO7n3FBwNmiLJFyFQiVZg0fHq91ojudRiMtxVDW
5gPYyMSS4Mx9A1Zzjycw2GKC+icwwsH8Yh8MKhr3jy0TFoisYbThOrijWJap36tj
1tsN8wHL093C6T7IJ8duUGkehNys9vtPfwipoCDbDshspheIFkZCii/tKk/X9pDZ
kkTvFv/hS4VFEAGi/cykjXf5ZtGZOHJ5pSL1XKOeIpSUoXsus3ZfPfipE/4fQAdD
GW6kk+7Q50rxynUXOQhx2Iu/VRjqwUAHOHZ9QZSa65UN6hzW0J4yy+1ezwFex7AH
RTD2or0QZCan/nAC8vSLEs5sRgRNgs5gemdk1cKZKnymz1KHc/fV/WOlMh/ZK1P5
/6zjG8/mZCF/PvBZSF/q+wVa4FRXup4L8HYsHTcvZbV26DhmDW8IN6BU7Qq/t8Xq
SttB1F2XgjHvfSXAETG+BTYO/bfflFnrsPlfzwseL7JC/DvB1ZJyl3UByCCht0ry
ELr5pCoDuKjGkLOU1KPYIQdcIEKUNw36IKXzgQCRoRKA/hT3zPUxk38k4bCRnc47
7aImiP0c0rwEXqvTdNvhcslqHigm9Nke9EvpUKdspVfvEx9cxw3Nlw8bVBlkREoH
xUga+fGSl20drsig7FZCdJTPxq3fQS1flBEoSl13RfUKTrj/IitcwNcQROqgws5Q
A797FFzdGBkBIKetLn5F2l7ev8htZTVbTGvYFqcuPQhSPsp6Ui8ZVZazuV/6KaGE
C01TDl9DiZ09z6q/X/idf1eAY955tNZmhkSPRCOZ5qL/zOUeWTZW9FlFqdgXowKS
XHFTv6kIYZrn0DNnOZym+lv0m87EN3CWTCAffIIMIPmXwukK6IFw1apbGh2NOgRr
7J79pYSg+kjVbXWTbKOjQz38MXmamC2Hes6ae6l5L+AJjSbpcWkEj2YcXJ9W4N5Q
ArQtXiyNv+OVijomedgmipU5MWE58faSQnZXTiZNQiySfD3aBGdcEzJMFDv+n998
rx8L5m5iwlmyLddNoexYkvlF8CrbS+frFhVzl0VS2H4kj0PYrgYxHRBi6zJC1ngS
U9xNEaH8EMXyE9BnFE9DUK78QlL9FGf+m6xUVXxQbwmJEp0wCMlFjut3z2dnz65j
RIbOZzbx403B7if2LIGjvs9yyVJC/vnbU5oAjF5H9/x6w5ZMC4s3d9bVjTrMSqLU
2wRobVX3HOOO772tMXhvlP9aM9IN19hBd4B3AC2Yyzqh/BHzXuBDglCXoasP9kgs
QxXSa4tC0JpL6EhHBwRjQybuvNucNDge13+tDhYXxYA/Vc2+l2dTYgoUwhmxeQAc
yoB0rm+7B3g990D6YHTwJzqM0AiTK3oFNvQNMUSD/hBsQ9aDR/HqrgXKtRnIl6p6
NSqMeqo3pY6xVPGeVSDO5dPVuWPFjePQ0NtIYEgysJK3b5O13NBMzlRCJJH0hTmC
hy5F6c5H7qwkNo5ganGR8u12LGlX8QR+QrEjLZ9EIxqjCW8BXTBROxFfUNlEY6Xw
Ic/u2eevmRMaPFdLJy009+eQVz5rfdXrcyziSh0jcvro29jfYVmoXpDBycP6nD36
yru8lNzzwOp+b5wirMz111z2fBpT0FsfQB9ySNk8bxX8ddGw7FsfAmhhaY7hk9ew
5Wn7ej8tl7jTKtzVE/kcW+8qcyFtlAu+jd0p682oxKOpi2kpOAXexTA7mKv1oLw8
X0bTCM2Tm0vPcyX2sAv7R9r4bYPf8z6/CD3MJJy97mR8zLeVrt1VkhSbU4mWVvbT
ao+L53PQTMaH+fGs59jCnFGvvzoBNq0DNx9qj+CJv6zc+PQfTQLP5Z9vN6LAD2nF
K0dXp/oK7oRLsmmAg9znXNJXbIG8q1LeTF9dLKW0dPM2fqoyxcIg19Eu3MAiJeF+
x1u+Vqy26GLwUQ6/gIKoU3ylpiqvwwoZENoclzxL4waTlblxV44e/KQgzezVSPEO
j39slSGKBu/6XVQexPlEsgppYvC2VpMC0k47pQ1hF97HQujqQdeB3cfHHlUAM0Vh
nLsVme/sTXF5e0P5VGIlpsqVQnzR14F0KE5HWkQ6hw2XfwyumnVg6op8S4+KRu/K
itgD5CZqbvJIc9EYAVVVKAjxYsHT8AwTW+TlFtLiXGUjWsZDDOFrnz2/RphRjxF4
k/+Cj9Fs2n2Ry8PLKjU4YP3jXgXX1uZ4UwBpTAr/OqfwAyjd+V81CH609R1ICv5N
F6pb+hlyuPmpgePyBAzsChqVUpSKBLWDIvG3SB+IzkFxzTnhKCcHz89U15hkOlmB
E3zhPlk9Dt6TRWyGLaPTLXAOJ6THy+IlAb676kNrkzIW7AbHsFvZ4CzLk4kqNbsD
S/JHRu+MuK3UBZm0guL3LhNXgKa/GzWrzqr1jVFYEUqsPYlm9+LaOsW9iMLZil9J
4KkTQSMXOqhT/kQ7AW47OL3L2gwalXDI94LNdSwnyYsNtymm2fcsYO752KyJJxYw
+uzozPQz9eeEjFAvfCZmCsl5bHpujgpAko8yAhL7e/Zkwuvp6QEav5EUAh6u9Cql
9OO8PZ/4UcOcqDvfr0WZ0InxUZvALAOpjXhSZtp1O3VijwmWDFqod8YnRxsYAYMs
gcMNrQbkquAmo3BAgcisWUfKBBifPZXxLGLD7N5/6B2JmoP6l9J6b7iC82Qeuogx
f/vcrE+dPTSf4c78yj/5iaz5i64hSwBSwrO8INeKq1/l6cSC0eqRsEZdEOKsb0XX
KdXane/14D5J1Wd5iPoZoaTnj7NtGPsfGYAvG+NVBb+PadRygw0M1l3AuxNjiUDh
dnYvM0ohs1ycEjkOtwkIH2wzkwL8SOLUZvKS9OzgeZbZj3Bgt5qTyNG3/1QYVvBq
r503sEl1yH4IUM+bCyL4OEJlQibQIoOIDciVlYPhjl/XPZmLrbzJ7ZSaR0dh8zpa
u8dKT5tZmKNR6KJKlywn6/I3Xh42RE7zFN/zUOF1HC7yBrN8DTLR3RzwPyfWuiCf
Ybt4OjIbykL7f/6zvOlOX6K9LQUCoeFM00+bASJVTYLO1RCo39bqEO2R5OhOea+p
1iySW7IaBwARdfFGTwMAJVnJqohiA+y9X6ZKRohHWDM+/Roc/VZJccU5w+jUT9X1
/9NxSA34PXGbUnSw57+mX402oR10v4dKdTX6hmVqjM1PLy3KyDsKevo7koqrNG8h
Wk2qq7tvQLkBCNbYM2rV75gus8UWSw8xsbW1j4ZxsgV4fjeGZyhSAHK4AYCnrxYR
9k7FPMkx0jNqhgcmfLuN4XOwKzUVta/+Bzc3TrO0aZCTFAa9jmXccWK59ymQdP7Q
lFEqXzlbD1YA0jyYNc8AL2ST/PW4xAAt1P2pF6Jl4ISmgDJ49IFqz2KjmGYmDjDg
/94GR8tbX5Wjv9wBzBcln450XO8rfIYQLUcwGME8MTvnGrV5gM1rD9ZLGX1mJMrJ
14JFEsdFAnhgGL5HONmQhKyjo5gJfd+oE5ricNFpWrF1Zko1Cz6HeGk5ssLuPufo
IUW4wPGyM2pPeeUn2oZn4MB0btAQ5grDnlBBuEwfK9x3ah51UNGjVG1aiBMBIkKk
syff5kPcBew3dG5+LramL0WAxnnu1NbFH5n/JdiJAewSMnRoRWJbGrF8aJykm2U6
41QqmgUhNtbgjCxl2wb/AsOJeJ0OBuBe7c2xoFY8zAiRVTeArqqKj0BigdHYjDJL
KM7qHPZ8XpNFiWY6M7BvEQQq+VVtIWi+8YWal0S1YRjmh/toYtNjD4iaSL7sn3f2
/C5CBiYylR8/0o3rBBG+/6cOPt/SHSK9caZokIJy53YYAIR5qUYHEBZyTs0lw1Le
+BhfB70M0M7AIbebSdMuuLyXGEBIRgfDnnnjgEKygObHGU/Vj90KizwwsXOmvHeC
OIhdS14Mj7obrdBZyiNJiDYweUvSyER+PjLRIa32fEc91ARCAWh6BfvbSoAueIOg
1889RgIjJcVt+LzmweY4pTRI5aSpQCLu+dG683Hs+/cCxUY9I6WykaTL+Y4qu8GW
rp5amq3ZaVcOsGlFhteLCtkGwxa5qPgv18MDvmRezAHaSC/lC3rRrSfmN7t6Tc3w
UE0gi5cFvSZ5g+Ktxc1W81nn1tp4EdF6A1jrCp1l6RnhoTITBY+V2E+XeQCPgLho
bA2pzwszFe6opGchDv9Gd3RPuHiq7DSwmrQxqyMNYz+nuCIDyu60tZbhGJ8AmGea
ew/3OtUSOh3ltnXgUR1UYDzowd/k87FWhnGDspNwE6rA34eR00u8U2Xiurjno6HF
N0FWKg/JZxgw6eunSbc2iY+GhCBo5kQALHadHAU9W/oM2Dy5mBoYHpK7zNhhKZMu
YF/i3rGo6YoCKemi6vgYmF8I3OBOPxo8E/sPU1inFeA0aTSIvRYpgzhWIIiKTbrt
dYy9P3W68iyONd9UFrURI9vVwwn2BHLTSoj+7wpBYsbX5qV7y3JWYSLTSnIQTZbI
bllqiJRVsSfRqQr+Pub+XCO+3w5mCbJJchjC6H+MBUgB9ej1F7t5PFUl727d6F68
WGErt4pttBnJk5wmkjglx0jnLbHE8RK4z6Lb6OWIoxCbAjFepaZgGbSWTWlXDGmt
r9Wy100vJLQ9fY4WEs9sPYfFVzcEaZ0l22btsdiBHWgxfIHTPtQgfG528/oZcFzH
HaOrlbBvqdSu3AJvbahUHlBU6xaAHbC/8VSxnP/eBuJOEV9Efl4MH5fa9OkgQrW5
lWAZ+K6fEncvAF0Z9tSANTUXyWh/b/EYPXC0DYjTPbelTDh6OH2hAY7HFon8PjtH
KmX61gdwX9Iu3Xh6lbsLUshUSFl1tpb/YQmS8nI/Dm+Ra/8kxTToxsSixSklDFaW
+94ckwxgdGBOmjajPRCSLnXugrIxzOL7eqRoZJ/s56q5j1sehrUCL/Ug/MldPGPV
ZrB1TaA0iAgfFWdPSKPwkbH8twKDxuIQQ+K8XJPaIOeoAeoS8uYbDRugrOn+Xbd3
ahL9POahV6ET6xhCzZ/DCFiWMvf1rjCIOKmYgGIwgv9pjYYhdBLmgHx7m5yl3XKa
yVd99/06bE1rviqx2X9fT4OkF+IPhxqGKpA0afHQdjYUd58ur/yENrzutLit8aM7
vVx1AXWKAjhfUXaCp4y4QN9eBeMO5ztVq+jchzZKPOAAdUOywYbNG0PLmDFpDfow
Oihmj5l02z84RwEFIcYrz8X2dUFqajcRBfYNeuVOKYD4xvngGYSy9Yxl/YKKB0TY
ZNn5RHW6J6Rn+rpD3CIrFaToj5MQeaHQoSx7JWV5nDP7YZ6g3OPXcqKkTVoLastK
FZaL2ItMhfz4aWPa/c9PkW2p28Q0pjbmyimSrvfnQYxpfJ9rk/ev55fUcuVDYXj3
uMi5FCU3G1mYLOyHgggtumdP4MiLpBeqBkQ7MFcVurFlHQnVCIugv/sSmYD7lzLq
sYBVpPeLt0qVh6I2RR2pAYYZ6/skJ/FtmvECleK5QiTm1PnhYGED7btCa4EdZYur
OgYUZXK85t5GP8HCuFqMceoP2//wcF6+c/qOQQLCjcreyvMfpQc/O1AJl52QQ9Wp
pDYIt5BVLdT9mMsNYBXQa9lUpjyWmjnuN1BvLtsBdpIiQK24xin9FWjVc8qEFJ4Y
qgL81STfQ8rA9DjFuPLP+0T+G5b/9Sc7aZ2hxSRUjYI8J0vGt9Q9jfMXpvTC8oV2
ftnykYi3fA0fyFJAa//T94o71JgvXB8Utz3XRfpV4YzCAjN7tnva6Vj2mD4I4c6I
a+6zatbyHez2uJQLoTpy5+oHMKVZuAJETfqyZLr8eBYicQFtffNLvNEZLYayBwFH
TdzLmcG0gp7fhx+RKfuuz1967J70u7rtEl7BZyKo21b10v4AP+vjIFMJaHTErNIC
wJv/Jxq9YvMbPbQgxp/HyUxyXu7NH9go1Q1LpZ1DOMb4NKdUXz89BloheAiy9fBD
QytsIAfhh15AtdQ5G3OMA1WOx20EsaNiYXebt2BIsOBEvJfKmEPevpt6QZ6rV4/p
ffC4EqffjGh6yc/vXUV+IAzKYLk2FDe/KgrvUCDerc5+gGdJEixqEWNsma/LDa4y
VGwh5jjFI/bC/pD5+BSqnfpDtyl5wi75VCkbmwb35BmbNZAd3LNVpsrDBJzn3iFa
ypcTK7DlibybkRN77jDscY3fzG7knVgOmWcM5awHyLZQCmPJcnaMsRdEXxNhsVQM
2tOiyMNweV6dsnltDAX6vFpzvhHzy4duzGm2TTm50N9EnZGBTG+n88qGF2Lc09OL
XEbT7Bz8Xz6L2Q0MyKClHswdwAaz9Kj9EmE5gtoW/Z7y4fiv8YbA7yU6yFTVMXET
9RtjfccQTtyL8HoH2MHu+0QGAAXjbL5T88BycJ+foUyPbFlsGqmorgV4U2jQior7
GHsU2LJGW2IeP5uekoSL0lp329SQfAWWLXIIBY++xROhX+gbNcN3LtANmHtniiX0
WBgrSKOsUBX/4CNZuln4mMv3DVwGfeSfHxPnOww0O290Bp3SqhTsjEyQcbnyWdJu
NRlKqeqDCD3Ckq5Tj06DDlq+EVksrOS96cErUb6J9xzikQucFoEpvj/aSnLH1Yzk
NY7T0G0xoAe9UR93u6ZIiDgYPkvYTOvhQGIsh3IT23Nr8luEgBCogGOupc2sm7j6
VPXTWNJ0jfjB77Uv896KPHaeeKbehJ+P1GU5f8yJIXCRdaZzQGhiBOpLJe0E4GTm
Y+tydcEsWa+6PHuFaHYL9z3O4d1qlRV1y8WL6HnHuYyR/lt60wYTwomJhwZUrusu
j/rsljmezAkfTHVQxBI9yDi7q9Rea40iOopF7M9C7aYAEEDKiK/K7WX5qM68Bsnp
FdG1lHp8oJClyoE4jI/bazi85cGVKOFUAyp8VFgmGd8euNutt/v1YKNt0xiAkFQG
wLhseTkw2SU9eZlYPbxfRMJH3vzAHNALbeVQOkIGx6ZoBT/wDaIZOkHecg5+RRS8
7QmSxoi5gOivuUyGt3XXpvw+xttWjlRSZZaXYcFeehlobdUGr7amXZm3DulccF4K
+GQr5ke5cLFnNfpCwCsZ+w7L3OyfskSzNhQTOh94nlTudaqfkrQHymVF1/WSFnF4
mln5ZFre71mgMRAw31fnE3itka7HYauFAE2AyLgJ/XOni0OegvDDGEnh6mMuZ0Qi
PajNtK/pPPPVhhnL5oKnldUNG5N+a/fBlwKrKW0Nhdq1VGlNecy7ug15xf+Kt7nN
Mq2D6Ysp521N8uYmaNi+Zn5vjKmzPUe0gdwQyxZ6XJMeVhRMYVmU67DaGLi84qIH
7MqPPRcXpAfkYZQ+kclT8W5MDyun1Xb04jfEBqS8OViX2ygV1rNNCpjM84EFSsLx
O3IKbB2YOJfD4QbgHq7n7Mg7AAEXiLUlaOV9mSCx4sxLsNRKcODJwxLymRMVG7nv
RatnwXqmVxCoESv/+Z4VFmMHCLJVg5mxmr4GqU1VzqFMkwDyZjZtEKAE0SDt1WEg
XUTZAX+ExvLRJKCr8Ic6GywzDEXYNE43VfSdLXF51zXdRe7bRoyccj0iAkjdpE8C
E4IgqSKS3O5fBXyZOAUPH34OEX0EF/UcE+tQppqXXvS4eTBf46wiRBOcFFEqBVPG
6ognDcatXCYcvrMaxDfqpTafoZLaS28lini95ol4ypSeawa7xtAB0BavLCnVwSov
psYozopBezTkPHEmCtlTYVfUIw853n2tgi5f3MrwjhMvtldA8vJ/lRe/PwyNK/By
GUaldrVHWoNMTC3ejn5u1uAZ6c9IJDjUGFIy4H5zYwWWtZb3GqLspuoIiD1hko1x
Urypu/0EicW4kbV73/tLPlNn2ERZcAwx0io1/UMlQ+mgWk+vCDEwTpqpumZWG3cy
WDezsHQglbPGHE4Fp91gNqFc659WOtIzSnLKXCoqezIBJC4VCfJm0gvlODm/snIB
d+sgKFJ5NxxoMshGdCsSSTQDu6aOMzvcNu6e5eo8umf7FbikcjGaSyRybDl5Lofa
Y9c11b+JdlLgJE8+qDp1Q2soPsN1XabClCTS9glxQX1psQWx5UdhpipvBUHvzBFN
/+MwC8mvOtPTZ/EyqS82T2gDAiMQwFhWLADHaUcB78f++sXlY+Ws2gKfztCrfLkG
ggjUFt74biWfd/1jZvV5sG+bL88D28y2h3FrdPe30eOXIE+mPHra7hd6MwTHZOYV
ujigpjnzGLYwJ69MIH5ZTHxFRWjPc9ZMtBpf6gkWuRt6jMoJpePPSBbrFDMk0I5V
aH66W0lfISDJPGTQGnavf9hPdHtjHK4oH7AC1Zkwwfd3ivOkfXjxkORDPfpi/eaX
EDaXVtpH9ZegTN8KwYeYSfddd7ITDopj1vBrvuhY5NfbX6UYaOmaoRKSzLNJXa9x
RHOqsH3ihx4jC6OMNXSFWxIaWrivzeALt3K+bKAP/rXcSNJb/42wxW9sVDqTqTAg
D8mL88lVKSw/q+dCrL3mHY/12BXJ3H/hKj+WSaam0pnP2hZ1ldOF8dPPTNIXId4K
uR3/sneOoDiKbu/YIPhHCc3An0FJpbg2VNumRIBmjR8RLKUWcQlhf26VXxEsnzP6
bSL6ABzSVF1uujEOc0/+Q0fXvob2RiflzpKAIICLG1U8pitspB3+l/nu3aZyOqN2
zDaXPLpIP9GRC8GmyPR0RWOVn2589P1Fd+lG/hfsBggwlRWeER4oVMzm8UN+0ChO
K8R0yeTkFcflCYmiP9i8a/y9Xho399d1flV7GqundsFajerLIBO2ZkCsY0FvPlmQ
OjYdrXJW/i/og0mkysK0x59osdafFZG5i5lFTGMWYWwWBKzj9Y7s2v0UsU6SsEse
dfonudGNLwPZYOnThkhDpuH0tw08cIr8hY0ROKBROQsUMx5TLAjfovy3eFDgpBQi
qQs437Dy188nCUmvCBgBvFu/3A1fmR8gNbYrMEfw0w8Ro2yInCz+li5cT2pymlAB
CPNC3sWwPrUrgzhfJac+4Wzdq+3IqNxqcggzi43iHqMT8vfyId/uAIG9rtYWwkEw
/0twDhhUpbrF/D+DC8KEnvFWqILhbCAwbra33uhCPzvucdNAFmoH+sOBDpc4Ahg0
UfbEO5Gt+2Mu6+EX99KO34F4UQvvGw62GHSR/ENRrCV20gYWmXo/ddpUJFtOwHsM
wVy77WscDwTOyQozV2qeYtMRZPjkoTwE0e3JKmdzI36aK0QY72RTV2/SG9rUVE+e
Cr/BZI36TDa8SV4kszQXUsJwqkx1m1cVPub5c/4UHA1B6ay26mEShJawYplbor94
yXZ9PEEYQgP846P9jkYN/kumfjKh+NDL4N3hH+UdE/56OeVeB9Kr/eN3+eRZ0gke
RETUQiflKKxYqOrUerZs7HZZ343Y8W7jg7ohLgqWEfjRr8Asvol8JmAAcnQVXGzv
H38aFQ5VXZOjFB1hI/kh+fX1ZxF9ts8plAmtz9ScnvQTE6rOUGD8dkWDvA5IryGL
n4FSci7f4kWcL9A0uEa7LHeN5DunVTzXL4ZiornMKtdJxuWN0GSfU2GUH60Y0yPe
GK033b6LuQZD/LMUyTde3GQtIJKUf0S2hel4ABBqj+zVlFRnSRzIFIsrwOnlwDtU
7p9AE8QI/Ey52+M45B/Hs6zWhzGIpKB7Q52vrYbYj7pK4OI7HHWpS1YC2quGIuaF
XhwZdwDbYjTf6WYmVht3rtD0L7K5moaEKarxTOxpgs6QiW7aWQWOMVJPUQZcbrhS
NJpFeI/PJFP+CHQcjf1fwIzYJztTN4WPhh/Gt5Hp1JKsxeOsBNNQWzb8TuWQx9tA
0O6dT2z1TS7euLWrrRpG8R22R79VHxVosibZoQrZnU0UL2VHR5BLaC3xflyFy4Kj
4zLJBbRJk3035AfzfPqSpbw9JKSigQuMvos4uUIdSM4YVa12BJ7KCqab9uX+fkFX
ak7CLkw6AK2Re432wu4gYUHvZlnMlVEUV6rXByTQy+LpIHXEYqoFU6UelPK2fy+l
Sj+EAypqXSzkRZ5cGN/PwPpbD8N/+ehDkHUe8hC5FCux3nZ8oWsOMMiRKSQK/V9P
ftJhbvcwcVzXeGiRLowxbXD5xIZCeoVVpjcCIpMFkd+8rHn4WRqqbhoo56Xsru1T
K8jo+MA9zcRPOMGTql8GpeMvsdt867WM7R3Q8oSUoE02rKe+Z4i8o2JndenIGzBc
kdmXG6XY+DHSN0hXyiahV1gpZTOo/zBrFxoi1WjwJiXoHawdtwCahMhEpYWsmuiM
XOVvz4szh/9ep1nA12yZfCEBzQcW6gFMPHRFxiSOgZBUblHOUGKzGF59eDIbPwpY
TjCFKMCVIQv98nn7dPEiE1WKotjX7umPwGAl15Y/3JCmAyMhpaaWIrwVs3geSCM4
hc6AwQP0fXe9nfkRcsbPVAvQzXN7Wi6VVe2SCw/CDM4Rpb4MokSt4CRlwrwebq6z
1toU3jWUdp1lX0aLtNc4YGqt0D30zNDZbheFdN7GrWikBdGPtclIMlc5guTcHT4A
i2Spa4oDfdgyIb0UFVLZmJHu0xEyNV8XMN+GvYWn4kO+X43P32U0UYSgSl2vnLvB
qAKLWqhyeWVMgbcBsdHVfo1yI5rpf5V57in4pPIBjHKQvlx6bzQHpPLExWqlz/H/
v2mUl2fXsF2aYebT3oDqg+JgHNRFE56NqFT08/4yPvJUryyqzqXZ2925ecm5uY2K
spahCXLhRtjzwaAux/e+N9WjUOgFwKdlkoKpcAocqNcY2ZaobYR+rUbC3jV9m1Po
tGp647NMa64BdrJ5MasITGKJti6P4kiK4WnSyxzSVze1Zx+7c3iGR/G2xwo4f8Jn
0Wx+smjekqXvhrCD9yU4yNm9kcSMJq15UV3TY8DU+snPodAF7rkzqnCqX+JKPMeF
Fd2NZ2eutxhfijhaJw+c5+3W3Uezncryja7SZpJDLssnl26CZ8qd4ui8R1ftk0ys
N8HAT8qFvY1l8FghkQ4NaRq9xJAFyyNd/juvoXnDfVI3N+pcLzsXXJLKzmK4QAZ9
Hur4Ax0jGsIsFh4aDbn9izURsA9j1QFcbi/+tZhHY9jbguTtPwCW7sl8w+U+RDf6
oGB7oqAoNdXxnhyotOfMdqFbkhuljovS8Nz+e1e79u5LClgjaKGixyDU+MCTHzKd
Q4WZRWn8Exvp3uS2cM1buWI9Zi7G5g/MvD0gD9ZF70+Y/NyQfM7vbeZxZKHQH1Oc
Fv7tNRg+LH1NWQxCmkj/1mBjedNd0hG1yu2LoljswBMFu20P22F9+M68+K6aS7vg
M/tnaywxBYpQDzzDpQd+0L4s60w6bdw+EHwL02P+mz1OO7/kyZHGOvWA20rYooHg
5413qJvAjyWxY1ccafyaHi0fQyzm8SKVGqqhM6vbRv8RKy44WV9Bz9UkqFGL0X63
3B2p07llZL6cYgWLMGpq9xF99SwiFJ5UK8WVsmaScrQOOa8SRg/DJikGv22rmwX1
DpO0cmGwpFb+iIcLCX+YuAyYMaGuR4nTqZP892R0MCkUhaGy1pMZY9kgQx2DowSB
ix3G9Ynix+ZBLg9k8wiTM+0uYALTVIWCGYW9bG18YPpTSRk4sbwtL/PwmbkHCMFA
di/wGHxJxKAYBcxE7swPbvBR5q9HySwaISOACYUAJA58S6knH9zrxhjFqNteOPPg
bf17znqdncKNhD3mmiHF+xpDqa5a+NKeHlsL4yUFaUHd8YargRUp2AES7gc5yKal
BTEuJJBygD6awGMxgAXwxo6mSNr+Ef3TveuJ04tgLIGNawVcXTuxg5hQxNuJpyhn
Jv3xxLgv22iQj0vjjvIEcrjnCKKwIN9jUKLaE5hB2LICjbfGlTCh0q/UUF2sKnTq
70zhOn3n3lHFDgR3aGFtTtxsHikwJUvF5IWJr7FtGCcdUuFqV+WQLLgkUoIboHXv
Gc45oNbrVNjlrs0ew/BL2DbqZrp3RTLsqaCIXeO/0zzuqTrukqClTXilrNPAcezb
ep7l1ttUQEK5Juj70hxwfFZVU6Z9fI8EzI/ayi9DbQ2DUcTepcg7FhvsjuIbl4b9
Sso0RmZDYemE+FL3AMaY3L+RAHRbtd0sXvgzVxlninOGvXoD7eiRJhNQTj8x2R9p
7ZC2XJiHFQ5q/AAWClSQzNN/psxbFKfqlJkZahduLnfggeYWty2FRA2+kie98ouf
2YaS5KOmVcvhFkl8bbxqUes50sAbLPBjgrUCK7Db74gQfp6UNw4Ebs+7UJAYLdnf
tuFIS+KE60r3yHctOxb1nGIv3JGzy3dYn7Jv0dPjJTVhdl06F5CACV3KiKqamoY3
LdT5wSXLvqwDXEWb6P2RpYv6qslf0o3lYd+Al6pf4+koGDN8gnI5JscDIh+JzdkO
OfylXV+wzOLC8MVpOdNhlDhh5qE/Vq6Nz+iuUxBbxHDK5EHDMeMBxT3mYP3nM38m
EfFBIGMRXf47BC97FtbMc4ngy02QG8OUrMFkOqtG4nVoBnvtk6GrN8Mmw0eooZvW
tXf3/a5ytqHFg2e7Obr8uWu93kCUwsivrZ+XLIETM6QBg0C7mUgN9140JMOgoWuO
d9za0TGAsOnvDvlh6AxvwrZmfuMfE332z7i43YK0dXO6VP92Y0ZKWqGTHIU5VylF
/jjrd3s5W9o50uArNIy9qYtkx+YYGmDZjX2QMaAi4yv+3JAec9vvak52ln/zOhvl
+fhguw6atoZtukNaJa2Bw/GGwhVVwyLVQb0Fx68a/pfLMBiBUPF8dBAEacNJAm/3
UBODBr3uhNBxPUQatM0Z+tNljLDmT0288KUiSBvZLBGK86fx3gCyO38UbmwNviPg
O5Q1FTOQTV8kj2cy7UqtMN2gwfuW7ZyCGtY1bpKdcWt18qlTLPnR/YVi7crCIuy4
OWWszuKfdFvihVb94WyRT8B/Na+p0EPWhVmcgR/P/dvtELADoTOwXftlosVcRTh6
a/nMJdTYkE4NPgb/K5AzzoSSWi78g6D23BI9lsTRBQSaHB6D8umygU7GQiZoYJEH
5yEVwXWEnAgMStuoG+WVB/w2v/pxSsGLCe9AqPTxXvu6u3g4wQURqo37mDkmcPea
E4YwaU4OyE5A1pgN9nGLouo6jYC74QrEgx7GIHAsjgbe1qV6yShP/E6MpyrLOTvs
Xr7oRZQOocyxbaASXTbSISoG+9iXazmmzaBvrNVtJIhKz5unYjDc81ta4qNGUOqJ
ATK6T1/XCYCerk7cqKstWpwEFml4DbwQCKwjJfQOymV/E+f9OLBYRp2EgyVVf2QW
/lYtiZq0XmeOEYK8OYj/FYaGPITfGi26L0TWl52ckMb0vqTK2GAbdtIHWPkczDpj
4lyABuPXNeErDsjzLifcCLDnqoFZHT7yBu+1yeOG9cLWbuWdUBtmCB77xqwQxVoq
EqNzRlLzECFLP2zFQRfP8xxliD3Tyg7HSgIMInx7fSQ1kHP9jxTFUX/BA08/+KIl
ob9OExuZPJEdQntDLTZFK1c+8UwjAXnGilWj87qEPMP/051TpGjdgSBAx3ctGaIB
oHLoIEKb3pwS+oRhCy/+qpO8XTl0adLM9FZRg39/Ul8WsHwO2WriMzTVK2f06FY0
Ql7AqWnaSmTfD/rIEbv3ToYDK7QnotrTNpv9Qkmp+/dtqWXBxzBsL+P4yYl22jQQ
lIY0PkW178PPZjWz5y1qKmP/6bACF+Ez6DQAprxVklW3NIZU8hyrLA3RgkNkgk7h
XCHa6WKv/TzSgl0Lu3CEkcTw+6XXZB8CspKG2cJoIklX9XG6A3BJfa+82Rx66wIv
VQX9lejMdEzMCK31dcxDUp6rI5KWzbyrafb4gRYna0szHNe1K5jPa+BxeJ8KK3B3
qAQjh74PxzT2pW4YH9NOZXNmcmJyCLydB618WYk8rdYEJoLdIir2+ZqIrDA8fIx1
UUnwYF91uXW3OeNIYHJDDctoxTClf/z6b0d1qYV7OGDXdrh7BqNB6XLpHYFVzw9K
Q7NqP2qL+R/M67tzrEvQzTxsWgklRmxgjFm0+THr+5lXaUIl4Wn7R2UxH41H23so
q6q2BkZO1qmX5m7OXXtRsiIiagdRbK0ubhi6hN9HrkxNy14xH+5W9F5n3sFuYGMk
g9xDHUdjV3WxVj/dRZ9XPENyfCTQ426xKvFFCK+wzOSjweovfbOTh9tqjR64R5jZ
OsyrGHwa6W/mMLMRS7AWqV1ABFQabuYyejxLrohgGqxJ3RZs64nMICQt7+Esath5
vQMhaXIVQIcE77u+2MiNuiIAy4OL92+9QyWZfM67SXa0wkLSlTd4sU3pMyzHVUKn
F3+CsbR4qGy0V423l2TT34BHZRib1kXqUs76nF60rpKaYRb6C4Cfs5JFrJ0ot7Ed
Yw8KEf6P+sCWYWBugDn+nu0H7f1pMU0UmsagZ30uAh8WejtgBsqnXIndo676i978
HKjITsEXqN5W0WpljBRsUHduP1XoXoszHQt6PWfGesI9mau1qZ+9BS7CvbheeU4o
NEHaVbvGW7cIR1qA5LjTwTiiigfGMA+glLwzPlqg7v/1yb3uPxHCgsSXwZ2LqxcP
gBPVOy1KvCGQ55eM+fbSLHC6tg8opx8Jj0k7A6Ef0aULpAta+E/pfIq/bpklNpHi
azddNuoKemUdsM7NiTnRU9Ith6nkQK8iGOqlvc6f7DLWJ5ldJWzdIF7HuHtCpqw2
zCayhohzKJyGJSTWaauqVjhXE7QbXCPY9lmtSsx6GcinRhYpEaXVwGStYHVLo00J
j0hXWWWrf+wR7SSGujZ3boasJLvYNt7xW2ufpw/hK9U2LpudSdIEa+J5tZ0J8hMV
W2bTe9BATUdV4xX1SyQrHb9Z/krr2YampMFXjcbjYHStEWlNRW74kL5ELKNGo/Ve
J9/Uz2Fo4QkKfSNiGI/XTECzYLxsPcGObILMAdjafGlR64Q/lMkChHFbjSAZRoYk
U/D3RvtQOzP/knQw/WkQ6cWttI4PMN33IMnF8iB/H//iMkaHoAR8mkBvjmAswujG
Zco3DI24+ZbAvmJJRWBS7zjX+rVk2zD9x+C1Krgv2D8NwiI5QxAzj+ROJz886mOe
T0gIuVjnvK5cRZEQmc89iRA+QOEVTobW5WBjWelUqobOeJA5m3UUnYpcHYgdVrdx
ocPVP1LGJdr2NI+EZQqhSxjec1QLmyGDD30/0IbMGAtG9Fbg+OmQI2AUlojFn+lE
TSNRD+no+G+FLl+NDC7kc+g9wlgeo60CAgLBhGSVtN9fRgexFJrb9x6kdnbKNN0y
GLi3V5Ilx/z19sTxzDCRB1uWhr2VxGfZY3rEAlo4mhA+sTZlglnGsHRI3rdSQrrv
He3TJneA2krUFY5Rd4/00FN48/rf3zB1Zvkh76tAOlP/bui9rvbJpF6MncCds3rf
Ysai5aHBAa9vD+oZDrbX5X4sNLZjIZI+LzAiVqrk/x3eZLpQ5+TFDcn7dCnt9hbW
TOINetMEyCV+QgIvdSToaxu3M5RumJLwldbUyJIro5awomQUHKCrv9TmNhnyioc0
LRFnSCOOPj4B13eQEBKc7AP3yx9X4M2fM5pvMzWafT1XEBqRMD6ue2OOdo+pQzoy
TABd9ghXuwyi10Ut5Y6UgnHHi+2GrOVpI7nxHJO8nr5L2GLn/huQKHDRkHefc8Jy
rxGz0ookldq0myRUlwKzOMFSktzcE2lDKwF1z+AUV6H2qNhzAAjaf4bl/MnVE2Xh
nWmG/0NNX0IWvTJgZ8lwQ2qdGUyxhi8CloIUMLbhsKdT6br0VhlpYi3OVZpdt3iW
THrg6zEnSkPbaPHIKxomVPRxwZ/c+aEs9uirExGwu8AMdeiRlACEtk40i0r1ZbBy
zLv7TZRp7WFpeL3/Zo/EzQ+Hu78KXfgzw20x5M/IljzL6ROQd/PCIapxZMi6Sjd2
FKlWfnhULcKqwfarYGd6Sz7V3KWOB+xXrug/HdJAJCDep4BHzQ6tj3Mqh15liyO1
UqHV+tdLgd/ld45OY7JUHrYzjfjLqpwRFmI5/kGDhNgPjI/UekPdsWHz0rY6EXrz
YEAxkrhuL8kth5FlhpEMaxQdQI26yPJs6dLfAA5o8E54hONckAgTMZTH9uBhqzqV
/WEBkmLaglJgS+7KGpoC5Sf3JL96s5iNEM+AagktdmtRfoFZ0fgOyIwSal44FGMY
TlHbRTkjozExMesgeDua6BLS/Ic9WW2frourMimbq/ojqzcVZIFOFyAjlM1U5diV
3pHlkAsdQjgIjt/2VKJHXpPMl0nC9o6SCn1TTcbs+QmU918+VbiWBxpJyG07YZ9W
FtFHOi8qsc6RjxhE0N/nvzYQ2QRaLm4HUQVH6WO/lcUapZTQ9WYOz/T48JeueW8y
QXfaMaI8/AwJ4oTH7UnVL7DNoWky+B02xlT9rMe62vZrlcJ6hntFyfkSdiUDhImT
DJppVGKqBNvH2d/Cy14Hbk4JZERVPPh5+IkysI5AcdisLuTnNaov0QaqmjQ2TOGg
SJ47Ibf90w5/2hfBH9dGjROKHa6NUCVZqykGH8fjltbDFqbzvbHz4riudBu0jxZE
EN9Tbv0vE67oLIpDhNM6h7y2ETBYwzVkQwjgKhTXPFjThtsJ81T8Bmn422VqOCvO
L76+8+9LIm283agQzbGbwRTWhrsO/I8ObyL88hWRv1g+q4ekbfJ+UPRKPd0a5UXF
2zpImNBtGoFkg1a7pzE+T+MG7fim79VKaBzMtt0VTXRK+lR36aLkQqeUa6r/GV9K
bhjuVw6253hSO/lSJ8BMHM1lkUClSGb/poEnt8QkkZ6534XS0O+ThY35jy0gYCo9
p9pVpA7VCn2smq/GTYHANKtSvxMCpJirNe3RCXFN1/yarEcdUlcdBWUKqaZembHW
k+NtsRffkaF6e354byWjboqJSpJhjN00N3X+CDeGGNU0vfevnqIcCMRLi6TSbmD5
Ufq0zgUUTXz6m7Vqln6kdMPp/D0+JdiHQMhJaqj87zhIAM8WPKR+zDkXGY1vqSZp
JeVsVnuyjx8BUR7hh6VRn0iJhzIUfTS3rVa8cMizgbELZYuYWqQCAWL+YmfcsM4C
xtiRoNi6pOGzen8F6gIk3i/8ktfh3FBEO1o48ujOCuOHHpPlZro42BBD+RUVQzgT
eqQpHlr+1ezGQznCYPpznMV9fB8bX0wN2Khkd/2iT1n0PKg2t11WZcjj4ikZnqNd
MPS2eCN9XV9+BUBqXu/g+DfimlUVZpbOWnG8mBbmLz0xfs+imQYGr4Y2W7b1uZYe
RA2zxsq0Urg2uZUkjUjED3oEMrzmGHgJBIvgZTlCpLECXVgPUkRMEgaI/VOwIr1n
hVAjMxCWo1EIxXfFuKSRu9ualZpXad0SVGqHI7K56/dtRjRsuvQypqxyLiFnZx07
mh+TtMuL+mU/tIAItWqudlJG6m7XGYEohwZKVLez3hs16cdzXtB1Lql83C8oyTJp
Kl2sf4lrF74s/3eZzLoom9dLj1xUDcfRQEj9gOpKlamr4//nKVpyEZEcXEBCMwo8
RMZPwz2ZXBE+AYI+SirNlUzC3cRCvA/hkxhBU8HpC38FEzfvRCIyjjMV3uOJdgbI
fEAAZlbCSjgGYdCacp370DKJ/Q7bcaBulcX9ooNkV1Gohl7Xrp1SeC29O3Ui8w8/
Tr0HxQ36iiDKfcCArOtFh/7iY1aNcczcVOGA3b87NmSCcUAJcaga7q8bUUY15xn4
goEFNyVAFO5WYHrGWeWnbZ8KFxePKjfXyfyi7YQ6v2qPck2sBzcc8LftpTubAtCD
NUsq/pUX3kv9W9cEiPKrx4Huh/3rw1iwu02y/ZOM5h3kiWMI9evdEy47TGPp8t5q
1XcINcQnxKvmLiAVGmC2wKMYN6OJrdeXnO5lfjv69pCg9gogSQRzGc8Yw/VTgFEN
xDT/3kvrefFt5b5NMOFlsYUwghDw7eoxNbu4qtKQSNYB1hOepnWhHZYxNcHBY376
FHWoqW8SYKtLS6Rp1YGBwWj29Ny8cGeuecHaclXWUfrRCrI1vRB4LCt/FdcznwSE
8VQDQkMiv+2mLQlNVV9rGIPGtoIKQLN18tFzCKT4kGzi6tMx1411En5d4j/OH0nF
8fyEq6Y1jvWIsliXJZKuJgNSLjuLmGtH79kTLyZv6l5KknfEAMHbUje5u5A3/B0/
84exYB0kxeZ9FBG+8Jj38UJVJWLsaN4IBEj0Bjs9oBFcsswg+IVdQQWf3OHNxKl7
LgCCcluLv7Nef47Mhhlbx2L48DGMdodrvjqByS/4uDCguMR9pSINCRef1nS4bUuD
2Ynws5bagEgLsCpRZZdyo5TmHguoFZcse0OVyJJMI8vLj7qrQd86y9liiXrk7/m9
zpyanU5QsRx7icQVPxPuWIlV3IlKhDtymrfvWacfzloTWZ+CvPdcIG/YtP8WpPlZ
SMy79m87zGBRG75bk+6UZkUgZ/i4KypZeEfc9bn89pUyT9jBPnt7tHcVZENhl69/
1KJnn07hTneK/ior38ZrD7o+SFBpTt00/kgQvrKVQ+ayR2Wr4+yGeAaxm65P99fP
I5QP0jYlojD14Pytovuc2kQeU40Al6aWrFu2o6GnpT8MnMMB+8PqDWYfc/wlauMv
4aVf8umvmofX3jbks8Pm5TBjpTbY/SQAAtgB9tyN8y5e/MKRBma5qH2TVrBWeSbR
3CjYoUvm6LR2jg+gS6B61n2OFf4itrksMhOzer3sV0evpuxojBIbbb4U+xH42sN8
wFxz391BS0YAt/SuHt32mC6caFDbGI0ydi88rWcoJR4aNJejpaktMjUarG/wrWvq
St/wNu8VS7rIWDl4m8FSdTvtrsysIvl+0FV4Azo8jst7pQrTxQQQMMtfvwr2pyc5
a22M+3WzgOAe3z+mNfhRm2yv3ZFSs0aNNXIdLb6Kgq/nAAAIuQ+vRmuHatQghgrO
qrfh28NMSy2soOeHCnxRAKySGYdxWhymt+XoiC752KKKG80Ok3LSNnXg4fYNw92c
ObpLQCEoG2VT1hoZnodu5E2xXfRewtvF6/ZHvztmg2CrISUpw0NcfPoRjih/tM6n
qbhd+3ByxWmp3aiHI3FyVqTAD/FZfyyb5Z0MhonCuKLRLCfc6n2T6syL2L9C3Md0
SCklaafjhF70fg6LLw7n8Cj/HgcSxYC+bpmpiT+pEClbPkqzYtP20r9uiH4fIyrW
qYzj0rgeEMj0duRklCuNK+JWvW90cWYM3YnIWNEGZadOEXmIk9QhSmEDWlWe/Rdd
1I0TvakmpptQr3aNlKGlYjxl26FTKpB/eHhaGrJvnmLfKvnzFcfGKvbjalsLRdY2
RhFxzrGnmez5GGwOejyzTqGjCal9YV22l637+RDVSYX0YVq77wXkb6Qtb6IBnNq1
uK/24C+kYQirLfIBL6YOwBLQaS2+XnQdYR575PWImnOQlQV0xEBG8yhU5AMi7F0J
YNudhAnMBDWXubEYKSgggHi+Hzg+vJsdhAdyqJeyPLlrAOl5td37v/YwLjoPYk/P
AQ9/rMhz3y4VD/jjvaYV+bzswHpR+PR1h1hOjSv27q8KzgOG8I5n/W1ewtFXKebn
8+/CNAdLwO45JtGhO1iobR8LliyrWeVA5/uGU+Od8sUupnKSw2hBwRnb2T+ykoUT
RUhchNpzfUegBL0UED60lfP6a3qZI2+ckbYraO/KCRIfeS34oIWAYI+jw30DJB0q
+xKEk4dNDXf7IPfQPfFrjPOvxEiII7Z7BQab4LrUhwgbPOpwHNvMmKBr16EkkPyA
+sNR/adC/+wEsA6xla65IomMqUNM+edP2eOIh9i1tVFf0pmC13866ba51Jy7eRFr
AJ+UBRwGUosJhr7LEXsL+6iDblaSJPbycE3ZbH8uIxUlWd6dOReoA9+xG1s5g/aN
oBFF7OiOu7WwBkMEC2Fz/tS/vmQmiZwmsRIB95QH15gq8BXGzDvrpfG7fj+9n7AL
rwwwdvjymSI5BtP47exAboRm6cunn7Ecwb4UdpkEkKOe9N7CqjtuHd6nIZGtmoeW
55RN+Bit5jvcs3vKSDNEJyC1pNh6UtpYWqFgY8qw7UrhfRb/25mMQCYHEq7t/U2F
7KMPiMt+NgCw2eE6s5gGnr88Xom2L6iTuTv952L8XOmM4/yAgqRjw41wW3cdXcgj
o2/lwNdplooBNLVBjj91zbGs2L2brZ2AKhvUQbVvleyPbsuA/i0/mKWeawbSt/3w
KFrORynpCRZAXlU7ayP5yPdxTKq953NieXoXGvDyPGUf2LqRtH5reTzZpw2tbeam
S5CNnv6Sd2+l2zCT1+/Yjg1aQcWNoGOXJqTYb/bE9trcSleN7yl+tKpN/ELr01dU
tRaCBZE+qDMfS7GqnCQuzSqejiO4rtHnOUAOOA4HyyWHPATOSJA3CEZwaXwKhkFj
q5cONF5sqFk8WulJlbFzi1pnZyS9gsUFVKna1JKOO8sGo7Z/39+lsz3OSr6QQAwn
1AS3w6EY/A/bojrNPVhpk0K5a/Pp/jSm3ACtQXy2P1Dfqk996SSr3IuHFynM36Sf
t+KDHyOroDOoBRNlItNfv49AVX7m4/Q3A/3JvA6XxSVtqE0uS4RnoUCj0XWiCgHe
+LYluCFgxx9Z4Qq1AF7yfuz9IT2f4wWJjYFtTCCeAS0qhk8RUh6yhwrLVLZakUrQ
7dDiZ6nG40JhlMomp0jGLDJ/MDqejeqMfRn+cf3ZtUoWOs0WesPXSnjYb3wy0ron
kRSmP0Mq6Po1bnFs+kda5EKinoLjyg7vyG7bcphw673AxdWfPpk/s/aDToWWtEQZ
hJfwkYxzb5WUYub+2xbzzVjhtF3w/VokppDB4MLGe2lkjZQz8KMI+Nuyp/ojeytI
2VfB2ZVB5kh8B2zPD+Jz8PF6oVgQm0zYs4asMiHmq+1IbuSslOBL36Jx73TSW9Vy
W98c7aW29xseatIat6egtya6yIX1tJg6g08+RC1AyUqNYsVZw3tLIHM4bYulfzY7
+QWgZZh87aJgxIuZ/5fpEFvihi2rV2gyOU/UtASy4C5eDSnyXD8FRPOMiefvvhCh
Q9Fb+dlGC30+jrbGksRemjBY+oGEDtM+RgpFJRTCdtW5JIKViRELKay03LByxV5G
XJu7z8hDhAaZsi6WquQMP60C9FXQII9a0UqvpHBaNGF7VjWBNu/ff9T+h+z76BzA
xeEF4B8VkvXsbzKInfUEIVYAf6fARBDjQRMRbDRtCXENt5k87qcQtsjKCVAi8XpH
0n84D359HseOTMjfBsuVO4fCsl6Zm4LuzwT8U7l5TS4OljgY0OuyHm3pLiA3ce3X
gNIj7uZVqodJjWADaVbGx97y+Bgxu0vfVAp8k2Yq4onohGjNwP9LZU9ph7n8Ykfn
NlAonkBQQ289S+GOYYnmtB+qDzvkzBnQxm1YovfEnMz5behALEyIfIVO+p0zxg1v
wsD7j/aCGUCwuSLN8xj92DlDerUTMRCnxu6Hvz2F0OPkPVZBOk5sjBcBUloTTrKW
9Ys0lFUxEqXKhjeeRPjBLW5vUqsX50Y2eejwF0t7BSLl6KKx+Q47i7z4LX/HI3WT
Tr83YZgognjeIuWYYsOIIfBG/vZYz1/iy6C7FMjKKGdRhiYqBIuyoD7Cf8GBFgEd
QG5Xf5kfuwNJHwNtu/Eg4tXKcMVue6JIdoNoHLD/616NzJMrv5b4jWfF4XvtEdpe
81tg35Q0F37gpbHNbi5LlEVIpnOv7QHMG7FFMFxrtSU13ny1BWeLXyHCJEpHbyvU
SbqBp6FRIStc0MZZfHqNMAoJ6jKbnGnvetgNVQWIDnpmyIsIcs9y3jOTd5YIwaJK
gZC+bWu6mRkGIWensd58dFds1pAesv1aIIaEqELkDov1OylgKVfF/Iu9lh/YX4pz
L0e3URKeZyv4V2Lk4/oiFC46H6ectoBtiXFcSZi//LHfHOUfCzc+SYFE4wXmHzHA
GUEgoUvC6JlyYrBHvOMKLwie3mh5+0BrfTLxgqxqc779DFBlw/OUhY9bT5hD1mVY
mV2/CQgZgCokACGv08Aqd1TMtddGnfYspfNMFY4cFmkrf4OnGJh4ay0b3/CjIlhW
9E4Ev0uwN30ffgo6Ttln/AjPNCSMjzAtGO6F4HRKkQ9lXyGjAHhhIYui8UUY279Y
Cq0cZdA9N2FgRtyhJhHkHq3t1p9THQ5H5AmqZog9XLxAY/vhaHIVFdI+GaCV7ZGI
ugQE6dqnqb4rKJp0OBeXv29225tyvVZJkK1eewmFNl5VMlEtFfXsgYKaQBO8jFOF
+zqZVTXHV+rXKdxfEtcC0tMjlG2+ge/8ApIVcM/vlPH8tFvE+VFz2eRBhZXGXNdD
F30BvDa2zAfNA0Gpyh3uSQh9XQBs/JSI21kGDdzO3SFysHwN7TgHMqfi7qi5+DfH
UagRPhjClD+ROzsaoI2Oj9n2bpwVirrZ91hc68DvtHOvj5wyQT+WtggczQR4WqVw
ajetrm2Cd32/9/Uokd/+LCRRg0B9ckmIjOip1A7esFU4AxJaxmei9cboVw7jnw+Z
3oAAtprCSOE72Ov9R8DeCLLpsmhIAp+5UxKZkHYxYHoKU7BUBRtEU5KmryxWt4ps
LXoRke6li9pO6QTuxdrV0zMJ9eei3XypJiSc2/yWnGIB2RC3MPM3zKLEA7AdxcMD
DiGmQPd0plxzGlmXvSdw0CZmBvP/Ne4boBhSTlDAwwTkOKJpbGJiwjiAB0wFk02G
q3YIr6DG5/3Oyqq74R/fgbB7wFVXlg+vMO/Oe9mpCpYso+4hyRhBi3SQAExjRjJK
IKjTBsbLtserkWtn50PmZpyfi97iUdGWBK+yQBeCwv0VKwg44drjsrJiUHa0AYkG
XEGmgUDzpvUgSGHCYS2K0XGkb2kLOM5atDnb1dulPZnn8nxyazL0j+5y4VYSmTxF
q/sUqXZjDf6OPDkTFlAAXoHUCATaDBVQB7DNOh9yOOlMBSRBRaIkCtFbd744XN7l
RvcQDZIdslwm3aefL914UN9k11wfw6FdEt8aF1Ue8NG/edIu5uKgM8fi9LtAGoOg
kH0UVPsDyg6dhbLpvQlG1DjyLSU3z64PfzByHpz6IWFiMNx/7VrU+X/SoNbRVL65
8O5XrGO2xyPfSR1gZ3nyghkSDwAD3nimhPxgEiaU8VvH8Qd1AYAS0Du82Ipl+ZU7
Jram/tK7SGtFljF7Gl55/XOK1o5mqskKjX7MmcpTAk9Xv4FRMIsBi4E3afo2Zq2Z
xF+VNe9+I/pr3bIgbWlh4iLgXsWWPuu0CgIZ7rX58ORf3q+IbnQ+yTgEWDFY3IYV
5Qs9ITHtOKnm2Mp1U2m62zrZXzmvTLKnLA+AXxykBIDSj1/GDA3tBTwLJE9UEAyF
2XOJ4XLUXpQO77sqgV7cC/X5kpZ4mILm+VBmZRNOme9aB2pSfrKlYMWkWna64D4F
q1bFk+NbEgJLqkBOfIJEs/An9ogbaFAa7VoW9Sr3leIlJFPEAX+o4p3E0aTv5oj5
f1o9GF06BS4DRoIAFI/JlUbYCAzxCXuzLCxrepgsfUREXrL19Vy4G0s4D2C92JwQ
xvcaR+d90SLgRPbKSXL8sq27pOJbdYVR4MMGj8bJF6Z9S/F4yv6oKNZi2BvCmE4K
vKcv/0v5c0FhJhOfUhQmSW/lTR/QhkgA9XIAM4lu9XV4EWNkGxwdvg6zCXYteu0F
lKBcokGeY/ErYedIcB/t+/2N436TYJdo8jV+JnMTPpEq0vUlEAfDshkEh64w47dH
dlHKiccTx5nkIeF0osNVUAjk/rVYzg2z1IbDPxI6n6PdFZdMvp9k+Wu5XuZTQ/To
DS/Bmz3iyMFOIiw0Bu8GNgYA98OOw8pBs2bzRmRv10gCLkPkN2t7GIdNGOQwZRan
JfhsfW7sV+GiSO6KDUZGNFAdN0XQtUmlucAgg5Gh9McuCclW6qgncdjNyWDtO6i7
vetdnHctqyHJ0T0j3MHeElkJ9RmbGn6PeTEkZhyQA2nqiZIgexx+QJqtxWtdc4mQ
7S6T4EYwSGT4pAC9wN5YC/f0ao0wbaGRmMVd5hZQUkn46FETJWLecbeWeHMkRVDT
rRavH8FEK7/bA4CctntGQXgI+sPkvbgRatYgvauX9Rp+Kr2WGtLpHbjUlYoR/AbK
8hzkfMJkJaX+pDrML9mK7ZAdgAQ5VUXoiJlc40md6YVerzD00RFW9tJCTLogU2LO
vas/gwxtceeTXajsvY9oktrkjDGEBJ+bY/VSwvzcydyRgoSYZLehmbf4NQ1eu6zv
Y2sT2Dh0skscQBiOczLC5pdbQXCitwKVhjGXIbJTH4je0IEUdfslb+HdIORoWv0V
VAaKFJyZUFI4TVcZX5aIQu2plLzHTjglUA30V5aLtoubwX98f3hYz5an/zI9EnZZ
pBZ+whs5DYnhiVqEQcaVyOWJRXwfOedEKX+UlXXG+Xg9cR8q5zT2YVv7FcxolKac
LEvaMHk/C7GGdPl/vX1YZteuzeBlaWpUg5xAx+CbymIz9KZLkmT6EoyzbOAL6EJo
jXhbt2M0zxZzGNom8hPK19s7Mfr/hETILtXsdWBkQcVeXVIIf1CWI8FTRJbkPDPs
cyJEhsYfErHFJsaHf1CWkIGMYGcbQBcPKq+uDLFKW/pQr0P8KZSPSDg6GtDOfiar
8bvXOjl9uzo78Ex2L/voF4oRM+rSlxjkxuYv1QO0GPWtRMUEz/271XmT8Hpxj109
LhcHUbUCxguKq6afdObDaIVwp8s288ktzdcyKdLzMF8HTr7o29chlh4FyGGuGNks
3CslzVV0353JisJxHCZ847ZpGrxG/NKdA0bgRZX5WEeR07ns8vSda7Sim8W8MDVa
nEWvCW+h7g3j2fFuCHkwyQAljwDKO/KYTl2Kw5g91cIqwwz9AUQAkAID48ftFT5E
OL4geoCXNhaVd7zfZXWGffqkLd9fD+P4yLYcM4P/RO9v2Wi1AqxWaZRtx3mK/0nW
akM/ZTieKegY1ljpQs9XTxK6kIpfxnddWSojmkGMsth7BJzIqlBYVTpqDOxCc4wO
LRUsntyEe0wKaCHpctQca+FERBJqj7KtcEGxVWE38snZx/JmF25hw/uBBKm+OyR/
W6ZC4X+KzGLX7j/4tj7w7lLO+IMdyHiGoKCl8eMiUw0X5+qycE/pbasaYSnbedEV
NIEistau/hhLwpJPIs9pnsq38Wn6ee/B6z9gd9HX8SEQ28K4dojeY+Aujp3gAv3X
ptdBmBUjbujz8gbqbuD8Z8a8nv+nrtTXVD70cezQJWtrS8i7v04wui23pnjvDJpg
KW4GR52yL/EACszxMZ2oBh8mvcaqbc8GwzdfDX8B2hxikfByVOqUz3qv2IOYYYSM
gfNeS0c6nKdtBcmwYl1wiFhTfKysMgYsfXvX1GdOfYNZLJ9qiQCE45BwYubrFo9Z
Y30P0RjiCYJr8CphJIKKPyWm+KnhGY1TI1/L1lAxhQrs8bsmLeWWkUfeTg0ygx5e
fn8tMI99rt4HTqVE6L6Uwjl5Q1T1HXIrCVTHrvHBIg+qKlxE59rnbQBGNRIRhU1y
S2FaIm8EkmkPPq08NdGKsWAIivcUMvaV4DNdGJT49RoWfqcym+YPEdz2Ob7NKuOP
Zbjc8+QUI+pmE5AWYYXNb0vIKlQwi5sTYn5EuprD32dSGjyWnfv9f7paobJgPJQx
oOoHCJm3vaZt1RMTrLBTbe9/9M4daxMmMPM9+aWnkxmGmtBNlQUZ8cLMtahww2A7
hGl+jFhhL2l//spl6gWWuxXiTOvuHf+B9KJybvUZIfIvIzufNY77kNrbFZthL+GH
9/NOFayHGEaqhCJgX9zzCjdHEzsuI3GRW97S8t2lPjWrvwuNk2rJi2yjUEfZKNFT
fSOYV5Y+kk5/HjhircjB72mB7Dwf2znDnHRL4NpIPVn7hFy/Fc5nc2NhvJhhXyCz
0uqecHEUeX2nmV0dyEgriF4oJaPAn1R8n7mgOmen9+D5ErO5jsShSyulShbQpmxD
+/cBneKj6LNlcU49EeS9h+H4ipvAGacb1BsFg+Yt6/2SmTK7Lgae9CsHdabrDtGe
gBBurSjiuHxUhqUEaMvWzO1rjEf1XsrMYQATNtuSV7G44/oDgET7FcwDtYrpN0RN
4qrorqCt0tl1lVkwCQKnT+BquCCR2IhccdgqRTV8p6o+9qyLcQRV3AI0YLEsNqMF
jOWF8S/5W5vaS1NOC9yFi5w7Y4kdI2Sx+YkiNEkv08H8vzHrOqpV4G57iLPrChen
6zYXHdViNAMNITCjJfA1TKTCte9BU+PfDiJtrhZe1lrDq7furI500Wv7+kvwxQne
RhB7iUaAlb30xItvMVOSf5M5IybCgtaPTOTfY0ec9T4dTfIl64rD0WHbNf0//AG8
1x3eL23vLuWPvIWQqY945PP9SMRy8yU3FX20/yNTNqNlA+sirlogaP+Kzt/Z8c+i
w0mEmqRTPXuSMTEKcvOnxun5UlOkBBmqv+t1ARF9/uTVJzmNkh7zGhQ+TLELDGIE
hPf6TOHmGM+mjS4qRyutz1OKKa83C/lC/vaHfsXFSA29MUBX3q2/7Qs90cZrAzlR
nGe912FPdKQX5+xswAnTFEpr831vL1IzcX1eSiHyhSIb6y9zGBC6oCOYKoXiYo6d
xSJShJjcCGukUb2QAdf+NkjBx5yYsAgZrYPEqmNlCqlyHdKUMxjeZSgXd9954oZj
fGhVRNmOWJv6Lqvgnl43HYsMEyTDYGx0lLUDEklKE98v0D7F0d3JEiO4I1Dj6OXP
rb3IgK5RHpRNp2ABg8eJdwgnFpEAgOR69J2d3F5oER2cfrmPT7ahKLAOmqwEx7E6
Lsx56e0v0/c1RZiOeOLFnY9eRTR2+KRg9pJO66qayadpZDePInnqm0w48FI8BeCu
5Qik9WYOmvJ4c74aMdX9/pLze0vaeNnid9ydhRojqzsRuJwX4Hei3j4dMfqJlSDu
2Dp2lZsHP0eFGfZqAzN/raBiew1Yxc8FPHo+kVa5woY2TJyCgubvdJTtKLo9sCUZ
mgkKkpx7HSDDU+KUrKmWaiyJL2CHiBUupLqArEYX0W79uWeEIARxhQOX36+VE+uI
dTZaBWSNAjbhpW6UvxiHnWyUG4p3DHxnkyrK8ZPTDmPbjHeoYzKt9xxqBOzf2Lhf
RvUtaTU3gPsW0VFl3r7l/szqtGeMLMYD76J331/DTE0UHC/oIYWHHltV1EMALgKN
lvYym31gZr25715eu8MekFT3j961xzEfNJSaNoFqywq1SELOMXiXcOGXWfiMMvve
mB6rKO/9x1tObkJYxrHysVXSqFD3jdYz10PKa1ow11vHhvEIFKeATKn1S0EwFszh
4S7M86KwzU9qePV/jHgWiNzB82m6l3UphZS0t4YaCtKRYtD9hkQr2mB3g3Gk/40o
oJgZzNd7NChO0AHsI1ikjuGitKWsQhg2fF0tRNlq1dHyyX/quTUmTBTvv1eKX7ui
wVDcGz2Xp+ocm8kVRBqEGCqedk8GR/RAmfhE7ropBZYn/JnbnzA0XkkZlK8uXH1Q
y2ShUcC9+uaMo0h8QuZI3mHH1vHTC5X7F7T/5GWejDcKWtdXdFLySaQ/793/fupv
6EeMbbXBFpZT6J/2WcUmBCVbm7GzXlaGm1ZPK+9qchCa3rRGIr7jR/U4FVjDik6A
U/6n4toOqEo/N8J4r1teGTBQjmVYVM2jJyKb3zoX2A42bCa7SXE7hBDaOC7QElJK
F5o39a3k/gcC8WeQuie0icv+ledEym8dFmAlbQcAY5lVfmFYksx2o/HSkWXSPxHj
VXEWQ+h3uYFu0VUr2+W5x6kKvSyHMtC799+YmfWDoU4BOBGbWSbBBuRLtjUqeIJ/
JTPHro3dMlWbfKq+bCSuVe3jV9NugnpMX388eUNN4XJ/Ii34+mccJ1rTFUJ4PDst
igEYb5JLaqKNAjtHyuVOzfBADVK1sPwhcx34z12mPmifq2TSp5HHow95tZtcds7x
QNC1ifwsUGgW7LP3lEEUWx5XKtAUKBwiC2DcZvTVNgsptFiqlEQewiFL4Ca3npqD
tUzQ5FUXxS9MF8Ac69CX81dgE2tSQEI2neQgSmXYKpIxtNeEi6HoREX0a7B0ZmuY
mIlTME7ek8fbs4vU1KTyx7MOnUuC95f9Bv+tkkuNAi9q+pYY+7NoUmDgmp6KGuwv
wP3xzZxBqZNfxrASgx2JFgqN0IXph+EevBaO15oe/edDSre65OEw/xC7QPmthUWa
7JCt3LywLvt4T9Kujgo3ZhiUfJ+NL8lj0I7/myVP1aSfcM6sgnBviD2ISSqYsv26
qrQCv7qf5Kv3gtKbcHQirnHctn7Zk59elFSTrEimZb/5yY9EBHRzCxp0RO2dOnMk
Zvm4LiJCCuZ1Aad1tF+U291xBCxY5MgtzONWefu4FK6wqt1Dbngk5hrWSdl70fAN
YrsW7qD69QdKLhja2L4LddUHQPtFQiMFpA4VD8neQcnlNfEPEHdpiE4lJRsWeZtm
JGEZ7Y5I0C61xfiA726hVWgq6YI04CVctuqKMWBjL6fLzoyYDtwNiDLsT9NfwPoq
oYYSzuKZpPtZ5jm477eeuQedmBdg6Fk+tzIQrWM+WpTExqL/2xcoTNaHdZvk9B2A
ts65Lgqu01doKkEHVZqKTZCK+3VtslA+Phsq2cnSDauCY8dvOm3Tf8zCKboVi5F7
45rquHxqdCKNmJbM/Btqwtb/Hpcj2ku1n38WHI+RvjPsUk/ii2C7UdpyJQx5eWCd
L+i/GRhUksfGXaWyfEoTOX8yeWHR3vTaO/TDwg8oxGnEZtreTZieeea+hzwynCHm
BL8Jblt7WycXq/3VklG7gz+aS590nn7gGUlXWfbHfQMWYqusR2ebzlIdVxZmj31o
yRIuTPJAaBKmPx+eyQcjbsMBTlGWv41nEjQw0FV5EAphLBMAfl67LWdmokjESePb
MsKuxuAfg4UWy1LzePau0cDBWeUq7XcU6+VGHyzPrShFFSMA+njp8z77e8dCxmQO
KQvJBh2/jai6e4JvA42EEqEY3V7XPQMEW3tOQtpKyzuZhmq7+m6LWBybMbHPBN4R
wdgUIzskeJ/00dL1mLIk7f7KjXbc+On7v+HIZn/0yiowbl/gPNFc4zdQqVU/qZZ0
fLAZwHn9e7jiyJEZC2Q5PLUdUQm3IUlD2FzxiDgyvXBvI06uKFases7fHUwSUNMT
LSm5xtC5t7iX+GTU2jbzKXjNkWm+AU4OuwIEPYBi8upkBLdVHTifkYn3lD7Rapsq
Va8MLfPWJXfOesdhsAYj5C6UA8fuT/AYICX8GCsWY7tv42Fm7W483KwJeqNxXOz0
Wpiuse9hsLSOb7w0vItXwg+LtmKbPEnRUKCTM3ezLpEqjXfO7Wd7dk12ZvRKRTQR
0TG1L3lUr2D/I9kA44fYnKz0Rb9/gAnQrN3tp+teXPtR9rMw3DOILQp6xpP/Xak7
9akD+nD9hVIATArCpgzw1d2cIa0bbkR3U+1zdoZBr+ZfYoTzaitdmnjAhTQDOqMI
SV9TcYuMVfaNojG6wpp+rUcFohSL0zNVvcfKQ0UAgEHlkR7ZI+9yfBRq+CPsN89z
3tpegOcTa46RIjhMF9Xrw7f+NuJ4msAmAczO/KNReF4KGlcpP/jxFqDcdLAe1keK
qGd2I1Mzsk/IeMUSzpbGm5Y6j83LhOzqqvSF3OvZWfgUk9K7k7O6arWEmSnFYZNm
yFnr76weW7pJjspIySamR1hfuMXeWoA98bfdhLunOP9puq4C4f+OXDkB5bGsHViP
n/K9ug8CdTLc+k5CHEOT8BRMATFTJiRrO2tS85tQthN+KTvcYrui2gdb4vKnQyMR
W0IsQJKCb5SPSBNzod4SLkJo+dVw2RDuDiAvJUDiTRBzWS4pFYtNGFbBIcbsSeGs
uxzii+xmkQ+DAobwq8r1m7qpBZohmZ0huUh4RuiDswRSNjg+VjvnHZsUypgRVLKV
L0N5p927xnnX8lK9BHW+cIJHOSMZxmzl96VINYdgDUkXgVEGD2ExE8BYGJuzZq++
sxZoWQPObMUEnpmP1RNKeNVkRNZjIZeekygUpwAisR+iewkQSCo9WrbIoHS5Hwog
UyZnzJZvewheH1RMPzO/gD7bNrVwxnllW8NpHGnK9Qbi8k6KiFA1WzcVBNzlR0Fh
Dam26IUki/GvPZTAV0z19k8IDeEgP0SxWct+rzZrHH2GHERkvtu9dv76b6R0ylMX
LwM85pgE/z5SMJCGcQLKbMcKE0LJ9bRlpziuwvtsGem01bOk9Ps8jA4sq+68ahAH
DShfPgADE/II1jjGZLr5uRdQHK+TVJRrpiEsp1fg6r57FGSvECoyiglLOJc4mBs1
QPaHqLcWiv0biYqDNapiDJ7ZCzgrvds3E42wwdoZzsuUgYByGSJpbS2mq69/dAC7
L9sHLtE262v+BSiWGpM08YOjnYQ5NIxDXvZPwjJ/THeR8QPpptKZ+Z9V9m8ptK59
qh4X7SMfoNs0rgys0tbyDbH6nbSivNoS4vJrt2YO6NO+XgfHkZMrHqvlcA4RPfnr
9QNTEKkKvIyJ30nv4rnd3FfUhgi2+ul+YU13iPuvEXAvtOApWiZah7x0mosW01wC
xsctUX6UlwesVxxkTTspvXjhxJ/Bg3tx1k+1AIMzemwlnpL0Y4mtNoXpPTI01W0j
kPYrB2Kp6896Vtyf2y2dH1oUb9vExoffVK2MJD47+lAj8c0ceIs0axHj5faS67iD
NNQktfj3wYJWzZKrQaI4R5we58aPbrUkd7fQaJpBnvy8hFLf+Yg5TqZ3Pf0HSyIU
SxyyaaIirECOdiDIS6edG//8BMcacGw50H2dU8ZwgA+8MhYRoqnLxDE2EOtpr4zP
YL0is+PPnNAkytJX+376LkV3GotCOK8jk1G76lC4MFPdV2/j8kridDJv5qgmFUoK
tlPGi9Ubyzk9Q8kfjIgXTboYwtUvvQeKF9nIaGqYPSnkjBuIszJLG1vJRq9OcXCW
d7yyviG7zC2ORIBh84r8QHgIxtkt22hZZYHNW2MEpSQlmPxgQwVSXfNc3sv0En++
MjZr4U86sxgzatAOJ2oQqDivxmCTGyMFo6pdlUSrflU2J/hzFWz17oV7rBvm9kNh
4x/PNOWJdmDPwpySlAtCnrjZDbnpZgds6Amu6Omm6Q+w20o43MnZppPmuMaxatvu
eR2TmdtFcXIcwu2lR0F15dLDY0WX3f9W2EpZ9LL5KakXX2RZcrlUI9O2GasJ7iB+
YkxDIrGq1m1gispXpZ0kPscFTCDhUTdCOyrjkpzNsvhPOUF9cC8MiLHJt055NsA4
9bYLsS+ziyHKNGWKV3NCowiXNhKnwepco4Sk8EK9NZ7PemRi3WwXF8YwMGO6ynIP
5tH2kmJ8Rz02vdIf/uCf3WXNiYUxsRam2xAjOAK/rKVSwSwQNYxbtiOYTYRIWrP5
Mz0DTj6dTdRpUY61dKxynOxmXPiWizR1pZat1oMlhW0NnsS6Sldd75wxG2vTFL5y
XxVCf6/E0Y1th0R6OBNooCX14jGlat4JY7Sl67FvZhamO07xITDff0m7MFfdII3p
8F1xajPzw8q5eFwTULwVqEsxyuer6P5bZoRaVhKurXNY4Wb5fz7KVt0eWSr4wdwQ
mLWGgGmG/QRNupbQfe6yZr0jv1agpe2xO3tRBeVkuglZIjPJfTmo+y8osI1Bs65x
muGdxGu3kO0MkwY4KbVi+MkJKE4us6lJGoIn0/XC63F7WbHx0YssfN0oOJLV0k+v
mXjmlXut+CxaeRfhJO1rD1BZtDrkMpHJ4lzRlDz3QIPqYzY6AlEKx0mVXq47Gv0D
YV6XWYD/+JRvheY+BpNwbK4I1KrNmrfqfJUOi4vjpqND9RgGiFr0qqDOat2565Ne
5KEXejusY+Gn9+vm2jdw2AgN2gy8LYDAX2ChNMuE0IISXERSyxIVDgvegtGEj/xR
/4VZ3etjNZDrHVvVIBAcrDCMumgSVMikjCTPNiqpShACYe4/L7NiUtTg2nCzTOO9
ugIS1+qkf+Epk43XZHP4Cxtkuuro5e+sTCxeVvU12CkpHNUl0Z0CAmiUeTx3oT0p
jGWWWzzebo5cXMrq+1ZsiudOw3JQKeVnBLttnm+xIDOlqCisIld8HyTDxTUe4/hT
EMZL3TRNNpDFlwyeFj2H53fyhM1DZ9GyxyOSUlmLF1IW6gzb+w6j2L9GRr/zl5Xi
8X0gYSo0h2OWDCGj+TilAn1j72EmXoK+5mSTN2qzw65USFkyfDC1grZnS+56Qw0d
wi+ojBuhf8+hwYwexW60zIvhBo1GEBv7QrmPPIfTtmpnahjm9L3tio/HLwtNe1hs
mv/WylWifL//meN9HvpzR3TwJZ1mP/ewLGC51Ye4rluJxN7/UhYTPwKboE6Z9kz3
WKls2XLfsUn4KlgXBstLlgyPkUJ7y/92Nzi6YjzSSjitxbxsBYgV+/PGhjXgrvTE
heUiH1YUVRM206hnP3mQeQLvO/BdzVLss9FDda0MG/L2CxmS9X4O+VCNCH3bH27u
KnIpF1BbOVUkZSUSqim+pmrAPj9BAaNEGcxgCcwTu+7VSdxAmUSJLaAG00TqW19H
zTs0L81612A4uqqiDsUTz5oMRCnZlbaHtx1+L86Z3P2BJlczfGYUwtARVJunWqdo
qkCxCT8blwWLMEmaBQRXqyVaVUqUTZ2H49zZdWW0qc2HwmXR3BrBY43jkBwFJzwg
gv/fVuLiS4iNYVbnv57TaPIUYqzaoCc8Yic+73D4Z0xdMdGXyXacCRaxTPy+f3HW
YyEfYLykAOf9iKZXroQksLLLvRAglahKABntpMnKJnFmipai68+UYgL5pbG7n1uz
s43QeVbDT7oWjQPunc5Dntxm3eq34/wxJ63aO6BfhvcbUS1hmX7hgJIVyEq4dr6w
j9+qJJz3zhS/MUaSyKmMQqVYcsIWKgHMeNP0lhIvdj+oycoJcDsu2q9uV4mNdcyN
NeqpwUS62Do3adF/UKgIWSKGtQeUJUwe+6a0RjWuoPjnNnLd4Ncg6ss23GbUvLhu
+6hbo6BZkNoO3SGa6pMl463KOI6M1LpAcDvhLql9VCXfUgZ2W6oJp7FMecEoIoMW
lCcG1GY4PteikppNiP009VvdTAyO3XjMNMRoY5QWJEIT2CIUoJS5pMSrsa8UGxY1
lb34YUaF14U6lgman7uZQINWDLQij9zk2wZIjFgWzm+/xS5cZ0irc0+qIvlLjL1E
khWwT7RixaSVDFfxWlwHAJjoU/W2UnCYSVxrAymd+430kh/wT0aB2r8wf4W340zO
p0dzEGUV6bfhmyvhYY7lD+zyN+kYd6d0C/tgvYEVgi8AUy70Cb3xMKsTgG3MRLLa
xEcdKqOK2DymuLsZMZZjgePP0Mk7W409maPNDQbh1+QpXryEhPmuPJkiYxQChiXN
lXoKkmfT1qZ2+AGw1WAgy2+DdQGE7xWuQrItZHZEVu3AWIIkHagKECjo1Jt2ePu0
xlRH93aumNX3p5Dy18joo+CuBBrfxNrn3Si9NBkCw1pxciytclef8ApoLHFX2Zws
meVf92JLF+f9PdppCJLHOC9oAxVhMWv4funqxvFVF5XNvx4Am4H2CED82Bk2GWvx
nkV3HwYBfL7eaOjOcI+n1uzpM5v0dHNadutgzvHk3/9+jp000lsWtNr9/nMl++L/
jz5gS0LXaDT4gE86UPFCrokH2KEPKISXP5v2uXv+9/Eyd2ofIKlpAXLuOhyFW0df
jAamwUvGq9q6hlF4E3h+itCRRJ3YDPNcob47g63P/ZLoUNiqqIrUIjEcLkMOnqEo
Hq0fQZbksy3R8LHAWsJdeI8EOPzGSpe9o7wzAusRX5AY5eYVbv3xxkcqNgnqqMxZ
a+zDpbnDa/YHYrcmMZqYUFTBkHnduO4QhJD91ParVSGViFLWtnZS3tza8LCz32ER
ZCwS0OnXzG73dd6qsBb0B/c2qVTbPw+DwcRGDVtF0ZtHE4RhejGBjWW7wlLZyLLf
ENcVeurNyVt0V3IDfhfX9WDEbRKkHR2M+gvQPM54J+dJ9GHZpeRKiOAZTA9XYz41
pMM6IbJDTmuUQvaENCumo8Buc37VypLSNNdjKxJwFVEn29GCtJ/ukdIsPklCICnC
mYO8G7qZXY0rLSI2ThMY8nK7sMMtw0o86uXkLLEeBoYDiSK5VryliPwqy17xciYy
kaFPTHLqdSMHsxYuueXhGLF5M7nCawHuNGkJ6/HFUSrnb5HHBU7tp8ymaTqHhWkc
OR14K89v6yevuCZ3N/fHzdtw7qvKUWHjykCRvoi5j0qVbfwHH+g8YLF6TmuZMsc+
lhpOM01jaZjGyFJYE5KOaPzhNYJ6UHIarfO2TnM7lR1mIZ7ybYsfZ0ki+/uVOGD4
c3zl3LRlxo36ghwwBNr/iSzl6uc0Fr5/pw0W52HjvYPXyDaUTAZA6pxL9qfl8lcA
6EKzwjuRW6Qliz4w2vydzro6+NVgoNkQtiO52exz9Fi0t29I9tN5SzGnQQriYF2M
u94SKOxsPErCi77JUA+ysT7/7+Sq3Sr0TJlqNzJFKRL4OkB/vgdrbmHK06Km/FDb
7qbuir+NwGv21yWx9hqQZwpK/kuKUG8qmEgySROHwcbDC0BD5/fUfu+9vdh69yJs
14p/v90Le/2vW5wmmtSQmj4Fh4uYnqXxYFndMP5Gg/lH3sqcrxlI5k1VyHtK0w6Z
qjqqVK7JNqKZ/6SaZT400MnSr8SD7JeWajQTByW3fjO3H7haWT1juglNMwKjK397
cEQSrHOgIs6D+lvPV83BeXQtUZnNQNzdf1kURwcj6E2G2cGzA7VS3OFInF5u1+PT
/MVXP5Nf/K2N//g032BYRjRSJR65kk/h3MdJba32cwkaS3F9AZ0jsxz9LydIPL+o
5JO+cAnnj57FUg1bJUH4UU6Dsax2O90y1aYsiPlo8g703sexxH1E2ZZ7HObs/Uim
3DbNS6+W5AGBomBoKKWvCtZuxc9ew3vbeaJpgLLjalwhaBl22Gl2kMDkCXGTKZgX
5lvnJhBVKqAtYxXdEyMKNjrVKMdT5Jhv1C66RCgXHjLzJlPJLxJVn7izxaiMBLT6
BFR5801+aG7D5c9emARowregw/F1g8kOyGNMOHARVd63MUyf4bomjfsbA4tyRqme
qgtQJnovrL3LaOSWqDrRZS0wCZfovWY9OKe1/7KexOhZQX3miitsJeH42DloDg7K
lVBqLeiJWq3E137TnkXeHiopL3xyHJ58NfWbosfjn8Y5IrXnb9ainYnKc3uuRk6R
dbu6DPUBXr2koHE3/XF/pXY9hqx0p0FpORWgcyWb4lrVhJEuX14iXxoCvkbp2BcC
P/cPNUJTA18EfUGq7d15ytIDyR99UY4HYkJmXy6ykwH2Y1q1yeMEy93AW6RRwuWn
iAudjirptNaoX9MxUsIgfb17OiqPx2GPDD37xy2Qgf5QQfbt1MYNzcZCDocUjMEr
H0zcEh9NvyqDInhK/FYgc/uzSmR3NiB1U9RJwh+P19FM/apn5naiiE0iFW1UqjGw
EybKmWvFPz5DZmPwW5iEh/LaMgrZdEHVpX08p0jJhjMM8ghvxHWi6RiWaRhCYk6i
OOXtZzgdBK6lucd8UKdJE61bLUeBEe50ffjgTyUJKdQN8mQ0T1W10Fwk414GZTME
aERMdTHH+/V5mlmn1oFvNpw0hoWRv4iHnobNrYzfqup/A/FuWx0+yw3T0XGgUUtZ
8L/DROhs7XTSepOPRMoVXFmsbkp2zxhhUxlVzEMxtVNdljAQW4plEhUIZ8S31uOf
we8zwFmt5hm8WU8/YkKB2Ou2LjO0TR4svXXJ/q8l07dlTkR0O8ag4jewI6VDGB1O
thp1FHUJxKBpbRBxdQmq4LKPYmNYwluTIIMZoV01ajPqP2cbsxuA71+QpSX4v4sL
ClsIHZIBiN/af4+qVePsIKBc0CWkHtaQSM8SPhIdqOxRql8J+xgXlt3HpkF4ZGz6
0Sm8F/YEvU0eTFYTTs5FkcsFVXZiCim33wRhBLicmGzMncgtM5pDlmSxKkTBhsHj
XQQQPX2TW/Y4LSmAAY/PyBZiVtxcsHHOCFDaUvL0Cmk4ls9bberf3w2V7rb72TPj
Z0I5FzxWpNFEchI9ODBEOm9KYCzApv2G5VajZ7LBl3q018HjGp/KLx2i5xKwwlvF
OrCnfVqSkvZ9A5Vgzy6cOujyvfk5+YWLREVwrbBqqablyK6cYJjjwuwahpe/fwjK
fTlbfGrlRSwJYSK+GdQIEMrJlOinavgtGUx0hnnhLcx6mGVN+Vw8IUktSgutekam
T/V+nAw+AtSqPxNPl5gPqkrJXJrbecCRmjx77EWDeK5+tzFdOI6nRMS1sL+wctq3
1nTEa4vzuqrTb/Ln81wDEQ4eMbD7zFr42shVy6gS52W4RGVMKdecuEzneOaaUxkK
eurlX6zF93IGrXfxyuimrr1beGA4FO7hJRZ0/vc/HmXxefdE1D611rAWBq3VJZJZ
Tpn0OqpxDAL9oT94/jK/7PInnKfyv9BW7pg9+oBv+LEUVBPGFAWg1sOeAqmDb0hI
s5UBgHnI5x8K49F/uvMnP1+TE7Qhuw1J3vQ+Q6XKSbsVziUa+s8y6ehYs6q7TkqI
Qq9jkfRWN8Ahqjpm9qUXuxxGVKd6PMtdwOKLcJLhb7u8w5lljUMeYWUdOZm+tuOS
FdBHIZpnnFxcHOL+4LyGML69ZWA9c296VQ68lFKO+Uid3eLl+9ZUgrbsv+F+l9b8
bN3vbB0bGmkE5iD2YdxK3r1gmtJP1qXk8Sx0D3nfWmu1h5MCVo/WrSkPpXmlsK9O
90DK6kFVTp+aT4K2eONbYFEzWU9cFvElW9ui6ZCtU089Tzmd5hi956+hSkCZtezp
c5HzlaUbikJRA82QOG6XJFOElOGmdNwTB1RefByNeah+iI2IaBd66/DjN/sN6/Uy
DumDNAmVePVcw1qmD4Qe7m2DCgY1NX7/UqNZd8EFpgbNTMjpL8/gEZCll0udUMqe
ipyzRsBxnKHNRngX2I7r0iO44Mx4lJtnZPDTY/dXArWBhULX3tZRC1IYXfM5sSxH
k33tALYlJu1jI2NsbYixlv8wrmOoebHHqlHKnv0ZkGsJpw6SJ2H9GNIrNWHlAJSB
IXQvOPjPLBvyIOo9gXe8aO9UbnmCDl1+Co3PTnvVe58o0LtH1vCDUFhHKIuxqar8
SxEeufFk8if9y1qdyUtHBynQDCy1Q1rLe7cseFQcqOdRbOh6spUFEMc1SeeeQ0kg
U9zEAaqUONK/0BpycZOvweVWPN0Ea+Vu9e+69yikSV5mTBetpOaSFxBRMXEDT/0R
6SuF1VlpzPgMtxB2EAhGzfeduH/5makNNDGV6OAYhBA+ttstZSFqQlgU8nAQABwt
dtEUc8eEPP8T75WHowLa0KQcSH0UfnhJSdRJDCRSU2b2tBqO+3XcW8q8iWntCSUr
MejawpnZJhDY7dOX3yvSjOTKd6Y3JRMK+OqMotL+yamM5awqvdx8sA3rhtxOCGkD
CmmmjLzBoDyT4LOP4eW2kwmaIyHjsnGfmFdxrk5xltZ9luRw74onGG5xFig4nI08
GBl6aaqFK1RDUFyO51FagZtekXtpgd3QQyqKdSPiQ9P4CE47aOHp2uu54KzURaKs
oxJoZ7F2tO7O+2B2JyQMSDGAcqLkYYawl+RRmhToOeuPoaZPlWeseNTfnvo9Cf0J
pqqbKJA3WKajaEtJM99Lmwl1MFZOHtu637Guk/S5Ei5Qjbtrkp1dXtS7m3hcq7WY
O5TYMu8s1UAAX/eODL19vUcMENacya6GgvYmqWfMGJiTgjQ+4lft2KyceId7ctEo
ZmcNZ+VlCbA7TKNqI3z96PST9Rt5LIQ6Q22Ni7vpe5Kmoa/tIYBafgg3dx1Hx9Ty
h6V8bTpXgkxymWsTITSXvAKre2RnVNlPt5VCw4E1GhlsvKl6jarfMb8Q4uOwJ96y
oxhFn9d1B7yZNR+0rEGs0SOdj+cuMvCnddToQhZzZkgFDpxqwWGQgdb0lIRaXIF0
RdJKbhLMF6O/7kkVW1Ybyc4FGNRq99DSsydGW+StQSJ7RlDqNKDdrT7Mb9TWTx87
IouwRSpQQqlviGge4nEVY1FUpIhLVF/VlSYfOjIFjDKFVtrvh4es6UqOgom12zHW
FE3Pb3xNZGIfOsyl9C1DeF0uxmkLaItZI19MQiT/K/WHfQtv0QDWhRJDPFcExiaY
WNB3ICtYAs8ZfLuXj6KCBxUXgSAVmKvwknOjIT1VcI7aL4VBOkH/H+eKY9vG56m6
CsjQ7Uq5FpG5M72OVAMOn7u1ux3I05N1R0rX4FdVN0RFc1Z2lIOqJTxRgg5jE1ak
MlMQr1CO+FYh4o8NkNKL/raWavhtOfiqO5/MjoSZ9GfVCbiekKxkEYxsKKO1VJCm
EY5t+mDFIcptMDeehHNaKyE3axFcRwMwGTa4NMrSROwc5JWjjL3WUywfusENaS6s
AtfTVTKZbwtzkOwld3xIWlOu6WzIuhHPou0x21bsFDDbfa4mjY2MVIa8a8cVfjSq
jpvjtQWeAu1fKBFOFBqnHUUS+wgEbveNUF7yCom1NLN59bbQLB8iyQGIGTKXi7fl
N6luoiq9LJZ6ov5lh+csTU9lWD7CnEitpAvWjpffX6SKwksNkhafUCNYhvEmvWDT
vMYG2Giwr+e4+/a3PIyFbIYAgl9clgkQAcchfW6RlIaheZYCdDgPTKIJ1d2gF/kd
h29rC8v05UG9e2EoV5niyJZ8L12TsrMSyi2/cCVk1UyBL+WGLTQR48OJauFAyTKr
Z8LLS9p77ge4XSvbBE/afU9/EDLdZyLwBuYci8Z52NtpKEKrDJ9PurB0eQciOTXU
SYyu0YTZKXYGc0GbCODjdamQCminJMj8Jz0q++8ufta2GUEqQ6reVKlv1Qc4qv4c
yal0q2ddDd7VJCNmCGg1SNCKVJY5NwCuK7R3CnwTWf1EzonQ3ZSgROtegKYKk7vI
dIhqqPDhWPpgE9WEuzFAQCwiv3ugmsfHZYAxa8GXBcnYt2FJprqLYCQ3dMebdMI/
HL8mBnX/cruecMtOpVzlRtqE6fHmngf3EFpo+iPu6wLYPkdgkqr+QVR5AF+ohUQU
8fA3cBWon39NsGX4TdQBuL0KeAzWczUSzCeMwtKei/rwi0I4hQZIKNZHUwoSOkWt
AywgWRrC86G3nAlgJYBH5sTHia0eZgXB6/jueBwziqIUdzbKtO3L+LZteOwXXMwM
iMhi9vEA64BZX4aQJfLvFaG9XNypTzCrtoNK0TshAkmkraULIjQr1Xaakh+lWTpi
NO08novZ0kWgbcN96NJK63lbZZv1Fwg6qQaTyWPiLMHs+P33Va//zNFWhQNtTLTb
seNbbpYLPtvXW9vEFsWR0wqvveq8KwymLJA8csZNUqC+fdUu0SBd3yJ/V0DczC2F
7qat79UWvVuwOBPd4q7IQTGPnOSscf5wuvIZgq+JRjbgFatWK5eQgwFEK3mETga6
RCCfDT8F/4gvm6kFD8lQYNcBBElJOGQ7arQQy1rgWjt4U3nLEply/UJnHBsGmSzJ
9wLsGUrhgbZz3YpHqVWmwpQU1xp9FiwO/JlQL+N36Ks1H9TChG/+AQiVcgipRwzb
tunI3hBEM40QzUMOicRYN3LHJZVqDs7V1MhsGN5EAPIUKsg2+b8kfj1PaaoK8F0y
BHowPdibuL0dtgUygAjMUJh3ytkoJQrbDaOxevlDnDLh9m6Pup3LZSLJUlTqjQm4
feY5Rqy7G3PWSw+0S6g9NhCKNwcq8rXuyFrWIcrSPqcuIivFOSFdNSGu0CIvlo5O
q9qAeFoZ47wwDF3a+ABmzA8806j2QcNB6xpkjGpY/cnI/Y+kBgx82sf1l73UDhFy
Y6cAWMVOfHT8jqxiGiHIlva5AOV7Hr5Y2FxumYPA9/U4GvKjPtniV1hq9f41F7xt
5lxLnhlkibV08/sFWJU/HZfpbT2bpnbQTg9+YfmFcVLY/XWZn7qwjUZs8Jx+kM2+
RjL4ulc77D8l6k/AQPXRC7Y08ZbQ8Fd8CJ//if6d1iTuM8R36zoHmGBN8Ht++eA/
27q/M+KAvmS6AMIEvqCYxCuoTGsQROY8xV6c7Km36KfjwTGSr6rpsOkh6TRqzAsi
mnb/X+nGgmfoNpBxYavtvsvI4IpLMx2OPKU6Y1SMQ/QWoCxpC84HzhXHGvFp9EmN
yUsOW6IxcWJ17U9K5MXinH4ryded5SQo/I2icV/Zt69Y5A5y8Hfgewuo+NZ46+Sy
6H5s72hAKaJZ3/+fQAHp2osUD2Jyvt07pcV7WsxtjBqbGAGlIVv/S7nIX4BVvsZo
wEIEbOrUdi3jKmTg9Q1zmTLgy+sX5sq5S+W+ejdIOTTnwJrtYlni0TeBT+R7S1Rz
G+xi6r9MlD1o1gEz1iUjC+YHUnWaOsOQHR64CWxeu4+rJo4h2AaMKUnEuX8y+QTp
czRLrIaaXO5m7lu9UxMYSqLok/H7LGy+iC5uhdcJ/9kPrKP/yjVYyDHogVFISfvi
t4QZ695oobn7uqG2MlJ4B/sqn1c7A2d+yogaKzAvmaoTc1oGLNhTFIObsN9+DwST
rFkKl4naT2hp53UruoGZeD/W1FxbrpgYxtYJJ3XT0J4Q3BM1hDUt6Myz+05vUDb6
aafD2BrV/TZc8cMQkFZZcgi+aJs1LlddOiWqDG0KGcpk2TS7UZsXYBhZ7l5j5loG
EM0Zp149eI70gi0VHAps/qaQhTRF+ukCVvXmeSyFF725Mk4+ol+gzSzhnQSlWIFl
U5KO+6o9FfVFoCelwcwmxbTicPtr6kfWPfxJjZK7CjBqMqvTv0L3CoLJwJOj5kXj
p/M5Dz9ZJJxI5ZkokTkCWbcARnD4Y9RiKdy9QimCbs/Ktr87zfkZ2cVWhggNSHEO
Jx8Jak7aptRcJkxd/LUnMO1tfad4GQljJuVXQ8tB+EPen9BjsvJKjioI8oc1hGkN
wsd0uScqmMWUhhnbRlCQhhNcAQcAxBArGhzoET6llzD1f/CCVJwpRh4x10fEr+Zg
j403Uin1fwlgb/EdU/+Z7iQFLCcNFOmeH2gnq4E8n7DKWF1ixmoY5h9wEBx4VXiq
+tV6dkJ6aV7Dn+inKbwPozfXNxNYezk/csxkjpL1nxkQeILuoQMZRaOaKroSF9In
huPN7Zvo79UdxpZsDo7DxTqGCKmC/YpNiYn4qUebjr3aqMkQ0jPuS8E53kmKjGJC
LuCYX9RIjuhWjSkXO+wUKmgD8jdLpEVmiAAFKwz/aPumb/HPVa0Y8TY8LrZ0WbPK
bknNk0LK02uDTArhCLATFi0o7zsxfg/SNKKy7OHbRKL9sxDNhgacxCaQTkDpTwcY
KFDowh1BI3lvWzAEnk1P2t4LeKGpU0+EzfwmREgATXHzdLEQVLPEISpueLVOpcwl
ubUH087HJ7NgWJ6nY2z8g/5VeoJdMWUehU1ydsv3LldMQkoabNCMyKPbXGb5i+wS
KoHTFzMnbfEQKdJj05l47t5vjDWelQrirJwxyfaLcdojk2b+18RFRVM3ILfeq6Fn
f/QjmNOmoxL2f40NCOQMOaeQgBk7GooYZ4z1TVTBog1A+nNUhQKf3g/sE1pFPNcz
Lys8gyXkR9DGm3Y9CP32D4N9CNmPL0ZjTQXEL70IpviIM9O5x9tmzVoq17YvMwkl
UeOMQd9B4EmZc7Wb1mPCoIMnjPmq+yVLGIAwpfMKk06gPrUbHcCxTSKZINU06rMg
9OZuUEA8L7LPLBA3WCwJCzGzPFQHSolQPt225hUGFSvxEzU6ADOrIK4WjUcbXo7J
Qfx93igiEMsEFA7c9hWPcBtP5FiuMqNnu+R/pSsqUqjbTihdTzcfQbCHxRWuLshi
+K12qHkWpTsWVSLYpWXLkcB5oph6cbJl+LrzvaMcbUwnpONJo3iT5YTU9e27wXfB
mAlcVNBNCSsLCmRkHwuZEJIq4XKdEsIt9rO01EaRnCycucRlAk044BnUBuFx5j/J
1jL/oemo80ZOG/EJS5TtEp3zTjYfo4ovonQQa4eMGpPVQCRwB621MEvJ2vp69oUA
1gmNTM5X/g3QAZga/Q0x/ruWsxpdHbiqJ54M8KZp9umJ0wthOtRaFczGlWXyRL9s
bUFpvLPXxuuzgNB8Fbg2lbpXMpAzrOVYfrP8bnPLB7B8cOE+mAgQ4v/MH8J5QScb
spcrLCMfB5jWiYkmoEpl6kBNPQAvpLZ3cB7bcvV0r6gpfzvPASsDICK7yFyQ8V5E
SyjQXlDga8v/mwKX/56mMIEzPN1zljXVRJB++x+Ynykl7GaR6xsPbyAdDEJscwxg
Bewjq9cKaW2lELuN5qsn/yz9rcngkPPqWchHoELeaJSLBYzIBsLzoU07/73JpPEd
If2ePAcT7BDlRQXUbpq0ij8YlWBrZxiFZptw6BAPFptf+Q364DtchKWSfUO6yq+6
epyJxG2HZu/2EkVdURRL52JmEI2fazef4r9clf8KqFaW8CcUgbaIGO3vnJw+05hq
Y2X5hj97n5XOm/e6U+CGv8uu/zRsHkqosvhr8W+z8aM6zVmK1Nn+PlGDr06ElD8W
0tc8ooz7vjR9rX4iB9dlFqVOBDKyCW6ojFCVkBOimQOAWkl1wH8TZdIr+RvFLtpX
81TXC7AN0Qr/vvUaRUmYU9SFvuAXcgTxWKKCtSyFy2oZSBH8PAupy3br74E6njHI
YJHc5OBt/XsxrdZyhbzlEJsdjWqxpFqyB6lcjEqTrBobUS31XzcaYRAFXxAC8D1V
/E/iJMa13LX54f7BDC3ImBfa6xlSmS/vVnZr1U4CxxBFrInZxjRFdTTcn3m38V0x
uY2rSTO0vVPXcJcLNhAHmy1A2k6gNmMuNEN/5pmnoi+huoVqfl+hVDkyt6+/XNqD
J6Bk8Omc7Su+dlObGcWvyMuDyPH1/xA83XE6lU0PxQ7JAWsTdNj6Rm50SbHMa4DQ
TGixPb+aHjBpnxqyppuuxqhSJZtSjqNerjXR3IbOqmTpakxRwqOgxuhEVgtTKqOi
M1+86ZQm5frfsXZWGTzymooUuhoM+WHA9HWfe+l55HFrldr75jzJw8C5oFhc0XRq
Nej86DD5rYygngFM8bZUxlK7aHdfX3XaAOWYubpbwXVxUNHi0yxdRLh5St8XMDMA
KQ/nf+IlwT+M7LPSsITlPYPsJi2ael/2uJfc0CZ0wlsu6MPb7EPomWV/Uf1aF53P
bnUOJW2ijMIZ1nAi/8ymh/OqrzG7DElbKs81KjJLZC0KPCyjvcrjXFW3hF4KA8qC
cw96WMm1glSBnaVQIGDxaU4XwU4BA+67GSTD+/NJ0qp2u+D9JfQUaFZxAJeZ7M2K
2PiIoi+4Pd8skalf+qvb38wPc9NllSWQPZRHpEaZu2vGV6+7ZUIm3bjvSjF9hkM2
kPmI/uVSieLbOut1lMm+cxcjt+u8CNP9DeFQszU2wlLdr3AUp3jv+Ilmr85hSTIe
DNf4LxfKo4KJw2WWoxeoCOx/A/apbtMNbi5AoXXB3w4NvCGFP5zOooyk3su1lzMU
seU7Jryg7Wu+ntDvd1k9i/rBc0jsF5O5fkgueoaD4G0m2t/SesJMl6isOOhVieVR
MyeJHaor2FWNDiSGrYgdPSUDEMunha7sTvKrOYl4Z87Q/OlLH5PWpnH4T/+69mU8
i1u18cipV/PdLjZuzRnCrn0BBgDU9q/5Z0Q1rumOiwMi9AqGdRL1Y/5tcWMBOwzA
aPi/55moUdiL1V60xRF1ep3z9QpaMcXQnCaq38IWGiNDLEyXAbEjFqTjHO7LfxiZ
qDXHh2nddNfiurLCeA/O+SJwmhEgTEDvbR8l05XLKCCaMKSMZw3yuuYDLNmC1ESK
w1nkGOjOYJusuO9p6WAgGXzQBttO5XGWRM5QxV/AwERTrxbgkI7rMYHDbArg9389
OK3jvQKHOce/wcou75FKGH2HHLt1/Qk7qBH0FrwTxIhVsDBN7J5Nh6V6e9K8wlhq
iAIrohjDldasYCCgaT2oJEspZFfbLnTqhvfrwfw4D/iP1sRYJ49jhEKM7EcYMe4o
R8fOyFRb1l0ErgGQ6Uzkzh2u597uk7UeF/FuDWzy+Ir1ci70Ewzn2kUrYkwr/SXd
NSxKSHIIcxTUS6qa/8fSWyjbvvEL2CPFM+s0m2Itiy+VSF4xISt4g36Dj9Bgt2gn
C1/9KDpZdtWQwALAFLWAihTqDUkBQYRi84zaNK4DCZCm+1WIvVdeNgB11ng3pYTw
/ih7f/JVO9QNXISLiVkXTK/sSeJ/7WRnl8EMM3kTW1Jq5ZPdoctTDjux9k/HZviz
pU33e8Uaal+pkPvtY6i0Kq3dqMNvQouUF4s3BlsdMIhQAbzhRKBBssOWyzitxAoQ
72DcxGisJicxeSqdZ7NxznqBh35BbxHrPYyqhIMg3amuRYiWibJRBI8r3/gfzc7t
W8f7OvNOtWSndJgbhI2YXv7Lgb8ynWHkGQpAz1wM6s1Zcxu0m6m/QIY3uXxiY4Vv
cnQG/ADGTwBzpuLtioKq0XEdhq8n9pT+fsCA6xBAocPq//qE4KiArTqXddFhmoJi
OWLw1sSD3BK2q9GuPmB7dYppSZU1dC4xWrLVbrhs/WlKLNpGqsDbCXfFxy7PtPSY
Flfn1ySVRJO+k30Hr3Rnj01DOM1JrA6CNiZJNsmrGz1oHqdNNsYeWRqhajoDkfWr
Ctb3g57BUNYE9SdJC5ZVSxPCDe1MKcZOAreO3dBYZ7b4Z6JzPqKkEEyiFgCEIwCP
99qQL/4heUskGHHmwnaZzh9738SnRMANHJBpgVeZsPaOg6nUQDQjcebweiiE+ycA
b/DfckKtZYV0Bsjrv70Q1jefRSYhn49edjOKRwbQ3L6jiOC2vWj8Hbte8U8eGXKs
GwygtqNEEno6uU4CU8oaRtRdiiyVGO6WEFTKcOTaDGvloLVD5TF1H9rL/fxtf1su
YFmcqkY09EXk5Itjd//cHOLlXI0yhuqn2ojEoBQvktiHTZBdhWeR5rHYML7HvHAY
mJxyN/CCsRvdFzfOwtGF8TPB/P04E8TSq6Cv5MgTTlE8sSr1tEK5/IZoXp780l7l
fwm6d5IQ0W4JgzDluFepURlZQ9Pd9CY51Bei0smCLJ96zHLIC5kFo0uY4sGVSY/3
px54f2saA8/HChJp8fJIaX+qK0jkhPV2rEaCDEnpYjBPaWFAfO+RZSqybOyJeRsL
W6koh8ODazpeNvweR4oKgnVxBHyBoIsvgdosf+iA0aHn8hIA2Qd1XHUQI7CZLMI6
ayLhJ3RudYXpFQUq/eVVmQo71PWss3PUufsQp4qjfqMwc94KljTSKHNahEHPSe+w
w/d6nE6Bb2l9W4tzj75kEV8U9qOJa3ic2QameE8IdcphtNWndHOvT7Bt9VDJxRfz
xDxLwtEItf1vxUUCa+2jdiyJk8DqzjVdRRYFhEFglxaM//6PpKWkTSAmL2JNgu6A
m1WcfE6Z4jSC11uzkNMr9Wr1apPUidYLCTbgE+pSmJDZpBKgmKrkl2AKUs7e76xw
85iqwSxU6dMY8R7h2y+lqDYgJOutcoCmwsHDP8PsMmstIh//CyFGHQcYCiYwn9FZ
YrDWDhPNCajQYRufedgi7bBOkGsUc4guZ0e8tpTWJUBCJN09vqpHIh2VbbVoTrb/
t0YjnSh7DQHchIajdVQ7wIHy6CAyIZ46ljdQWoQv98Gb8KuICENhm8xtwRz+ZunM
E2YMBKSY+PulJoUD1P26S6/xaF9GZ0vEtgJ3pecwnqAXpr/JDWN51DOXpwCY7Crk
j48vmD7rsRBmEaUvMgY2/A8LM7UYTFTQjKsuNKonGJ+4aChCd4KHONpl5GQLqEjD
YvCseFg5rXlcSrT7NT2aDk2Jt7ZtHei0myHRU4r6aCP1EUmyuCDqDxVCv1tv5ZPT
U87VRpWCH05HQXCwyT80QSJtM/Z+cQDQWFL0k0N8HNY81SRzgnldWgKImlwI58GJ
sl1LQfN4IAX2gYl8QosZfhtJ6dlAPEquqy/by6aRV2XqN+Lu6pbuSD+MOMy6OsrC
n8RcG1C8/Pk/s68hTCQj9Ra32RJlHED9K99vqkK7gPSnIWVdtsxcJOPE7/o7vFfD
CyEOrus6V/6bFeMkv1CqXPQ4jcYTqFfziwX7Y/2pLFA0voU7jyda1mhiPrb8Ug9q
d4suSb/GRszwUMvXjBn7JJLcVzJC+7DMCrF6ksFosUPLC0tLkB+A0izEOfrFHFRP
x3AfY0nvGw19m29po+20czuw9emA0i5PK0LwYH1y8dAM0I1/t13NUNFaUjE6KOhW
kEdvumRS3ni5Ue0y+0hzGz3uilVaLLTOn/07WCpNbpqd9VWa98Rq3acWdm5SRGDw
2tIJ6V8AHNQLByX0XeDwE7kEx+Eqcq+RtmKqusbaaoGb84Uz+fRyFgwOufgcn1KW
p/imROP/EnCPjMJC/WO3o9/QSMWCfhyBTOKq9NsSaogqRvHxgo28OldDQlPos1pg
PIu9zE3mQ53HH1LEGKbscTUAlCJ1Jf6vM1xx+BpKfdZW916K4zRNMa45rrixOztj
WQg050m47tzKZji7g6QEN50ber8oT81f3fick3ztQZ1Uqc/EXrTruwsWmE1xCsK1
49jOJkqJsb5LJwWHPv9v4npqAdYzVbvS4V//6CPBV0xq/lzecrFaQmzV1O+e7fXl
PuXA3LGEOxWUL6BrXA9MQOZrurBAN4HoTmC3mOrGyCXQCk2A2t3HrhiOW2uWtJWW
VqGj7zgVoZXCRbBSe39urHsB0MsczC+nJJfV6Ipuu/CiiMw2HXJWp/4qqJQ4xiYJ
SXCaR3+IgAmDNEOjhlCaIUOVV9mClv97UfXe9FeeCyUBNz0XekMxO/tNR3E1owWw
ZwsuYAqqwuMHS5UHe243iGbVN0wZwWygN6oZu+s1z84JIQgKh2oDHJN+cQx/OA8G
Pd1gLl8ZQM95sqvSXc8xSEpRywj17iGuZB6j4aFmMxtX50aMd4aknC8rVt6J5nvt
xMXimCg2dq4r0/KBgIvUfs5c3X2uxkdsP4ATKlx0EtrwRNfehUemPrWxS4TnDTJe
Mgog+SUAzkONhTg+zWEn7fagK/cKBXjNNVNnEhwiDnfGL5gkqFc+Y2Eh95dLDiHF
Kmx8phaOgvg7ekCqwzP5/71u2BRZ3v6MxLWJF5n69k30C1OBFeKxDUOZd+TKcTbb
88l8BvRXhLNwdkSzczFOi4/rarAMCj6FyBX86PkQYGJYKw1hkINTEOJqWI2O20N7
lyjt/XEq9LtEsfPQsBGoVDyZCPwx9oIjqqI+G217YQLMFq32j8TWVEEdINWQHBXn
MsQH4qv564xOHAHMYOBKWF+JIL3+zwszijUTZIR1dAxutKil+APPCY4ymE/w8cvz
Y7b5H5svAcA6zoHOrZXzYYCHhF4OXoxP2URseYU35eGuFtjhQ3347rW0EEJTJcyb
/veiCVNqCFbvLd5gj2UWv1RXOkXmC30GhPmCOujsnnxcKrys/XHSxVDGCxtdjV6G
POIKGZdIUvs2Sm8P9X+aFVyL/bAWJdjZym9dF3RR87NzKWUmWjuA5XRAEhpyXi6J
5p5SOqChCxnnnf+5fOe6CWUZm2Zs9fZmp7gWZ3OkllNzSJzHclwiEa2q0i9+7fXl
004IWx84rkLo8vBBklkdCDH1I/s9qK7m8hPLIY85+qaFYaU8B4SgA5uy44Qg+sTa
K2GwCJ3udwtYooUlbCrEPdWBHNDNBK/VyuIw8xwfOO+d1OGQ+wt2he9g/A3Iz7Je
bG4TUcAUc3ewoN5PD19H64f4Vq/bNV3DuN9XkY00UjdbdxRGuR8dtM0iD6r0gyMh
uTHT5LtyDsSsM7FbZThZihrHJugG7oxGDJIXS7ctkP1x5kLl3ZerZWYzGzfJI+qP
4IPWCogqJ2wEYoty8NcVMpGerYWEI+ovnaqrUyamQlaGX9Jy6BQSwuUAaArj1ffk
c5Qcshx04DNvRyAk4+SL68iZ3JvHPLpsN65WEvZEJ7kHmaqfKdFKpu3HL735QuvD
mN6m8hDY05K+ZP3R+c1VNUYLh4JY8Qw2PN4dJ8sPtXPwliGFr/er3WW0fifgn/EA
uzXsb7zvAsN1xGP2rxP3ZdW8plWQ1M1E83rKP11CF2Uv22wsKaTWd3grzqOivM+U
UDDCrXvlFVGa3iER4Dp9JO8C/QpxSZcDhTB/OlZx5yHQTl9zL6sSxwdo7eMVB6RP
RyHNNSFj6J00t4gQadcnsZKHCqTU2YSNm/PdFq7eEMVnzTyuF7AmB4sMH0guKWya
J9Lf8n8P8E1P+Al12PFjF0Ka5Bar2HkXsrK4NrDHppelR9r/Yl71kp2xLOQgh5rl
vExwGb80q4abmuGDkVrHNdVANC1DbyePCbSiSo4YepnoeCpMTLXTJ6tgCPDPUV5F
CW6ICYjdRNBYPCfpgGDx2Xq+07zL0lVqqvRZJ6caz7mcI4JSC01IE3+PsAWmGvBw
4+6cEcow+r8dlUf4v6aAWWVhcffUkNtPZ8hgLkRZGLbJJxJY8lV4DXyfCD9VOiWl
RGa7wFEq/8yZFmNVNtO0ayH9KZIIXhzgJzQx2NsQSKklSVHg2PKIWQqSOMKO0dT9
yhfqZrNf7WthbeniVyADX6Kgs2RJvBEhVi9JniKyIEDzaPDU/sj1EbF6stq/oZKM
D8QotEarJ8T/F7btEZjqEuhliTz9xgN1nyuJKUwce8lORKrVYktqPEEMuQTpZGmZ
s+fs+H9rOVNoydh6MnVSRjj1ClWPIBvnz43SCgxhmLf1JYRChGb/c6QniEGWsY3j
jsqd05VX2ylryDf1c/NuF1kXpNRg49d0NAck5l8cMkXGvz4puU2BbA0muKalJuCW
MkVV9BRFDiJCaWJYf4ajcMndcHJVb6oJlywFWGN2QP6YwqDRQ4tJu1wJSSnketZ3
9avqBG3jf+OYenKhl7SvtQqp/TJnSfWYJHR6xZ0Jn0Vp0kv7++l8QOS730nJSJqP
pUS2JTBdWPhKDps2AC/ulC4lSb1uYx16mwMXuk1lAe/oQfzOTpYpJOmTvNXXCtOc
SSOgLh0eyM7g/StWtLgKIYgz9g6xUt42OBaUY6WVu0n76B0Fuhkwpx5Kxu5LznTa
ZwrRL+1NJgYvvNzRdpsL9kLj54tv8JWQ5frFwBfX22XwVlB3EiWIXYr9zz01++Y1
XNG8iSzK0nJjUrSn/lCIjBDKhMYcRbGNC7nLJRvfJ8uruIaw6Mx36cJYQNw4/jFb
XwKlU1CUFMd2U9/XYx1BQw+EJ38Z3D0Grw17mTF5HE5elmXp8joiZS04+4qQ4UaK
9OpbstsjXcam+wP8pMhLLl5DR0uTi9icMn+U0NJCdoEwHSzE9yhhPZt/0gQGzxBy
ngpb6ZeyblzOJEwAYY+LOdMFYJ7g4gt60WoTajqLojLkf95pJsdoxebKtJfmrPHb
lrNkhcIBidKwo/MbstsgSApR7dAYobPEIX9c6UkCvsAPnqxR1AwNIjlL6A2TNI4u
I2oo7AxK5duqjFc2PG+WjpPwS6D1YaOg+gLcKiZuKzWO5DbSSjtJpdAA2hixKAun
7PSn+uY214vQuz0rtiS+aHV7sexnXQ0hfgRjJpsxiSh9LY/kCs52IGdxxfKCFyGn
L5GZUm6wVZ8vH6IRSXh6kmudTUEnDbL7+DIuwbaWTAbk/9zusiLsqH7wm5Q5b8vR
HkuAILEZM0Bx1ua/oL7lgvHTwLQrNLSKmKHw+2coFS8jc/262Gibdvzx5isnHsdZ
61L2MkGUDbmfh3exR3wqwEHIRqau+kkym854phBDfAsQw0T7gyiHfSKFIrZb62uo
NtPt21SIqYLHkEsVIhxD7WcH75He9wtliJdkHK3EANwa+6dhG12A5yMOVHS3HqIr
464hLRYwQrtPPjBEGwdPo4qZJ4GB8M5cgRsyFvhWrFSPkJAJ6Y+oRIt5oVxSQ3oX
0eisYpiw4/uu8ojEvoZWvyLpZhV3/PQHVa3nOqB6Y68Z+W+4OqXonmhT8TgV4IR6
BWW7EOVJDsLTpTt1mVFVsbjEAcn0M15PcdHdke47SBTuqWUNveETNwIQUhPSIuJ8
KqnWHGLi81qxpP5qxCHHdfozcc5aADOqiASNWtXY0zLhs3+WqAC2BTmGXU5Ivwou
MWimfoTXnvIGdswxeAyFZMTJxmZmC+sDCgL1l9BzQZmQNRPecxs+1Y8mUv5f4nH9
SebcjVvPKWeDDlmZoUsWnpT/NI78chE831ghT/W5OQnp/OVyKF6mk9E50+5rpm1v
A61wzOn8U7Hvx6d2LJHoikxUNtEyoQKOvDU6jkGtFP/t43YgiGlCUigCkFhDUOQA
ll6WDJ81ybOm1TVUk0+zmayz/e76auk5XGM8BEPNN6XLm4XllvKLM5V627LE4hrc
vBwowTPfzlg/2QwNhn6vMje+1g3QKYMhqa4/T4kmNhFIf9nplGJM6qn2YB4W4jbz
ICqqgoQW8F6a9px+eJz7KuW6vhcnwU9alo4iPDkYKrWeCkIJqCmHMwgRnZbmhh9F
pD2QmpeHL/kLFOFLDrrFI49FQlcMce+j2dP6WYOEZhLFlAcA8cRrcLunjptCrdlD
azxC8Fl/R1TRS3zLCa3sDae5Hdlgfciy0z9uyDhLFmvsOEtvDcWOZHEXuo4YOmEJ
G7jR6JE5JoUAGoZXXj86BSmhqq4hpX6WwV3ZfkwmzW8S464+YjSlgTEM+5+4Olti
ykFUsvxW09Ot54Q18wai6JxXHaYCa1/PdiNEzpq3/BZgiqLyR4u30hCQhIpN5c8E
RjS04EP8MT75I4L7Hfc2alMm4mQkmlZcqbz8H7/9vEL82ngzR/t60DvVRZ+XlwDG
a1bilIfIgjZNcqtG5TDDhMIEuTT1IkUJUMJvZn0I9/AQikK/RA03fH8ta87WDJkK
uVHJrhHPWAm4WplDmiUmCcu3TGYux6x7jbBnplMCcmdzqn6hUSu8ptOXKOn28NCv
XFT5rpWy67xvl3/7ZcZK3IFBvbhWoLNXmvJ8JwliL77o5NyvmnC+P//s0YJIv4Uo
9pUDQtO7u6ha2Je4nYJDnxHFz1EoO5e+sCbCZjAyhQgeuRThI1kxCIojA9uB0fBz
qIIFE6pHCx5FKLC5SGkaqwe+sz89w9l2OEjuI5kOZ70xejqH8+8iTsA3CbpbeuY4
Cc+MWP7+uolaDMp6LQCZfMMVwcDleFcMSVejheaJAhbRFuk62BTHAgGqeRANcj30
GDuzPwY9GN1+n+2+sZcQKKMINgCP7Z4pLUk57yQRVD9xpSAyjGOPOLQgDL6lAMZ4
9gJiJRNDMFdjlyv1I6n9Hp/O0QGWOMPldw0Mf8r3TiFLPqI7K+t1ygkW7O8tnA1+
maDpRUPi1inA7S+cLx7N+a6Mhg7v24tL5ld3y5OymY9a18tFUjCrGfshIekMrB6b
bxynJlAH9bd3Ti13MUfVciP68q1oFoI1ni+hsoz7b/nz94mRJi1uzxFjHnsbK/yw
jquknmwaKl0BwHWfxlv2NPbZip7RmAUJv3NAaEYAGhexOpKU6s1IUXFceWTuQPVJ
PSzGV6ir6DEJEfkrZu3feGw91NlXrT/IKYoqhSUWNovXrXziybFiMcMzPiw8sdXm
AO3fq5Ws50vAmDtJ1GTbf78nCpwpQfqA0FHkV5PVuuygNsvJ6bEOlNTOxJJ/sY2u
BvZyAlWzUF5064B3JbRmFj/G70z+BJjxwM49YBls6mfbbL6Psh3GnzMR6K7lRB0i
SMvK0mMpg2YHeYwpflAE0wzxvCyqPNOlu5NtI6w5PBeIiVdP/oQKAih+YLn8jKwj
o0UfxZNwddSJbkaK38eWZ7ONIU8SzKODErsYIDVE8tBhlYH8IaOgqVJqNIzzcf0K
hziGM6kBSaJ3In7fU1dxXI9os7zAuF0UMdVo7Uk/rZMBjO10/4NxcFs/gETe0Yn0
bTPeI5G3JA1NjBW0wsOoxF/mtTEDUBGsq+otn28s+qZoVc2dCamKtt/jSZ76fnpA
J7uBEems3dWdgiq2yVP6fLhOrdsnjW1bVHF7oApsMUuZPGYNrbyDpFApRcIG+HlL
hkuzUEh3lcdQZB/B9R9NgoIqjRwvv3ugHhR7tE//Z1r1cRBY1BcC2xgrbWNX0MQl
8gi8AU3MiQkIqaFnYEUVzogIEa2zFyjIVPZ5O/jPTvVAf6let4lJLhvY4KmoYQmy
5VaDu0k2cIKdTC8kVqdp6TgEgbMqwkA85T7Z6EB8G/Zk++nSHj/kgIz5U1NjWqqm
4syg8g/J1EnNpiV5e5uCxMft++1JZ53ViYGj4nea5vV+yVVX8QQY/AmgPanRO9Jo
eT/IvyKu16DeVAkdb439XUP0Yo7h0xC3uZPxZaNOS9cRzwOL9tN5UrIPk1w2C/AU
Prfmwh+jdYt55SLTP1g2p5Ymh5iSyJ+7DwFqc1nRwYFg6m8nO/L9Jp09r2o+fFIT
qjRAHm0Z8F3EBpmsYawgkaEcBtdQ31h72mWprbqzEJSR6Y0RxF/es5RSEDNy3geF
Gieel5bKQdx4E7JoYTlZct5owaKAHBvRmahV6ismXKXHRYf9V2RaF2LpP4G7K/IK
75Ydhf9sXXU+O+cmXDf2DNOY3m3xUOxIXpXA47qvgIlrS+w/H/+Qhm7eGZbXBX4I
YCSXhKC5dgBW4NiWujppgyIGaJfIf4ZDqrZy6Foqu9LHPUi7e/8J40gbhj2LRJeQ
bWBPtgGscrCUIgyWBSiLV6TQlusn5qtSIOxxd9SfAdk4JkOX8BECrQvTtowHf0OK
4pmo7LFur6GcHBol6XbJhJqg02XdvGSLpA/qKX2RvLhCSzXq1HhngDayJNKbV+Hm
a39R9fPCd1eNdN5j1FDedLp77rNNAsYo21C3sleMbRdxvdEYyNo0t2AWmKry0919
1SqicvydR1EWOFcroT+nismzKLKpOVn/bbi9VxFjvhV8E6LWZejarbDqsK5/OuT9
rCRhkw/4VJ+ZikilNY7+MG1v5AEi2342MIRc0rn+c0OKMEp+Pl771BzKtdvoibDY
0+4JBU5syViRLrapRO9843czxK+81pL7suUoZzLL99saNXIqYIDn6tRkI/2eFIKW
bTjt72BJYh1ebsLkDDEUutf+56vBFa3WAyO/0PLHew7V0zZ0c4bdZHDLteyJq+9e
phpcoU9GwS8LLQBRk7vaVMUbJP/jclgJ7meXhKw3mMXdRdI6n087RyMQvEF++7qR
lTlgm0qCwudjpqU0cDmDzMmxcYsr5YrErl+AzltuhNzW+gmEVAwt+9HneWwAlFDG
jWRSWl0UAY2kc/M7yOAdRyLdlDQv46lefqzd6iPz/ZapYHxrxcYX40raA6bGsiPX
om13f3L+PqBjzEUund/F+PHIxhXMyQ9ocLQtjMaS9fUE/YASI3wJRWZ7pePh2jn4
A3hWT5CWMICFOEEjbGvmBClGacKw417IETKmv++o1BbU6fz4+lvpeRiiFXKmg3Nt
KNy38ykI/v9NcHOQ5ZFKOpHqK4jxGALCIeblCTJzyrSBEMHK9VlRoV7D7i3xGGDV
ENk/w1+6sbDruBX/moy7e1O7Suypom6F3yh446bbRN9HfngVks1EG3Y3DWHhgpoN
cInYoON4f5IXM+lesim7cJmgbir3u0pDuTeboreKkMu8oAVL1n6c31/i4+dwKIJu
Xein5inZ3/+uP5/XPdbYnyHwVrvLsc6VyL0et42cVo1otYp+JDouRL9S6TETQT08
89cC3F/MezCHVU9N3MsVLzajopBNdvyNfB+paDK2KBTSMvlTvBDiYN2YnlQRzh1y
rQYhxWzCIDiP0pdXlwumFuPweuuz+ICMBwRhPDTRc0z+8y8HUc+pKxjRzb0z4zvl
TXJrbb4M1KfIF0YRB0XOrv2RGg+rc3oncqMvdehKYcghQ1z+d79gL+Jq5OeSTmfd
EZrZQN+TQuVGffDNLgp7yf9scLSJBZmlTdEAJkvvP3sc/0CP8WVd1gVVKKey+2DA
zYZW1ZbKhwo97UNtwzFCuEINn+wneEfOMg5DPPps4gCJeKFs7gnWsX4HrXAyxJyY
2FzuVtku2gtMzmVbSUxlIMNfY8ytk/y7JlYgJKrGGCwcJVzQ873FPDjplguQRIte
6ky/OcNdL1q7QLEflLcDdBtcrXpLapSxYzKMfYDB6SNka4gTxmHNSnw++mckmzQH
t5G+GHxn6e5hQMb1ApQN6vugt2XT6XetH8xBnIrOePGgZRIciEDypzdUnzAz5KcK
9pvMAcTZa0IoQmqcIeH/sOrRTDQrTKSx1vf2TJpjX+Nt85ZeZBxyEE5LaJD/kyWL
ywG39higA4fztPuhdF/qYY3DWSNV2lIKEgLW6RXPSBg3LxpzzBzJk92R6L1fHiz9
Lt2P9VfsXSl+5YVAZ0WYeiw/T0HYANlq8hhBcrnXIHDGoZQnn4ghC3/wbFbLi3h0
JyYoZyZyY8ZIxvHJT8bw3rYN4/HWRUfxB+/QBgt8NZP5f1g14n353oM4OJylW0LQ
ejat/0u23B2ELyKnZdusky6+MyY82eiBa6T2gG6IzgqxGSul7RN9EMuVw2ZeyuIP
8UhI2Fb0B12EUEbp2Jw4Op2qP4oAwD2A/Jvv2B7tBPXgSCTJ6x+PKCwWb3EBqeLS
eLBGR6jSfze/Yp3DHrtjcnDVTEngHkBovS3lTJhuMaUKkdETxCkM+f7AaW1ZtE5F
4XgsKYQvfiTJakkRg4o0j/H1/s/DoCBEKR2W8WqxArQsMzD0nuKPtwgMvmVwYJwW
89ST/PQWlO4A2PfD++D9TfkiT1pMZrmvz+tldY6oRNlBPH3BI95wV6FpPdv9WG1Z
DhLX3fhoawZ+BZaufOVRftvgCSpsxnnlayA/nPeJIlEVPkX/xb+7gisqB/X4kbVV
Wli9pdDCia8wYNns2/aCP3B/4r2gFEqSfpmQpDnhhY7RPiYletosAELu6AeFQeB7
GAR6GicmBpLQaR6hUyXrCU+6HEEejdDx7nKpVpPJ7wiClmH3fyI3z9217k5NvGK5
+Ph7stNhj7CQcYEXN/3hhadh9tbCW9kDtpl0U3UfDl0HcOlemVKgYv1KuvinfsQD
FB8Yey8SVJPAWh/oGX2EU3tC2pjKmCFsNZ3fklkULwo838YRmFktpiywGcD7wLPB
43+2jKbn76JMyg5Y2+VZxzMjLUUkgtzam6eWu6N3y2NWBg+mVTx/vDu6TmxOQcYM
SUrAEkk17o2ROKe07Tqfd80A4otlR6J5x2pUL1jQboRMi6MkhzSBlHnKl7J1wLtP
Ahi4dMtfYwTOaAMIxytr7Gs94jj2aIE61a/M1t+ra6YVB6HA4D4cHCs8ujMimAJ/
FULsfM6e+qr5gWOKlnAcKeco1J1lzG6+Pz+c6oXXpJldwkrAdqWT3XoySEH79XjT
iQplsCiGm5LeQRGXYfAm5dQiZqcz4+8V1XxGyEHz3aMA02xSXss6Sysz7nSEZ4IJ
yw4rTOMdsQNyG3nICKoF5/BaiKkzj7aSKBOZ4AsfCeOLoPf/Yagp8Sb77ngR0SjI
EN7cxYTthDqkw6L56MeIMDtCwzJxsvTFj4WYIQD0TBX/2roM71cIKStzXB9NF4wc
fiLeAp7OQhMFuypaXCLmIqVUcfEF7V8NaaZF/1oRJeSlYtvMeLS15e4i9TYfCtdB
yqzXoMNiAV0RW7FDIsgl7S+GtgrjHyE+HlFhi2kNPvxhv4OUp56kZNFu1vtI5ZMJ
bg3dGk2F/O9YAGCaNAJV4KikzDMSap2ELFlFadxg2V5QYQRq/kDlIRrzk2Yj9t2J
/Zqh8QRsxxYy5KYEf+esmVLFpfF7OTMX9c4vskVLxp3B4LVGE3wLbGDRu5gWvgOc
O7cUYdxJMizBLToQe2DUtAy9VCw8t/+pGCcoTs+f7PLEOCe/iON1rrF4KB+ZrreX
YYbGALAyGmRa7mIvYDoQHHyJSujc27RQ5EQYiLwi2k5w+dn5n3UShfipt5pxGEnp
4czoffUa4B5fiEzBHwb7+/H0m7ZV/qtMe7fIs5M1nKRegQTONBl7FP2/ANmoePN/
kXV9j4Qy/h3lqkrKRNLQhXgglWGswWms0WkiNJH5SJGg9LU6LVx9++HZOI4fSA/W
Sh1qiexlOl3l8NiidUSeQhvp9wkG8ZgmezyiLxJfuI4LzBNgE9IMEmiBa4i5lEFe
r4UcTYIMRxRIPsBrkXDFEVqr3yQRHbQHDgDStz7jFcNkEOoDf2quK/7HAmyQT/ts
+a8Z0znYUZIFlQKvOsaG+Dqc59Am0gbueM6xqwKfbHqaLlNP7UazPwJE7vgMQ7Tz
qLB81UVEhkMfTQAWIGL4N3KlXSlBbyBUvgVryBgdBGmuKyhvYpSAlg05SP+0MEal
fsO/ZqMGuwn3mauCfk5ma0SYUXui3W5WLaRYmD9JGXyb+iy6WVRvZUVnVyAhGAoR
ol8XVejxn3xnaa31UqB2ALFVfVKFO3GC3dDjKDKdD9KGIVgDC7A+T10VxIuE4kXb
ttnZ1KW/fSrhIrlc6nlODbcudPn47sY45MKLc0t32oUsdrYzfUMKc3PhsX3Ijjbi
ulXSqcQUl82R+R3omoVJ5yGzJSP4U+ejbCEoT5g2+oU8G2LiI7grF9vs47Xftq0J
YM87s2lrcFEQshqV1zv79RHxompYfpWNQu6HFWn6sMsfmZbqVen1vi8FamtemnO+
Enaq7dk8gyb3z5nIXGRgVwkFCP4GNph1jf5oz3o+Y6/9VV3n+AMlQXqt8gVQNwl4
P+iwkFf/YjA6bCc+z72/a7bfwIDsFkyorQlQ9GQANOAI1b+zvl+Nr16hT2P3zE6D
Py61ozx5EfJPxGZo8A2phmerw0puLS9afPD6EVSk8badOumldu5fcyX1lBsr/a44
Nvqqs+xA03Vrno5Fi/RAQc49vZK/KB60FI1sdOiP5txMmzjfkTs2Do89sippfB/s
PlibUX9/BhwPM18NA/IhhNjShuJWEFGXUpy0pUQe3VewAXEXmUib/TUjAkIl5ap9
+e7CRXGqpWXbcSWzSyHz1af4hPQSQFPqASBr8MW8ZqhQ52ths6SpXHTis9QVLukZ
4yixVg1SG1IWxL6raHn8iwcUkQ4e50XTRzNrbvxejhxOlZ1jFpmMSXDGZCboSexV
kJSXep/dYN1lj6jFP/N5wVgw4Yc38yJIzUQ+uYrtACJ353krXGbZc+D9UgyZUS5C
3BeP3jNrBepveyHQg9SqKHTGuscsrowFmlr5jqIXaixbFCAgkD/NV5BqZNKkF780
v1P5s1RwRUP9CqF0+Vm0Qe0Wvh2j/Acrl05fmzT/K5g4RcyEhwyV4ehAzCmUed1T
bAh63K7xMZ8xq+fHCI+Ys2AB8K9XiZeR5VkdELNbeavfPYSDJBUxva8L9Duakxlg
jc+CisYu+460AtODGG4YdBc13juAYLQ37GEdG3cMvonojxwqo5qk2gCgmgvoVgAQ
NrNXXjnjE7qRSy7vJg5yP0CdUgMFei2LZsvMbk1oCVfqU48EF/pZOyG1Z7L7tnUZ
MSZfoUEsFPwJl9rstSNOZ3e2dc7K28bS5cvgeWFcCMAvEf076MXJh425NzjsICaW
0GC/veMyQkQ3Qrxey0hNpvdMxRE2y8er6ilJpHbw6lz2ksxTJ1E0w2iru54Iw+yJ
dfRdPS/LLiprjxihUT6fFy2qei4u4NwDOp/JUInleCKFmItcioi7q4PdgmVG75ij
NkzEhgQylreOUqt1R1vh6CcIH3bWYp+FS+D3Lee2v00819in84cO+CKoXnQNLlkb
BtMYUYZcLCm/6P0FGx1xQHAHxlYAKpcpT8cbXlfTdm6Pta6QNl0NuH8x+4qH9wI7
GDlD46zKPxsIYrKO5hm7JNKkX2lfMpD9Ewi8OTMjvK+A011FfFNsgkvJH0z1BzME
4OWRcgyCGT0R08ipgErb3XVLpijH22hJHmRidEcxH57nyNv9QSs5IPL3IkqOWBJh
6xpnd6Cc6AY0KtNxETekVp6Ud5aqXS9v/NZShNo/oqQvctzjdVSIOoWi/8p9q6vw
F1jPeB+232/IHrGmcuYK0vium6KZnvNVKyO3ebO4eFurDJt3pNn2zfO5xIKmmiFk
XPqZcf7KJ7CosBp0/glEZFYf+fJxk+F3Gr3M3vhnt7zDSRTYPI6LrbGKBa1gExp2
2MN2Z+fF+LIGqoU/4BoIiukfInUN8M9QYvROqK3miAdKQ44zrSvPfMD8RB8fJDvj
0m5N2vft74NLgGRpfj2IzKG29nKWsGFvQk5Qvv4kCBgbsrc+IU5YfHGhHPr/aXaS
kdBFA+hCp+f1GXmP/KJa/gq5HawMEMYiDkgPhEmq/rem7aGkWkTSP7rTdlVf7x/w
UV4+StNtoW76BtUyvpYHf/FPmJGDYBmCt5eqWqmroqHOivsFUYwKGUib9MiNRJ9n
XZFiwstBc1pBOX0clv6JeAHef4atQviJC6R8sE6QpybHXgSNELwiqlvsV+/dPIGh
62Zd11KjEII3HEDQ81EZODqxdNpT5XDtBaHqHotQK7bhcA2BYnLlNj99kgF0A58j
tFNx8gn+z4FLKnBwgEtpkjJVthO8QpyP19tNdNJcS/1viz/H/MSwFcbA0+LPMNX0
1ZFYV1ZIa+C8mwcqh5EgJ4p3b5565Uan3nYAFCDt3GeZcs6AfgdjgkeRXan2KoBk
xpbvORWd5P9q5PlDUB+L40kZ1qqFcaQ9yg9WEqcCWX9iereVhWjKeLWcXWbGXp7R
ti5zu6DyKC75WvLj7TdmeYIzWDsTw/mU80lbFXoz1nqmFz/8SOo5bB648xQQOUFJ
0cetICiJMdop/jpoyWD2vCJaz3doF8nsrJAEsKi73luOhLdOzmRqxbykyWoQBNzE
NUUEEcN64HZzolRaR1xTPO9Q1wLNCBDFqh0yc8XNjriHw9iYHhiHCkq5GtvJhEDw
A0V31lwdmVnCl0LC8fo5Irlq+tsYANgUJHiC4ddIAv4HyysWCLL+456JceIdsNpV
/ooGSBb/i1kHhxWfcch23cR3FvmutMFOel7/HO2DoThAJga7/uuJg+fZlifCBslZ
YHwSu0/GLweLONWjwfHEhVwb72c+W6YrKyG9LBXDBeiLM2XamqlbpeDUTY5EBlXr
tIGt8HZljhz21cFaDvIkcn4sb4fiYdeUZiNe3TvrqnjChBcGiGg+LJ0l1yMsQPxx
c9Hy4wX3kim/sUt+Zc8/vOKqu9a1X3T7zpdZ4maUEvfOlpm0MzSQTauHCpT21sOS
FIjJPhytCNlKk2FlUpKj976+fapiCT3jsQWjsFXz2v5NvyBiEe4SVBJI6ajQwN+r
Njx+vPX7wmiFw2+Yusd8xy7L4vl17zqhfvf4O6M3wctUiNRTfg1aITWsycgMmzQv
vovqU+yX2e/aXRTpaoBauMMhtBrrvzKZXNBhsxg4K1hL0ePmaWV+jqlV5Lv4IcCu
DiRjab/SKBdJwDihh9gq5Vpz5qSK17MqEpg5WJeNLjnvJyJbnt15camFtrBfb8vn
rbdbDfaXxH8QKltiEegNPuPhL8G046rtdCpqwBGaJGI4p4auNaEywQJWFacjTpEy
D7H5CfOLxLoRt8GMK6awiaKZE4bs/mOW75MStZ31d2P4kU4+3cOO0DyteqMqgG1p
iB9NkYRFqLS/wNZTbpmrfAOR3yM3t+4SKy8kAhywsjNtofH8XoC9b43+6+CQHjFo
gL6/k6eHrp7AiOfQAFZKbpEfMK9LCQ6CfKksyUauhziGITqm+EHPwRoqZOJaGAY/
Yw4gmpbUMCens7m2l4nuFBBbQAPUah1Mar0xSC1Uzzj1UoWeaX48LXFqPWMpUrby
s4DLIwUWa/QYJi6R1ay1XYfdSbgYUZRqtlHzCod0OF44s88sSTLz++mpA7+fP0d7
IWjrDkSWsHdylTI8p+gmspvqb4HUOgeAaJdVF009dEu0z0f3By9DyoD+ScCKhxqy
hN8909h8LrjZ0xmsgz3VT7iSks58rd2tjhK9xDl24U9CW5tENGw+If4c/uTvej/I
gorTQfSqGs0FeP0KAhmUJcn1VB/Ao4wVHTkVRfXWKnOjlrxD/uCt/BXYXBiY5KCf
jDgXEmLmtiYkbutFUWocTnbLKfS4tMDlVNZVo7+On2Lr7ROadmurehMJmhrr6NVJ
uqoxdTUbUBZMyFapf2jR4tdLkMjetwBkCU0pwfytWjFkHdp5FKdBqqi+4p/nhb1Z
621tRA73loJtoBPRCyuBGV905l0BJhMVxsLr1HymliH6ah84bY5FANZEMvOwctRl
yX5mjlru3dGtKQ5mJXmkChN7bBvPxT4yocvMyo1gjnivp8qdRmCkWMxpDG0k/qjd
1mowtMAaoBopm2af/Dxo/Z6JMMFtBsOblH22RigYuVNvQkyIrrrmuskrfxECUKJP
CRD/OCBiTGmgizEuQuYqbmcHbhuXc8hvUa0v2r+G115rsWl+Z0BBa6QCPSR6ETGK
A7CEa4i1KHgENXiGAmmCQV53LNKcTIZr/tNPYdhxep3PQ6MgdqT4nQg7b3b7ESbe
e//TYqEINCsebIpigoDzRuhkMucQN7mrRzCT7q6kKBLIZdq6+r8bNAgRD2OIKdBH
6Ag6Z38swVtsJAuerlPgPjmj3mlaFU8IV5ZzUpgKIKRSscg9owxN0W/X8805pna6
RzpH0er+b/udkSZFasKrDnfm0sxIyy73PFwBdHTsScxgibjSJfqpeiBsKP9u8MeM
6M3802TqyVBUUwmQi2wNmxk/DjTKhWwzF2qqTnvqu85tv0G91dk33cqcQW6PaYV2
nTkkbB0FsWwGmmpy4dzey/g0gIZ5nlABMRaw6h3DHZqN9ktQEZy5GQovfjZME+0S
IOBvw4PjazNuuA208aEckGlJBasXmQ5HtvqHV72iQz90DPxhX71Yav6VArauoqJV
4E0vHKPCcO56NnktS2urdZd52AxGkRDJQTRZKeUafuebXfmFTnz5UHS9ggG5yirB
euGApCmtOGouq6lAyiPI5OGfUkbyie4R0tlUDdyDE9WzAhwWYCNtHKn/Xi5e9nor
34e+WqEqBB+jhvuijjgAaADNVZo6JFuLJw7la1kfB2R0m+/Ea+gt2spZ0Zb6QIu3
G+ZIdpNe6tYCOr8Jjv9PTyO79mDAnbFCpbiBdhV3diadPCJQKqRlaWsATuQcWBdF
fpaReaUyrPRkHOTEZb6lK51MXQDNnZCltGQaGuB9jcG8Vp2kUV2WR6lOIyjKniK8
c6c0Wmk43a12yhxSIafCDN3BHa6uuDtTh2iFqcKq7WGbAMZGMw075ibPj8WTBZmq
LiKq8T4roGmjrJ/DzhjYIDjlr0/moE9fDvuO8CLeKu3z6plT0DGc856S4w4wmbfH
7MdhtRSWZndvpJwxCaD5w1tkbOyM8b6ngpa01+uJtnRqf1YmjbKettDtaBtFAmzb
R59WxhajiavJqnRbi5RFzpnXdeOmUPxQeyFZPnVACbKXWaSVpJyvjEQdRWWhq4lP
/MzjJAFRdBLnA6NyBkKrjUOICLxEMLo5By/TsBLe9FBDP3QaemEdxLxSEcC6fZk/
wizGJbFtL2+Y5KM8eDMKc+Q1kvR8zP/EmeSD2DvAoALqqN/EfbIV1YfA6eRLFC9c
BT811/yqxV1hjb3oR7yMdh+jOQPFSMfziFY5ytgjcIcBiSNhrrZYsq85U67onPwt
3tunOtSyk8q4RA8qa82/JKGJrs+yVJykIDngIs5Yd/Btch1YDZcs+UB49p4xGYiG
LultKMD/1YvX1Q4EnorRyoHdzDIlZ0pIDZJ4hG7lGPktmXbydLlbKhjcNjHfOlYU
HkCxG2A6yypZW/GUm8cUv6mO9fHN6oU01OT4yBbFarErfvfek7Pec7ru79oFWYz7
gQrG6wOI2oib8pKJqrSj2FB/EWx5r61h5os0dplRqUAS0GqKI9boeV1Yq5etMl1Z
IU4gUcEv3bTO/7VzyZ6EIYji59zN48K13ePKDdPyaKmPlK2I0laoTXyRSu/vOz9m
kzel4NKPyFGSjg9OcjXcd+9fUU7Hb/A2gafE9foxODx1CfskYuh0M0NBjY5hHzeH
0k6+ExfHcMCxb9nfPxh6HJ+cQcPl4AC4idbEDUXlxQadwayKdfRK6LXLcxOR/NnE
of1fyw852h9PytXRn6tSFe8rzGGV9rHytxvWHV1ezZKQ4JMl8V29UEcuU88wN52G
KmuvN1GBR8irGmaV3hRBbBqhQPwBDGAsH7hvbW4CXI5woiGuUqR2xnCLXZElvXof
3zC8Q+H/2j6LPFyyKK+s5yUODDdWkyhTnOkFQEMwSXd1Q4lf5Qs6RFqNTcOZ58s3
NoCxCNM1hIJSKhPu8i7PQpCCCCCLq+pipZUhV84qT6aFKOd35qLqtHncYjgV0qAX
qrgGmZleITAsWnwKMSYMCH1kTTIaQbFhMpFZ9APC00IdOVRw6lHwKDVqDR608g3v
C6bEmQIwReI9R4B84t/fa7WLAMPnTWSPE+K4GPuETnDxoK9qKr4qWpvB0stFiBCS
GmmW5Dx8+mYq2IgXQj2xl8uPX+pf+ovwrPLaJ9vaGa8YldeoGSs0N234U7zdlzKD
9Ev5HoPyuNmZR0hfusAgpTS7kVslGa+9PoDO7DZUHQXxJWaxhv0esmB0UXs+G9+w
zY/y5csK4VgEDGsNDDQHkcu05PHFvce3w4zZSMCqVTNlNj2MtzKEC77rmraumMzP
wvcuYPPFPYDigCQjwgcBO3i2fAohpfQDovW+pNSiKD/tFhQfKUc9RU41ojnIZXF5
ImF7nuJGaHmK6Uzz285JAUjWQUISjEdvtYGjG/dmyy5H006uca14oCNWfopSGGJP
wYNE+xhZb2khrYGLJTA1efdxJYJFPjeWersmctOV/pP+oNikWDCzpQa98F8Ws6k/
cq6ETVxdKT6I0qmZ8mQe7TSqBzI0rS9sjh/cufJOmvwpICkMG8oqGxCWi7IIgKKM
XZEPYJ2XNHKk5T6LJejvKiziHu3nXiZ+3jZB78iDJT31qt20SlPpsj30slhCQYGO
QYu3XeJH4SG/NBlUIBSVWjkDWvjQbyHI+ubwCdPdoJs6tN79GxZnxOBs5xgRb+MX
FoOXZx07jQ1fAZGptDXb7yXRz1ngcnLOe8k/0jgB0AXKP3x0Ga+KOj/7FmxpNBQA
vi5oiDbI55asQd1kC5Z5VdbyTFUrll55Q8dG2pX/YOnakwxbRlsaLvp1CvlLYulp
BPWghvadN9YoPe+KXdTqGJdsDA4JoCB00JWoXL57acpT5HcWJ/ixTjO95llbqvp8
ZJ5883QUdskxXGOnG5r2R/PLB/HD+Mi+gNkPFnVxhph8rf5oOfqw193wwIEt8f4V
TGyvTjLq+mLxsmpDOaEKHso9wCaA78tQtDqgUu7HFPAx62JllbU+RFqZ+N9Uj/AY
GBLeciC0Wko5iKOEIAI6sdG5rugBm3bOj4BCRaWcLOioQUPpgrhDgdbigq6X7e/S
duc+P3OorNrAIhH1dFof3m6tvuFrUhsQPaSfv+DPxCCmtYtFbjZmGgtW8pGlZ2uw
4ExLDuz+HpUNXpj5ZX8rseWdnDpKx5McRG4TggG9j0XungyMtrs1j8ZpTLhRxlsT
e0oTtoTlOT+VOTDVPGSrog3hwLP3z6viQ3F1jJIGFe/VS0N8nIKipXWksG0Z53a5
OLNy/oKP8WKPvjoxjuQGPCHkaVy7TZc7vqkccpVP9I6vrGMTihnk3tuVXijlKHL6
ONh1kvEzaZXR6KN8WaH3DTIVRlnz+dC7WxgRYZruXr2lEuZnD+VmStM2ONs6CSwt
fYEPLvsFKsOK5DbF8zFhgvEnnJ1JZn+t0hX1JGFCmbBsD5Zq96A73r3Nx0vIIWU5
6Ce+I3ylLtgrcJFR7HOw2fpwkOUwFCDFzi+IAwQUbq57gc1b3MTFf1nnnazDZKhu
Rn+cMm0e1KjasTRPY2HtZKHSZfwMBjsVjuiNCabnaNe0ZQ4OMw20dvJrqHeb/PvD
sLEF0iSRzxG/choWTlW0n8nWAwy4VFdLb+uLU94V1LABYCGHLNKpBWNujQnb3zOX
Vn/duGK/TLyxXV6gEOCpQY/D1WkZJbgkZGrbURW84hoebUkNQS+Nh+BSsqHj4dal
k+1fLQ2SLziEu+DZ9jduZlcFzwuS8mZ50w+mUGNCNQPLK2Ea8kNzKdSr+eLRcJ+H
nmZArtmTF71cnnUQ4KZVZYVEgm4KyZapfvyjOCMYtRJtTsAKV/evs27a1Y+B07h2
BBB8sNynaK2sOVBCwQMgncl/nb4tZLMjaJJclJfB9QTObzgy4VBeSFlQw+/EfJBI
W0KX9aN4CTV4uIOFDhKiNByu1ICWvSCEo6CBz2Ai6qIBY8HVBbBzcoIzeZC0Ctxl
nh8LK/I0I/cgzP6NrNNrRJ27w8ggD8HSPRNcy/9pgMX33tULicoeS9pBtdiGsugB
HgBrBY41LGMR2GHF3nXK8q3WT7Hlf1VpozUg95X4Yh2bmBz8WeAHNYN7MhFcXxee
bD4FEg7d1iSL7U4BpKpjeg3POTF9RZWkUtA4bsJe9NJI6tW/X4Ll61djmHDZqL4L
wr2flwF35kOUA3RUYH+UYWODrwTAjEPzqZ2O1zhVjHPSicdDDcv9ck2FOZ/e3apv
WIwc3gKg+G+dN8hIXnNK6mz2WX275D5dlb3ZEKxlLtRRlErd5+6KgaLL/I802xaG
uhYtH5R5rJHQEOWtnYVNkH3mZdOaQeLOp6kUv461vFx0DLhtZJKsLrI5rBQnM8wj
J2AGGsJ9n1gjxfGQMShBSAW3d68Cdbhb4MxQeX2xV5I/byHshy0a4Bpd7h+KSSax
poOKADG5suENS+bdhCkmbcfXvqvh4ZMEZXgCnJGaWwsUwwJYUvjxbEMqdmHn03/B
tz0ZsVgNa/Tzy6pKDzPXtMBH2uzCnuk84R3jF6X8oHwMSh3t+eW4sgZxio0QM40e
P9ORCyOg7lZdxYGX+5dAd5ZMSihqy6NHdWGjwGMk/So2EzraUXMP4dnYQLOD29uk
QTu0B6HcGqDcKSA9gvCvfiVV731PfdXqvu5RJDCcSkLjGnEGe0rcSlbliUKoy8G7
ZkEmpkuzMV28uAWbLnNmH8PSUXZb4E5uCUXpUrtyJXRRSjDtjVscKlp7y0Yf5KXs
pR0QE7UX9CBoX0nRKafBz9W2H4/Hl5MINCUUyfm6oTgvRNvGe8X2s7vxQM/Z+9RP
VL5KmzaynRV6IQUWi93UxtTOIfT3xzuA256C0VP1FjFavcgS1ZAwRCTVSHsS1rYi
CyPc2F+FIJJW4OBVuIvCiBfx/4OJ4vYba5rFEExK4meuK1KVuCvURAPa7c3H7yP0
cpJdibmRccfVHJBhumDzZp5QxkQ2rsvSFvKXL3rp2VXawMDGlelKuM4hCRXkj+uh
apn6k6BR5EODavbnwGZmMIZiotwW4g8NXZKeV14iHOoYJ81kiJnh/94Dkmtcguim
eOi9fnjRJbWFHOIfGhbtuSOJVt0pvJnkbZZE7KPkFxBpmttLKuuzZvWL5NaGhvKD
020LGq2P8g4PPkPvh2CX5N0jUIJPFahTwp3f+aZgCIccCI4OJOjEsTgOVV9YUPOv
P3+Dza91b+WpIdOAUO4jbFvyqOBaKeDJyNDRwIcrzG0hVFmlvSHz97+TpaUeO3qy
i4Z/HTZI5o0LDLWjATdbgYUpnneuP8spnoauKOKGtygiRYALCa6F4C+fuE9gV0Tu
/jxhBI72xQPF2bqprdPLdlDVIUjwdTA5GhqQjVPFyz1aDt+fEf1ely9FbHRSNqBx
zpW30VoK2i8CXF4EfXybpe0UTPR/ZbmTXiBbiagk2D42BscU71Z6XAUcgYFkwV1/
w2Puofwql6z0OEQecSJYrEdL6SABmsKDZDdz7KvJ39m768tgC+zXV5hv7KbqdwS0
cb02aC4rdjyLCFWFzYC+DJbsogX0c8W4+EeAjH6KZxP3OmD9QLq/Pgkcwi5YI120
hgNop+TNogF3k0DUC4Kd2EvmKB4M93mjvBmXR9beZnNyooRvXgAK9bNLyVFMaznJ
ouXusdGtOYIYQaVZox8lQ2cCTA+i/5T45JYUOBeraLmyCBPTS65hNwElX08787IK
kDrAMKPI/sUPM+dWGMv1fJ4iQ4mY9N8AQqTWGjdAC32ebFvWUQsOCLmygP6TRntN
27FpGSqYt1pe00PXw7ey1m9CpDyPDJPyerLfvK/w+JbtAesPojmP+VcRE+owHUeU
gdYPUpZy6kxZIJE852YKY59Tx8Klwl6N6NR1Bu8cUo5FIWwXa1XlZvIH1V4aD5qS
POewqCg9IlbcTx/cb2qujFVomupsB9cuz279xKpp4S0OvGK8jrSHui8jrTK1OJ4m
M5u2k0jqa5nSrkj7aWf5c24lA2n1U66sQXoR3Mv8M3DIYIgD8ZoShmljGdZTMNzJ
X9fawiS4kuoB4vuc6YyCtC+IkzczwjWwMrkmRKzHl0sxuIxnStaBC/1d6BxTahzm
cUhlu7UofZ+K7A84jRetjqUH1A5ChCr8TWPLTyKKWATBF4g7RHzqs2z02u944Pif
ya8a0FFpUgQpm0vCU8cWsoUS+zfy61YDoBIoVqcGEYZdjMAevFabNZiZoN4f6kvp
58HFBIP5YMhRB/hX9vRA02oRWmXd8c4egF4txU0pVn8vngPo76RWx5TcJX9luHFP
4DJyNEC5Evm/X2XvsO95MsFgX6xIWxivYLsgkUf38zYtWzwumCrQBuX1cbcM8ihe
k4M7mKt6GNwqMnTzM1VmiJK2pkEwNKlm7D3mubxIZIBIADiSp50If+SJMMWlgJQ5
cmknHL08qCD4PC6fTPvdcyOMIsOTvVXYbDE1WRundEjMJdSn1RdjwuAfkaRG9rCH
t62yszRmIQljWm+ItytMIyTE+1M5beLGFMpJGm6eYeeyjSRhSSaEpSnZogUDhPkJ
NsMEDW1kkL6RZadZcdUfOGbweYyKlaluwqbbkOaFzNFLZ8L/j6lVit5+QBi4NiQf
L6T0RTIe+rwN1WzVvAlHdgiT9jXogvy4BR8MEtTK7TqmiVsC7AOBzuF+IcaE6+4c
9g/IekV7cCm/irNZQuvGl4BMFzM5HoFw+MT7RhAE6GG5ylHgpjBF1QefAphjYaNu
G3pJzoW7z7lVy3bHzxxZWr1Ym7Ygwq5Wqo50yvtV3lt1DVXy7dc5cYe2eyGBRqA+
/hBmzl5U7WQtSQW55lRpomyhrTY2Zf4MWO7QawheALA3KhOOPWR3y9jcu1vGX9lB
HCkHTqvIar9NzU9vl8+FAcScNvbhyB2wsiQhgVsnwMRgaHmrOJBu3zFx8kpvVBWm
thygWkeKyLDWu77bnQS9aikC9Ww+Lv2ZXKvARqmlJzu0rMPFXVqAwBlNsTGAIYrt
IvrXPKJ0gp35gkIAICfzLTp4pseKdVyzFjdW50UWtmQg1rqzcOyyT7M9gL4cgjmv
8hi6Bnomq6uG/v8sCPWkxJ9XVZYEgxEGwkI7rHMo2a/wPm8ef4/ApBEzgyM62iuy
UukDSwVCdIs4ySSRgEADFdx+sc45OyJiOwCP2smpw6AOE1W5WKybIyzNZqxxIz0l
I9MyaPIEnwRdhK1iCs8eObkAQppupJJ3IuGR5TpjPdQadfmftof+P/T+UWMDQ862
Y7QTb1zdHhWv/qm5FQaIBgzybkAx61/EvlSgB/eCToLXUdifnwxiW6R9C29WeMox
o8LvwtUouGjK+veB3nVY0ZUjjSHeI+8fw2DfL1w2yEuA+mymziO8cvmDt/8jvHQD
FXS+LCRxj/E49xO3qIw77AZ3vTXsy6EXiPsWkKY/Hp8TiVqmdJrZtVZAm1VNsQN5
Uph6UCSRNnMB4VtXWEfptfRfHxHFVkMQlWmSFdOoJn1tQdeFRo8q9rK0RZXox68M
bjLL7MhoAAejtZOXIXH2632xwIHIGwFactrXN4DBXOlQlLhv/H+qej+/gryCjYSt
lO6mWP7eATpz5pWdYeRQKQjD83hbyVVvS95WpnlDSdf2z93fBndzMTMUNXF3Lh6n
cGVRL/pDpd69GBY1mst+zfijScN5+7DhkWmIpJDyyR/5Orj0p0hxocbWvTb1mQll
/Rbe6MUDwIWsS3inE6oNd4BKvxKfpmF3/mp7ixm86LiJ/EouU1k+P8vfZ1yxlU9u
KUXfH2QvVMtbQCV3Qn8iFwkJlWGj/9zT41FEI+N9wX+Ev1pE3nXmcl+46WJMoXpO
62HD9fFnSB9xj9SpxfckRXkX6v9FrThOtl4zByj23vVhNs4SmNVeybVnL3Lr8cW/
gBR8dfYAJoGvPRfofK3AoXKrTJGKAtRflsagyOJHhMwZP3WUbS/pXRkKkFuIXR5Q
Bayf2X/wC6yeAYeBHsD/ZtgcLTx+v4Pu97N60skSI32SESV4uGTi+fXkOyeFjC6d
0c5zy6xd1N56kTX1mvBKl5MyY5JwgoVRPvwLnWMDq2opgKamD3GWnsrf0Q00cS8Z
3bX/iPGZIRi/CPYeYTHIpYWZ4gI124MlSC1nZ3pBv+P7srn8w54XE70i0Dn7Ji40
PK+y2ts8AyJegxxouNZx4uzvw/3rwd4pz5Ex6LnSv3tCbAMasj6jUNgtZq+FrArP
DyuCaXtIQekQq+GfQB697BnJ0ufiQLma63QEgEO2P0b26D/vcYKGyckPmyeU/aG3
Eqzyo7aG7t0X3/m+D6U8MxHJWCpj7Ypzt/hiGL4Hk1cUfvY/anjjeMQnZknVtASU
cGlLxLbSeVyjuLUU2BYp5QN7WGw1wBVBRbes6roGSWwzJFGx346McKzGfs0Wg/yU
0/DFN5Kpduj5x3oS8+zfDA7Xu4Q0Eoqb1fHEn0FLe3bcg42Pu7GG5hXPIrT7FBJk
rml9ttWWXBfr63rfiprqvEv6IPxsYuwORS9AAOhorpCBF1hQYq0tDPoEGuezccQ+
VO8uSGQPAGnWpuVVpFffOXlUljEDShA+qlgCrIINo4S/sd5nPI2oinvC04PIw/O/
kwiIDFPgk30vm7whpQ/SNSfwcjqW5B4YA4f7EfpeydT3u1ZIFU/DFch9uYHZEt3J
AyHh3MyJcmjT2kQMGJ2bzok8DrVTTbhEjsu4Bz8uTHsN/lkSZAQ2xO4Khi8BXH/U
gCBCsRf6IMuJ97cyVeL6EsGViT3sU0uuNrlvTNaBjc6oJxtHkli3Xbhye08V66fD
i/HeQ9aCtk29D7ouOSaixG5cQ/WeeUcl5W6+HkhcaO120nBQjzjQTxdb/52GX0y3
ZXiTmfMhvr9WBMENcHvvc36PdXO4Q78EAm+AUmqJOWfiOI0BQVaiHnBnIKmb0III
Vw/my1QeOsrX1JP3r7oxddI/bPIrSu7hzOverGC8NIuCURNJyuHsGoGK6wTSe9RX
MuZRcxSUJZjJUvmNDJq6WN7ABMPCZig6ztTLtmyKub+Qf0YEz5ClEiSfFIX1G3oP
2Xj12ntriBgw5pJdwH5dTgdEenSLffTNqnY3yxeAq3n6XXxTb36V1Yfj/sVFASnA
n2dknWS9TJ6IqELgXdXlIU3F0yCNFxAKZV5ifWoxPsD8BUEUB9sv6/MDopxL+95U
ZJfzPrw6ibGS7sglFV9mpnrm2HOpH1MB3QvEOqpy72dNWpmpTkfy0Q2IzaXOr+Ke
6sTOWNX3hrsHWfUtVNDl9awdpB7gHLIXDL5Cu1dQnkt6suqiqz9bbSp1YlphxXj7
tb+MQUGGEx6MGXK/T8UJVJK0pTF2QcRIYXQXtCV8ZgTfiG/luthw9lYw4pDgywwg
z2Na4Be9wiDi1uF/cYj9/Slc7vKYFHwFS6Q62YzXT87KuBGTsORYjGN0vGhK0Pjo
FxWsLkTTzzsltNdxzdbLqGr2TFY+52d4n6iaxGq9rsTM5nxHYS+grCNNOyDpV3G1
M624dqNLhlHXP6ZGWhQd9voXGD8aoywUCoOObF0iv/9e7r2TX9rYiltNJmF4MUAA
YPfWLIgl6E3e6sxAEujHEfkSrFFD88WvrP1gbCl2/sIho3TwHnln5uKVJntZ9QQF
IpdG8cuz4g4yXofxkc64pYLERDC3QNcTozV1cpXymHdRghKYROuESa0MnsiNnQ4r
iRi7WNuSrXfH/FJX9FLWTdkckPC0fuBgcnut9eB7nZ0m9s4zx4WX/cObF4O23NjX
57UsFGYLalU6OkVoshY+VjdF531Wx+VzDfyAeaMiakf4wpkrXB0Z9/rFbn1fJ3Dx
nfivEobrKka6cxx2VWll0CbhwOcLai5C+0DzahhqQz2EXxTAP1MWHttBQ+dT1tWO
E9UCPFxoKRv8ejOF6CeO780X84+4uvpHe+ZrTDRiJzuTyEpeo+XV1VLhPAWREmG/
b65V0cbdPEA2nmOWCjNF3+n89ozsrzL5+/gx/1RBYn9cBankPLQmFSjiFz0XSfAy
V1XADYr35XPGe46gR5YZAS2xSNh0JQwjjh0hygG7Y+l4m86LYgE7sBdZpS9qHeAA
f9GfomSi4f32rAU9uCX+dCSfBMs79WdUkLP6ne9uBnlHOTtklSPYeXmH5YDDF9S0
XF/8GGvoaf3yHKuOe4jF7z5N1M/ef+4wjnbstjqfA2Zgz3Zz03vXKuAfYCyBF1NJ
nazCxfq7t9IHRIVpAUXzxzDNy90ErwzYa9Dupie6UGktEd0JUOvcEexSvWWMbFlA
S0HUhWtSa+PoBh3L+XdedJ4CkgEvf1z0V9nB83HLpIHkuB/jdKLpNZwS4Wfh71ur
bWRe7E4DTNVP0O2zGnjaYLSniyf7kmUXjBPiqbP5TbYe+6FLf0J6fDM4+lJo2YEb
a/5aNvpUJBXfanXFChPHw5BhVVfL9PrrmXOM1Xllc0tAVnwNspKALQNZZcIFA75U
ZAckR4sgj97BkrFQe6NUk2BBJI/oPxcFQJfTdlv8b2w/pLJrwbP2YIl7sfddT2bM
ITIIHydx1d9QhCohwoeVvzD+W+iXqag9cBcIHiHG9dKYpEVL87hVDJIUMxv81VvL
iAMZa0d6xLcNPP8j0GhTe6wryfhlxa9P1x/XHvy4o7OyMcW7QOsA4pM1uynIH4Ty
ou0Sic1q5f1NfFAjrC5y9MBeX5acT1YoHs9gch5hT+DwxufaRL1YJnspcrnLCNO3
dfgiFqnGXh8ImOtmK8jgwE11EPoKxcyn6wxv8PsG+ZmzvfvZK6OaUPahGHCWE6gf
Q5nWmBlXSi3ZBbI8t/LvJy/Q6hTMURppEVLuG5X29Rh9A/fmMdsjiRHf1KwI99ii
hPmwsifV7bemDIgSkLfWFxgq9hsoMJGw05iWDwatqaZclAI+Nt4L9bFi+E61brUw
IrOT6LtCYYNs/pnpyTziwrv5dUJ9zdUhBQlILmfP8jqt/aaDUT3Qu3LujXBz+mJ1
uyMIkJpOwvGLdSeTnEia3bjK0CpS07TXVLCHUIrviwpg24aTgfdxariA6JRSN6UF
XjpdrO1rzwrkBEwTIS88Q+jodWX1oNm+h+ouvGVnfVydO1NJufWiLiD2s1IdyWSB
CslSu2FfGE5p8s6E3tkf5DCyY7rWKHOndQch8o0MyRNXdglAMyL1+0ljqWy5t55e
tKep96iCcmFJKonyaTZmyh4joZ8jGL2aJVZo3W4HZEdPGUWVt9jilelUWLkJvGWw
GlBhqFammBLNNq5RLnihvwW1nswpyhU2G99RpkDcaQ0ZvRWEDJbYxFrx3bVpbrkF
hDzYS1/ntZ8IqrqKvQAjBZoo/ookdTi5k+yPyllJUP5GatvbplBmrfOQxxgwqj08
CwZ87vE9O8pVWw4LGDJ8SlVHChh+Had5sfMjOVuUVec4jJRUmofjZuc7XUpGw/si
ZcZ25CUH1ete80E1ikxTLQvWO3iBIFdY7chlDnLV2oiXTml3I8cvSgHUrV+c4yQM
gZceowPJr9Ne2yAeGvPXtB9lUWHB+AxDKswU6sm6oNpg79J7Mf+MxzOoxVvCo8bN
3hqEUbDcvYRd8+igfRsRXTmgkIAdr0EIm9oFIOoRAjLW6FcstRHdL3dnh0VrDns7
supc76fXe+s4A6cxH1gcqSsbkbMo0i0ec2pJRYDAaN2OdFMW1gLvmLgfTsp/A7zI
6GairekPERD5znOsNifSBSKN0c6yzDikaHZqL2noxPVeIuPXqhWyGrmslr6Xe9sg
oVZY/UxquPXrX/sHXXBFJGdbE4Nt+MAhJIHPglcw1LZ9tvmzhewHQvbJI2Ln+CWD
9+o2wjS9wZLkESgjSwdSpE/4wcUmWJza0orC0aUJ2xdtgAQ8K2WEHmYnkDn2KgOQ
uZ5jYENUiss1ZXaeIgHLBdrmP2GYRXqm5ptCdOqI56Plf40RGGwfuHxqqVg0VChr
ttGo8CtLpl4n/fyOHw63CYy0HlXftwdqqoMXXiwOLGwqzqENbUIAESTPDPyphqW9
o4HW1IGttc/swAxs2s9vcPFjairs0U6mcoLh03sYeR4vu90j8Me0R5G4B/Vry0z3
ZFPcIv4OW5OUlwQDVRTugf+0IQxSGYPkk5xdeIUIbn9Qyx/U5r2+r0ctAjpvWxDY
PdftqrHqcmWlmVWLXTSiR6SSK2zxhFoo52X24D7OxtlNibPpdelpNZ2PzaBYb0EM
L4MeASBh350QVZRu673eO1iDov/8vFQ8bLnZnip9bq3Ny2Mu1HRFltC6gGuvYOCk
xJJO68urDv80dAPaZAkaiGMFwIm2B6I+bQdDWz898g9I6h0BPtu+1zbyOgS/ZBqz
Ik0utIBKKMUHwWkTpULBYPimyrngMzTLTkbi/DrPamVKxM+C75WVqA4gm6c6G7hR
b1y3numa+p30L9PJ3VIPT6pROmVcoEdlgIobuZvgG4duhSFd2GcodkGuRfXTQ5qJ
bGim29tgWxPp/eoxvGiX/cSHO+F8JgSwHQdNyv5qfvjyl//PNr6/nmdKk0mgQDE9
vt1N3BvVAhBY9Tdnm275j54UM8AMdL5R51EurAXmrjrRBnh0duhBOpMc0QgTiNz8
7rLws0LHI8yO7E7ATGD0DRODt07gESERAmshktwDZqDJp3/vfXXij6HTXOz7PVj6
GFHPRm4hjst2lednk8Lxl1RWLaEMcUZq9O9aTDL+PeIsvw5KW1hwA45JQHJf+3cR
FL8qMzddi6lFdIqHraQP7G0m18DRGQlXvGFGWpb4e5mKthtl1hc+10fJBAR6tR26
K5JEb43zvkYgea0YzeNdLbHgp9Uiy9bhhj5H3rCwolYl6n6X5R5N+gZjGybsPYMP
czDYr45tVVBm/QT6ljqaJpjHpbD1UAmCWi7lK7Qbae/xYaQKR2ukUXoGFSx10w7Q
PJYp0oBCSiX6hlMQVP0oKbWjt1moaSuDoTKoS3bpDhfdVBde6tT5epCc9TgXxEz9
55Kc+V4+qI/UM2V18p8buwP3miFUxZBwTtlpG/FumavMhs3sKdZyfCJyhlACXdbL
65zoqZGK6J9wK68Ws1xXItkuz6CB8AOeG5SOJ33tbLf9QQQS7yfmHFgzYQm6Y8iS
PqCEEMNWqpYTZ/RUm2zgchsIJnqsDX2scj5ipH4MoGTla6ZDy7ZIUx5wy7et/Jdq
GRvgz/3Bo29cL9td40BGCN9ENWPgehvyhbly+LcPFHltRHH0ZbkMAT1VnfPtMRcq
cHFS6kAuA7NRt/4nPo1Kx4ZCuPQv+ZLFt3pQyBw5UZRWY8inoxZ0rhIeaLD/l+4o
QjaJshGBkpecIzbOLMk7DyyZeH1yA1No/M1LSkBUFSaM/Gh5iyrGTRq7GtQIfsy4
Pf+JfCBrDrMyIgmCRem9mq0t1Fd15FJcvZgs6/gQB3W7gm/kFn1o0Gjo+fMsB2TI
oC9eBmvVSHAmoyCUTxILr4Ug++x+EatHm7+sbx7LCos1QpbHgCbLlIJDi3Kx4M8M
+s62Ooriuxi84q2f0FKnb6h2i3BApdjhVDKp9kSRScwjcZFnfG+bQlc89VBp5BAt
Cn0fenEWNNZEcU9cY/bcJ/syGSL+uJuAjQa5BV3/L0taM3EJlszSmZ6O//w/jOro
xjQuzEps7dYalLeo8U7EDEqYIqA/vgxS1Nq5YAcShmrQEqtDusluHdPvDN8ux1n7
IgE8bFblw9rnnR53k42XFsEc+X0wKyMM2tqVI3RupeO2pn2ulmb6zBc+CSjbobGl
0EDuJd3/Wa4C5Q2K/FlwCXg2iL/Al9VcdGrf2T7UVvweatWOqYOQ9A1SU0TpKEuc
N8jzq7Rpj75lcLoJAPtFRC3RhQP1FS4iDHdmtcoT/aCPYx9aQp7U9CeAHVI36MNq
6pchiyxJPgoy7WELNU9g6TbHVBmagrFl1lKCh044p7VPyuqq+yCqDvNWWsLXdNV/
TbBLyhF5fQ+EkGUKS6Lg5w85FibMTG+1d8XZ5ZyJBfZ0YAnZBgL/eV4kphFJW8yz
2WeA5lIsjOu77PNnlckiQoxyMm9os2OE5ZMvleQeMGKQYUdc/FYRoic4RM3wW1Gs
9DIVCGi33GtUbmQpSN9EiGoSYWUkok+rashreUkomUpMbqcD0Vlo0Dz82wChg4I8
Mj+LxGuX4hLJZdnijH8oGwOwog9gokEm/zqvocN9G87GAoypVcu5ptXyMrVoAOz8
fHDY3Ybao7/H9PGbD2zg82G1Xv0z8aVoYSSWkYTD48LV275uqquRfTZuMzd4UcPY
RtworC6bw/ayogqVbvdI5d21TA6JhSnGNepToIOmjqUVlZA5YDUfudbUJw5OwBRH
A5B5EW9rKuBtppVB2UESNy2XMCfoUWLjL7v3n6q/TqP9HFBZYFKJstfBA8tBHW4q
Fzcq8l9vn8YYlHDvJF8ELW6vQE7NOgqCluCIzoSUezElDXrV89U8m+UgvEh+nIjP
lDTaevHuUVQoGUnbrfVq0eml7KIKb1nDXkG1Dt1kSXXm43WU5YoJi7OYpqx0cc6P
dvkDrfLu9RMmX1AUECPAndqXYT6qWbFlmFwM2+7a4NwbNDFax8diowZHvs6FV1bi
RaRNzbqyqqjIiJdjOec/PqxabvHM2dbY20FEL9Vbd3zcaRxIicicWBGNrGkkNoUt
KGNtWkDp89Je4/n3Re6O9MTd3ecZmKg1NvIqsNkn9qfcqp0eUl8iIYAoB+49un6T
N5bvOlRx1GMinwyqWw884kbw0S8lHFG4GbOUDTfFxMcZ1TTYcJIrN6OCFjAmm2RG
ua4N1voC99dng0M2r9vP5CJS9eePhTpmWWp5clTu67097CVS5VYfP4i9nwpFNfiS
2PtlSlk525HvkgDEwYBC3QoDvEPmGHTy56b3lxDH515OjIJtkoMjAIgDIJVgfN6S
LDfiDVlvNI4v8IbLZbdRzuBpAW/+pMqtimTfeLeixLRYELELd4GYxy1FpJGyKPnH
o1kFs/cLPOKJlnBDpHkSmlbOwJMRrx3dQp5s6a3JSJZyIQ40rOxWuEeWHA9riq5w
Rgqv1cwvFLeTV3cNt0Gi7iiDrB2g9qRdai4Qkus1uItpnnhW5wa6/QvtuiPjglSy
FNLqdsDYWFMDxdq8WUzNtBgQCV3WzPDX0qBkSJ1fYmvkGIEvsHO/TSB5nOoKBSM6
k6gUnvfHniwLdLImXcIklSLS1y5RUnbVNpVgm6Cd5e4EO1cKu0Z9Hh+VfkeL+dkG
M9PQ6RfdGqVL/0etQb8McPP3LM+htG6HtFBURg/bMX5pYOngwHbzdbakmJSs3eMK
nbUH9HCVTpitZYkBj1xxcF7hnKRJV0aOw1gYoKOGE8x1IWS2Rr3eFX5cmm8z7NJR
bWQgA31P4mD8y1+bDzv/7CsneKWbjB7Gqr+pUPk/EuzEq6g8OdeuMu1fUDtjyCKy
SLd2RTrV4ozrpUnVfwhokseLaNL00fbMJl+ULs9mcZOIuuEk3uqzF7SI5m9VqK6/
arHt5G6ML7/t+IFM6uXGpTGBgVgtVxpctmzxn6tU41uItPDAQCaCNrLv66N8v3JA
tsfu6ouzHE4w5l8y6lX+wRSsp2pdsScrZwNTskqcOOc7ZARZmP8vGMRuTqDT/iDq
WbIXdRWqYAJM4UW6gqMAqJdW9l7vxWyI8EvaJh30j0ys+MgnbfY5XMdPfWL3Ht4l
vdrSZZS69rnHoRQEi/J1ZNPcWNTj2YnU0/9NMMwPcEgD70yCEAOgEOytGeupokhb
xtKqpgSw8QK0NALaKTpNb10yo3ax9+dCt050Yrk53igRpf4vZ5CcGZ4qGjdzKxJR
NI2KpaV4AwXKRc2DO16s0sji4Y60u87qBxXvvVadVZR8TSZ/zqCFa6vOFYy0FqKL
7PVw40SyYgGRvDWty2gNYIA8p7UJmiAUrUsMPSHeb57+qb3+uXl6IcFzGt64V2hq
h7mXRZEyR7LOz54dpmbt5w8gh7LlogErR44/Kt9llh95oLWK5a7tT33XTL5IunAp
NRUg3nSJ+ou/7F/ijn/D40cq4imjPQM/G6f/zw84UqGyCb+C12d17h6FbVICnlCE
wsomr9/3FFRfKDX//aldfhWZScSSwb5Yqg/hVSjTXq/gIrYcdHB/Cd2KdFifmnUm
liz3rN9DnR+52M4YeWfVbvoybfZzXgMxIF130lP0eyLfa4OTvLnMMYYpCC9rRe7M
01i3GKtbXUVNYlWTcyuF8Usw639aYH1VjzeY/bnFg9oqIhvpI+FbgAoEkZqgXuf0
fyjRMdVPF/G85D59tqRgw9liVN4mJVOPL942DUr3Ss42UIPp3KHc9EIGQlHFCMXl
AeBLruXuQRNfvWLpD3+v1Y5BX9TfF0e8WV9VHD9E5HKzBpLok/bl5FLNyiY982cp
nXo8U8cjgIR8dB+A2fsou555KBzNUcPB8A0vWVb3ZJXBLio1QMghqVYjpUHNGhU/
fuQm1cUWNyGrI3Hcb1T6lB/hCjvl+FqZPT7v/83uzjXK+C70jbRg2RpkRDHU5+Ix
MqSmo6sigHw2C/N3Z46sH9PxJRYdFBiRpc5Yv9VYPE1kWr9I9QTWSOxudpMSj+pj
GXiEq1OmPvSYYAHO94BSTsj7XI8/Czrt+7lW6LUB4M18HSnwuZqRuUkUyT3dGRZl
XnVv36PYSeuODcKnf8asZ9d2jIQCUJrODYRWTxNSiyyyqMpmjlspItAtOfgPOm9W
EXrYBzu7nhx/uTYYSUL/UScMLrrZ+kiSgKkQ+3ChKwDXumdomgbderqEJrPeM9QQ
m5DdPuuvEkovR2aTswcT/79zxOnOpTFAL2j9B5yA59DDDQtfFt3K5XBxan2MO5vs
A7xPte5+hMi8o+kM4VPXvOdZcuXtj5+nVcbknTWNyWVjmuGwsoQHuHhh4ji0c8VI
wx8GXqaq52XtFv858/wMPHnyd87zMxb+GFJfhzVC68imGiI/WVfEBkK194PVX46t
5aVRjdaIDz2q51H1CEJF02/KmAQWhewkq4rozvT2eYfiELmYKy9Bqctpv8+1vMyY
X2I38TO2i7WT724xx/LsuxkNlRpFpedPEi2kmvlpSvhu7GRvwPwmNrc5q8QzClKh
5HMjHBm0SfxLbzx1NOzHlaT3hzqTcvuqoY5VmJDSaXh7/0GggQtPqDHv4cimhh+Q
AK/KjhghfzP8wdMqQAz+DQO9CI+vGuFzhHpGZhXNydl7GpHhYdbxfHSFGX1WWxG/
9b2iUXcB+F2JqvctvH3rstAkJri/WyANIJtQsyJ00RU7ZoLC25BhQESp8PRMidPM
e/M0kRxFH5LuxV83VyG6u63j20BBPq1gn3kmAURIC6HXyprLLBEKkXauA1AnQDk3
tFEaH2aEm56ZxjGvIn76p7HV5jruU84PCY+cxSla1luVa4ocuFpGkc5f1HknAbhp
5G7c0zL2LPJxjBBH9K7Qk8PoMoZlrKLUZNVO4rE4t9339dw2t7bug3fCDbblJY+w
Ut9nEAYE36VCrOXtij63XuJlwfeNGalLStUf9A3RiT7umPPZHXR2wVLRjJguWuLY
BMui3tIIh0QSl7lhoCpY9ouEiu9pScycZ3o7YIyELUDupD5v57bMtPrkxvdiH3w2
Q6G7iMgruCxKBBHqbSs1dfgn4zs/ZjdyeP/G0GfeYkogYxsE0q+58pczUvSgH1CL
lcvEPOiwgx+uU132Ob2MLboPzZT46ZIT4gndsfM4E4vg+xTLYR29D2WUhI6QEZrN
J6eSmCqonKYF73Ix6Qrgl/aWIJ/PM8Hmc1OVBsPf3ds70F+iWuLGnGx659mS62NV
5QXLHOtgrPTf7OTy+T18znCm35geX1BQSobPo0g2njgFsnRccr5ro7zv70hdYBMt
qMBXpSw8bxxYXybO4SqR6RapNT45wjjefwSdgxXZmitLwCGJvThOnYwWML91rehq
xataK2q33bsNr04T8oXoBsKats5rzPKA+fEEy+nJlfWJq9LOf3Zg32Y3n+ThsS6t
jgQAAVms4i45/ACPu4v+rXGTBSX9RB1vEjOJQVuCiCpx/eU1r/rvC6s6bpPAJFKm
OyPkJ1DrVDoG7/2jpyS7K7Ar4eAJzMoYwy0krpE7VM6bMvaf32ST0Et75FHrMcDt
9jk3yNob/xM+rXgIuZbN6Ih5lsPVGJ2ZB1D3BOkqYzqS/dyfcuk8HCWLpOGDS9nf
u9xSvDR/2yxdQr7gujWpfaI/IlFFp6Qs7UpTAI7EoNpcoEFQ/ekNxW6xKKuCasIZ
kohXXG9+bnuAposK14F5RlXCjSsOMBSpqSBy7Q8vKWuwjy5smPo3U4yJ0Z11J6Kr
lvFvm5gUiqUyH2TSOPWhamo/Dbki00QTCNNaW+/fxLU8QUS4gAbXkLIP561ARoT/
xvEry18EQRzR5Roo0LVAx9GQ+rypbonjeimyju1RGMdLiNIrNu6EE1zei+pJMIxi
zk517+HpWh923Xu9Ekf3KzvkuoVOpHmiSgnqq2VbmNb80AarYsGmUPJyyyZBg2Vt
2qEUND9RVollo+qslaKDOIrfgvzYdzhvJFl42OUOz/dIWLPSAjW69yWD1bIvmj6B
xQKe/ZCssXHpSnvbH/Q/Ct6bsIugOvc5eLSXEI8gehFPEB9DaMCvTvkRno2L+fZ8
wdZn6wkWaiCAQY9N8ZdYffjUM8m9ZG3YnRGZzY3D8Qq80qmepr3P8PBRJupBn0tQ
tC/lNrreLZgedmUD2dsZx6l489NrcWQ0m59RBZ0x2a2OMHhpumUkF0G5u0E7aFMH
bhxAlxWCIxP4iOedOf9Zcc8V2hF/jtSCUMBGeABHtV+HSu8P5Bbl6ULVHcDTKOYp
1zYRejNQ9MAPlcz1dg8K7fDvKgZlpX9yB3oS5WviqPnFx52c6eXZVK8Nmd5301qv
Q/bRROQPMHZeOEi/+ywNKC+W61jvkvKTJZ0Ke2eshi3nVjh7EZDC4h0uHQK+iCpi
Eh4NNWh9FB6M/SJLUR9MuOCHBJhlGaAYb4shoEj+QA9INQUtc49vvGfEAuoJ8h+8
fw87QV4aAivA6hoPTlL67Tm5E4TZc6Qc1kPjFsPBE6+vrn66ScIqL/RfXHuBT9zu
Nf4QQ42VOw+vBbxIsuFsTDFe5D5i7FRkaOfXzHCSDDof0l8SgfEhzy9N0SzX/zXw
vXQiXjrfy6clWUdgZphlj6RZR/MwkuHCQxgRWUQtZl8obZq+1zHvAtpbVFm5VgYW
Q19X4uRvv/BTeRmWuiQ5qpnl1fCgc+0Qs+9RVwdvyL9w6N1g1LOHkOpvFMspDARM
DDZgVOFqPcdEWH08zGKyNU3YLt0jG1fqC1wXM/SkSmn0132LqMF1IjGDXgcibtSm
fV9MbYfDAwsHDMDlhDWfw6rVK1tD8e5pdElFmYlIzNdO5xPZ11HAlBx+HUCYBikX
hx4MujhLm0FTW+L1/1pZJsTjeOc/+YmmMWCEqiRWBL9X4c0+ptTOgUvj2pk8ebZs
EdfLl2YyAciAFu4450OE1f6mGX6UZcOCxIfhKjqY28a/bTyR2q4QzLgDhDh7dH4P
GtAyHC3XzXUZpJkWib7w31f1FGi6e0cV7lw3iR8FwxHEldvDLfTtG4Qxu6CiVbuq
LYtG8SZnyTKd4QUjO3vUq3G/f9WAmD/csM9708x/XYcurWSQ4W1+PcMX5cnt0Syz
PxXeZShPnYkA+05dXNJYGWdHA6+eJn/3cjWFKW3wxqWAYqRz7Ikig+6KZHZ7gicP
DqeKKIDEHu1YQFYZyCgqZCNHXttUyWomTGdrSH9yGyxdDAYpNdz8MhyOUJrt2Vxn
d9UwU4sBoPC9B1Sy4i9jo5KaHvAb0k2+kePL3fuzHJIwrlSc5bAjvUxQw4dFGJcw
R8uT1C/DZ5GP+kXo+iEbm+fu70DoBvvt6sFyornzxUlElVEbFP8IuX+KTNkYu7YV
uFihXDeCGHUP0POPBlWFfIp5KpDY2xsz5jogwdhWpfJei5EDjmqfUT3itpF3K5FO
Gx4hl0cqOcvpLj8ygPzkX4/hc28ZwD+3PAg2MKOjsEKGVAahBP5vXOWB/UIJyoCb
zI3Y6tl4I23KjtX3BL+aN5iIfbiowf4gpZv/d+SOh0HbrruDfSAxjPbdp4A3yPgS
H90E+iosSu3/LJgKlWZChLmGdK947FJGJblacKOrXZ6qihtQgm5HwjMqHN1Dz8e2
m8BTE6bAr8GvJIii83vq8UkD4/qeFjDfs7w5wEdBtCp8/BMSaTk5tU1BocunUCgo
aK1ZL6dcoGenCvxhCz+G5lsLxBgPp//N6WwmH/ZlloMa47Gi2iRkDs2ti4CeBUEd
k6atrsmEYrF7DbyAj96YwH6oYU1IIPTG0UlnI8B3vVhldcxjLg+JFmWIqBX7l27i
lcyyRsWKQU2l7eRxnaCel/qpxh5cnelDM/rr6ICYC+DfqhTEkLMJFwwSRovqeKyp
ZEmLWcfvyuiV9Cq7PCDGh41KGHHFdMSR0IDaFOUmHHH7DhK/b5F2Q96G1PnNzN/+
ClL7s8qSDfk900udpQSbkspv45RFJ4ubuyotsV0d1CXodsJzY9AK7SnF0wkuslMH
zG1POs1ZSG2Zb5SFE5q4TYCzrR39bj7J7gsaxDym5V1vKkQm9mXm5key+vOiLaSb
KVedXTle0QXc4YvKIEysbN8ffA4nuZDWAd5w+ri9yqcdODEcRTWSpkYProvQNWhj
LzR2qh98kE+arISel9UYyJHzFcdCWKL4d+9p6PGsRZET2L4nGOsK/0KUB3QSNaE9
Dg4e2Ve57Kab/XzXG2T+g6ug7bJde9CgWEhGKlVTgFPq71dJ3lAh+R3gk2r2/w83
4uhAdcQMrexUmJrPhotqXln1IYMNdWZGd67ZFyggFtp8fU+HPIEQqiifhwEe3bLV
EXyBU9QOU2oLwiOPlVDfL9UZpozutEDcwWzjajhJ45jU7vrMGqO12z3VU+JyT/eT
TMNiHyVuuYkszgHJFDSEaHpjJdfWriOpr1gaYbP/BdoC7xOIqLJBgw8SuVlRa4PE
cuQq40QqVOhwYdMy8LnEAroDEqcUqv1KTiwlsCwYULAqJZs2MNi/9Tdi9OR97SIS
95zLV6mY3r7ukWLnVOz7RVaC6+Qv8FMn39orEMx/sZQyJE1aIuJiBlaTnTuDpX1V
cM7I5xcEBcBKYygAbXPp6bHJ7NQ24rVgm1wI0NsvOXk7zHdIWZhV7GnoE7Zav3mi
qj3jWwFCTVSVzYoZytzMJqb9yNa4kozCFaVtH1lFqs6LpvCNGxkC4Ev+R/N7Bxpj
xyzfxboBDYdeyBTcmJAMIjC3medzGJiVynHuhIrmERz7Cqym2wjKNbRteJ6dkYyh
sORtrF73QIwDphy+yX7sWd04ak34VJ6iyFyY96cjcj/+W9/FGzsfXl4TdorVJDx6
ZxHoIz5GtLaUw+XobDdrp/S819E3ooZDl8s4hPyxKsMDISdll4e+Ewp3IQWvGXi2
VNaas0x48mqScO0G/84sEMx2kkdKKsa83ePN9z0jiz3kqUe16K9zrODiebMq+2qW
As3ARLWIwpWdK6OVlr9d3U/CO0RcTPlAjHvqIr+qq1vjOKc49Ca2L7klZlMqopFV
s3vJauzi6g5SIggINg3+snLySQGbCl1P4yDHgQCdZ2f5qSn3SZ5mO/I4IEosoDU/
HY4QLxR9KI+5PXxsdKMxC9001f/Y7wqHnpzKXSR4iHbtcQqBVQDZuHySI2TFErDJ
BfNDr+gKDKcm+S0mbTkQul815A1MC1mmLPjBABEx14bxhhfHQTDSH/cLCjRRlDiO
OadzkoyfPiG66So2AXzoAejSrWj6azQHUOyX/Ys/12CtCCHtMRz7qh0Fmnev43Mi
o9/mAyl21LDFn8TKt+urgFANc1GbPkzJQS83V5VpCKvV78a2+uMr4Wq5SNpGRqyN
fi8+8Ewq5KeUzynfstV8oIxCEATaix6wKXJO2WqA2J1Gr8qi7D8khS/4VTv7SapI
nqMse/9IiJwGRMmoAWtJIf8BOpF+Uy06Ul8z3/dv6HVFy3GmRUUe2SLylGIg4GKU
iSYMSTHlySJjYPIgmVzqwF54wM7kvamL8yDfcoFsAzUaXlkiDqtbb0OPgtjeAzZJ
22XRqqgH2b7FT1xM6R882xTHbPvaGNwPyQpHmCqUxkf4VnIPW/cTP8cpoLG6YrzE
sb8qb2NUBUXXI5dxCPXyIc67g7Ito7OlPBEe2qzOsk3gaYnHTTFI2B0DyWfzRDzI
oFvg2PRmhUvUNiF3SCj9jDgLUgU5Qam26bCLWoyO4iGhDIrgCVxjcj2wm5glYb4Z
sL0afy1+hScykhvNLtGyATAQVo6HSb23bpLXa4HScP1S4FiNJg40f4oF6ceLVSL2
PVFWeczw3Jdk+IiTZfivOS2paDpRXY58Z89KAe1NK5IPdqS1h1uTSR02kEUgBeF7
MRBLYoy3hl8oexNN5tn0NAeFP23waX+Ff+hc2/FcRPP9DHpj+ZN4XnocRnhoYRDj
6wa8045Kh9TcJNK4aMncK8n+nbEJ95uYIeXicaEOFdhs4Illg4JI/g/LMrbU0UuO
ktm8uQL7qMY/YUN9IjEPNjEuhC9XaSi0VwWyBl9Lf7QzGgrd/0yf3elm70U9ngve
6c2qCsJV8wI11Gmk/W9+lajG5S6ri7BjLo8sDqZCBfVMvLdxDPKkuHfdU2iPToCM
+m2dk1DhxQIPy/P8s9G3sNavny+gwKbK0ftIKTmLPRo+Y31JE0Ukz6e4/bJ5einT
X+a5zG7x/2q5R+yoe00GdomLJXPPCAZgLVBfrTEDe3kopS7ut7smG+w/SCOh6UMe
NWzuW5pNLGe1nNlcFvJ4zGi1JwzDxjeBKbGZ/aOIMF0PEvIAMW76tsPWggogU7pB
w4JsDxFnr0//vbRgtCrx4aN9UwkwzDDOcOF+Mld7oiXEHDURfodqxusS2S7SnEhA
40JY4BkNmxuZ+arRJTsFXbbGF57MuSMxnyLPfttVjygCSrUDNtz+TvfErGd60Cbp
5g0rotEO6RZvjOCMDBKQ/RlNU/BzsD32X/v8y90E1fXpglxG9mmtMWW06XY1xobU
ENcU7jb11Ri1e3k2JZ/TlJB+mjCPLrHIenHhjCRH8pt5KJhl/Nd/MIYjxoiE7XHc
q8g4ZMbR8OBFkS3fBhik970a/mbP0iLk3WARiBw9TkspAZ+zXQH7IZxrE9GFld++
SHAPwatvCAPCSxraJwMFejSD2zfWNTKzdUF75iymawBEE/sM4h7M47elBpmZymCi
259k/pANZuKlnTFf31YlT1T8sP0MdV3XWqtcpHPZPVdZTSmV3YAG5YYt2YkFKxs4
YK1VwdQqBu3AGtYHjANaONINSU73YiNhMvqVpc9XsDOXnywbS0z6gVDvfYzWcNbc
EPc8FdSpA5cTME3h4QZWNQomtYKmFK39QkHxIv5ClFPeEc527JfuGBSLDDn49xGD
LsLXZcqdhg8eS3cdyiHqGfd4TmAe3KlMVS6iaUIi5Zbmjn8QpMqMUnwwtqightRp
63/EVZ4gASZgC7BfnYKswOry5Bm6kBjfMr6RzJNOQeyOWoG2h4+EB3cw96Tag6E+
TX/ZmKmkZT+4pUYq05ZtDKdSXYaDFA890R4ttOqBwx2vRhehX9ZzKwniNIx3rFU2
/83D2iKwgKBbnKdHn16K1UlIYs+zEkYONMC3y4e7GHVhjZwmyBXMTju8P76uI0Zi
+Q1uWOEtWd7LJ9IILqeNlQgdjQ8Q6yGS2TPUrot1oEIpvzC7zce9rV6bk5FOAp8h
fZH/RL4UVR8EsIWUMJ1J1g3CnwRmZliQQx/oDci8AN7M3F7nHghK0xRXZpi6G9NN
bYL/m8ovN/I8Sc0eXrYbsiwF14wTYZuX1m0/P6qFHQ6278WA4st77cJtGLpGNC/U
lvML3KgSFNN2z5h2yi/aZEYd31fOjIeFWk6Bro7zx/Xc50LJ+FvF6ytptOvF6IFn
cRHJQ0D0eamIJfKvARaofsyMps0csKMaG4CnxWKmS33pQE0fFKoqk0mo5mmkGKch
DvBu5MArs+n5fOzrCu5oI8k5NEiyZgdleYvAVUH9yMskG0+MQJXEqP4RvhFrMh/M
BNdeVLfKcIrYZ7jqaVG2ED66PBdIWSzHaZTa8e2qozjIx10KCJfYeH1BnLu1AadR
WxvTz47gOcyGRmkUxqPkou2BVK39pAeQBy8YtoPA2oabMdytwZJfbOLV/qeWRDZC
4icriI3t03PAU24OHOHrMGZVc5vnRym7df8RTYN8Es1MxlUlb4wVF/Tfvz6/G22x
CTto3nEd9JZhsABrClhm8hIPA9Twig/h8EPOfXRFkuiaUb3IoxsC2aBioLHumCPQ
TYIEm2rEDhFQlJ0h0Yt1VrVkL+ZOiCAYGHSSyMqpN+Ul4Y0vMwE4CbA8m4GfQlq7
Ps8bGkH9IDca16NnETrMbujl3p/fR4MnSzGZrby36qfHh6P0nIxQoyg2LJYkgCO8
kXAA4ZIhqv1DaYR92/b3Tt9quJCotxvyILfDqCesaYWM8Gjh5iovoV5FvMWuyzPi
wtMFGQU/9HhfnchOadOxgNv5jt33aniEDed+8EeqP9Zf1IYC92S14nGQQZUU6eVa
/Wyg2OSBrK7cpCtHJyqP2FcfK6PPt3WSTzae3mZEU9Pf4DNEQ9JqhxPbCAqZF4kY
hOboI6QmpZLt81diCPBCEA+Q7U67CU4E4rg2xbPcTiQNe1C1ALK+o/sxTW2NXqsJ
Q4YHgKEa0RmMdTL5DWvXrJqlGUZecXMkAa8NlkBGR8891PBnJp6zVdYpER24w9iP
hlk5jJlu19zD1LSYi2cfQ9jaXxlB4MhxthJy2W3ZAoNPfXc804cr9BXg9hSbVvXR
1i4IUBHHUmu6laOzLMwu6Dlvyg1frls2I7bCr3USRGGuqFnHDzatn345QcUoy7dT
CbAkMt60Dc6FXlDQBDxai62Hj+SOMx9NelMCsYQF/ebyesSjIvD/iM88rp/4CfZr
cGwJ/7cEAiDVuG728YTPqra2lBkkp4ViW3Rj/mYmGS6GxvZ+Hpmoetp/T/HxNsCN
wyslKjnkouMBG66N2U7SQ2B5WCRxVmME2E8iNjac5sCjVyG9o/nXSuQy01xHMBHY
o7DW1/xFjS9yjGRo/1A7ba/XU2PDFpsYJwPMYFBDa1YjtsqBqZSQVS+RmuuFEPry
qDoIjlyEsPTgD9J7pwizjByC3uzBo3+rS37NkMPHZ+Qs2/VWUp42TGvW+Enue45x
88EvQ1WGpyRQQM6G4R5VizHYgQSW+rUUcSemSLR66Li9cYBwFPc+H5ZrQvHqYfAQ
SDR+z8ztRUqqtTBdgDtQjw0jC3t/171c7NdZqG31Yl/rX9N9kaQykDnVzUIgG1PN
mDFHB2DcV6wkeY77g4e7ic1fHK9AZxrL7TItKDAVIRu+x+Np2prvMFUA+wCWp0eU
DEx8RHunkoD9oOW5nXC0uU/rlhAE8fEG+8BebHnlW/y9qhbWYB/EKk530IdmZiQO
N3uDbo1jp6wuHZ/6OIu9hWlv7bnuiGb80i+DERgw1ujeHQx0wLdsJrt2NGAJ+Rf3
ncHwKdEBtdWULNg/G8H/Zo6bna4jXMGO+sfGfTucH+MsBfGfyH7s28tmBAmN9CxZ
FQHUHG6MpW5d9O+uyiD9n7VfQORzltJNctLOVlOON51dZoK/pkLPie4SaxBBAdAf
oSGor0TkeOScekzMWvr2D9wRFF+aXGTo7w08MIqI1zaaUDooJljhvxkQvTcduZvW
8FTGKB5YoKLCHluI0qcDQjyi/mEpbQsPtUIS8ZMbMoPJ3BbT8Zys/M7RxxAO1Zlq
DYf2vIqHbSveiWxfbiBtiQEHv5F8O9yUmk5nna6/3+c0Ulydt6N5LcJMz+2tcF6/
s4C3kVfc5CDrxlDN3eMKnTKFL89jlZA06IDv3Tt2wgkAw5uBhFChWoyGIETYzbEa
H+GCSuuRQsedcAgiNSpw2n8qnRLDz98SvgjNHz3fcnNK2uOXRR7MrQNClprydnzL
R4UZeQWUO1Xt5CR2SHQphBozh6RGkBVva+Vgq3mYYs9Lbzxf0GWTPoaV9s+QqVp3
EIeNeoX8I1Lxz5ZMflhXZapbvWd3KlZlZagi1qmHTEny/7wNv5SIL0jNRskcRyRH
Eie/WuifdKRepPiiX0EJ3RoWwiyhd7jW1NQTxx/xP0gZAmk8EjUL3YlXJFuQRLFj
fjhlpGQt5xWRg6daAQ9XeHfsdOdehIZlpiNoczILOTmEicvbdf2Ejt1eu/CUOsj/
YCAXb5bTR3H3TaSaSAWdUv99ppkupTXB6/MErUKPfYFbavejt1thfTcwSvBzkhwZ
IYxC3KRNlIqRDzPssTVvEjPA2yIIdr/Cq5SNd9SvN79yJCGXzIzs6uRW/o3C4ngD
ByIR+km+oB2w40KYlHMMTwdYW+dlPvnE4l+ojjJ27eta9EcwgSvfNBOw1QDER3fB
plimb37nWXCFYhyOndFGMLhg0g9WZ7su9PWOU2uePHLen0CkSL3mGccQPKc65hwY
sCncVJx2OyS27b0I2V0Urt2wZWktkq3712+hIIC7sB7BTnaQfMO7vSY9pwdvUnVR
bVOW4sPcGaOL/mtY2+tP91FpFi9bHhp4HQDA96LAy0eW/7O488R95rEiBlvm8k4c
4z6Wl3iJ/gQ3Q9JwX60/08ZNTC7YznHt6195jf3ipwFcchX1upb/57z5SyXR5xHX
j/kirar3APjzD4DA2gMfJqzXiW2CgpuWWrPBzLIHkf2oevjevmGtQWCsMTnexWt8
FB1QUdkigQYoUVQfEXhns29TvDpRirHzUGdHJLa8z5AZwo1st2ddvIdtwX5snnu9
1rwS055pjheE4R1QBPL9B/BYKmPYw5aHyNeHeVSiB2P8aK79w6lk5glbTEQGSHYE
pRd5U2mAILxdN17U0CJCj9mj8MJNIiH+PhRMsPr4rzp6iBzqN7xVSgtEKi3uf94J
LC32EQybAs0v7Xdiuy9loC6uILuGDAcrpvnxfdt+OAtX2JNdruP6z3rkDDTyXWem
L5aqYm4OG4E2e/dpNZe8K1Zo9FkQAaXVGhtg3JQvkxg+ErhkgkDV60CE8XSCjHtN
44tJLyiPCU5ioBhlNiaMyQou+8WZLVM9sQ9GBzgg/5kufATqKuzQhZ+pp156xWfX
0rFQrI2jglvsPFyxOiVvTRVf7fmrvY1CxIuk098oBAhpFvYG6OGW+ukzPP3LF16D
zVHCQjFx85N2I030ZqrVgpNuKHXYuNHpm61Z2qMuFjK00gsCWcusE/mM0oI1j6sK
GiVcCDQPY9dSmu9eWploiM1sGOVcJlUJwwhlC1mUgou/kJ3VviQJRqonpwEP7vfn
vsb5hS2sYwQctzQr8MGbw8e5vAJ4zjnIADVRXq16fOQpEHZIxcAwrmBCoXINahM3
WlWwVz8MMItK1/VUn1u02p6/RXDBNi51OWgmvz0S/Np+0yxQ/I2mHBnWcbwh4r4b
ANEnlbp0cnSajHmmyOKbaHgOim0o0gk/mrz8nqRcPeAK+h0cJVB/0rNseh2G7j1c
F0c6PCktL11IjLIg2NKf1PkIHLjaxoTtcNTdB/ExUVBOZB4/davTfH8Oa0zrE5v1
O75HWeCpw4yzLBEewWkfHm8omJBUCb0FzWFo5QS4RGc3xyM01uIQPiPWdcaMFjSW
6Ge0PVOKF37yV6oxW2Is3VqYlk7591uX0tivbeYdR+J82ESK785eHzrucEE7zOTs
lzzmXz9u8OzLleUFeRKsBNsRuM2nYOuQyX+5CtZ0aikhDF7KI0Fn9wiJ9J1/XpzV
vFShxYEFeFqa1jdjTujlbGS+RX89mxIt6Lc7kKC3znjb9ZJTnDqfXVgmxXwIpi2E
gBLEuIj3fKZQ0CWZTwzWxv/Sq/G7qq3MY8MOZ2bit2Vz3HL8nLXNyGAkK4RUkRgB
rxKcDcW9Dj91Yk3tk7TZkih+29ZSXqJt51dwKPxLQXf7p6Htvb2ogfHMkCTwqJRs
UcHjO/SnP3QV3eUBY/UBhZNOq2i5UHtHtdX+x8Bj2qFUouGQHphjZtI4h7l3zJ5z
4sleGcFgu0gH+7cOLuTBlR2j9cUuDPvweIF/dVCKU/JN0TaOsFhBgNIkXBnfgymE
PvWSkGjzO0oTEaWhdpvM5ksmWjbGxk3WRGmRIS1jcw+xXV8HEDCb/limftvS7329
UeXW+UAaY7mSDWr4nuNjQYFau4BBlV6evx5RSKak/SkPQoFw1EI7qisZNkMT6dI5
/MzVYZ8MOaYDGXQFiUHMZe2RrNrAoHP+sBHOUrkcK8WTlR37T//c35qgZgF25bGy
d1PHYkzoYbVMJ/kL18Ruy8WSU+fiTQbxm/ukTzxZBb1nRqeF/UsfvwYl+i3Z/3pW
gx1CTPWhJOftlNN+kQYknxuMRRxonC/cqeWKi9opJy+J8tHVg3dZO70EeYw0OfPX
3Tfpeo18HCQxfkX/ou+XXZIDtD9wg0C+kdV6keD14+MrkeYHLbvy1NtqdquRXuxT
809tWHT9WRlhyjGDJqmvU1yIOgap+1Tvl0Vd0xpxKQCn40kpvGcv8kJJz4pj6ySq
2GSrtbobbt+nLgZSuSIXMIdatylma1ZnpkbP9cY/hAYxYLBCQCB6nsgjsj21Zn58
kZLRGSVjKDeBKpHrr886HtpM+7EMbd6PXT3k8y0kiVGJXk6FP21KLl7+eLKlOn40
5ECUzyqCnyvEiznycGHh/y7eAU0sl+8eFeZLSIKlSDgR2a452J86SEJBGXxcnTS4
OAxAbJ+iHu4hMDW611i4wJkzfPQCEqtXTeesY/jAPfxu2aRAmnjh/mbLOn5IoOP4
cn/XZd2VvtieQaBdINYxEnyJqK1CE8RpjsoOERG6EHStIk4KxnwJWYGs7HSlJKhh
zeLnfRNuTccXUgMuSn0Vw0Im7z7yeTJR70tvthecAE94ESQ0bE3SjilspZEWSQks
wZDidFjTwUpryAfN/0RkIUTBPILW8g9GzcPF2C3Pzd+P8mN7RT4Ti8N5dk2U0B4w
o73sntuVEeYQQAgTD24ik/2mrjsPgBBS5Dv2V6AJf6ERnBMfJbOpE2Omphfidm1y
Hp0N1DC3CFF47aWJY5FXROoZ6CmD03KLxjTvBv702jTbWMfgCL2Jj4srr3N/gaD+
WRuFu7l9BYDTQD+yy9354E24ky189j4ro1CgdU+C7Z+vdM5rtyOoW6GBJxsW6R62
t7YOvLlhwKfGvlTFkvoAiHpO7ctCpziHZBZrtK+Hh5bw0sx2gY9CJ5EUFwIZ3Wxz
KL3gyUSrHlEQGoINEJQJPiEQDBjDHEuDZ8POyJL+A3tgyOB2ZPhyNKJgwtpPGmCw
KYkbAeAcPJRb8YmQwCjLsxfxkWcb7lEo0OJM5RUdYwtgqDpUMNjNplujcub/3hlQ
i72rSdgj1vD7SpuWQA1TAT5t9mWYhIWCJNPL/LNi6Pvtnd6+1jC5Xsfx0YcJbjhn
72M9KFnJZPCpRE8Yuwyt3qEUOvUWw1OGV2QolCklsvYSbnRzDKJ2gbbGgQLxiud4
yvlZ/0R7cu+MuFiNtn9VAIHpZGpHLqk6yN2cHnXasEqfGhdMgGCcbEdn43/RGY58
wOGg61GKF5Z7bytWXRGsrPKua+IchDgm/ehRH/boHxc2Z7Ge8+CLZcazbuJ/0hYy
j60L2c8IzQKvERZYR4JHC+lC2E2LoEmUCoBTqAGc7po4wdz0jlWAGMUmLaDVBVVM
prFWslqS3h4YjjvVcXJEp+d4rcC+BdRiVqrin5XLAgdKjy/K1xGLWHLpvHaJnZbj
vF4YcXb6CUSvN3SzNomPc2hrb+WTrM+xaDBKQce5p0OekdiG1ZZbj3geZf11kWdC
1KsCA9m60BhZnOiNL24vy0KcdcgM3rSt2xYnLv/vB75y/w6spANPKx2i/DSpE3nP
9jy6AHLBrdRMcdggnchTHl0wwWj3FOUb9+d2+xT8HcZ/MRebO4JcjUXCgicnMoxQ
9H1fLeN/1uqkSfrEJl3fXQlljmt3w8XhrmZfeN0a36p49b/k13ExtUUhJzQGXG5I
L2TD0n3RcZ5H0vhoq4nb5H/ZvfHswBeF4Iqbe2a4ZGvohCaWlre0vmKbQP3Ic/4n
dcYHhblFrEGuOK4OOx3K34rtowrfODeuz4oUith2nvAPU9EiqzYpoD96tknM1jNV
wLepa9l3XU5x4j4bdOOqO+X32pRskP3Bgs7O6SMgRjQZbmx//zqtNu1tBIonDS6l
51ihcgF9j1Lde0gn/oX8dFcUaDFzLFKnmgPCU6OgpXoSRvNzoSdR3hlOhStw2mGK
sOiA1fAYNkVZPs9m9HCQ5iMUznh8DqOvIxefVWXcHS+jrzskRYai6CgQi8GpCZG9
RGHfwzwqRwoya886qYRGNJJ1Vmm2lTXvyWehcTP/zSdoecR2bKlDpD8hxA9rmC+I
as4LYofMdHPogGJ2SfvCRZx/r5BAdAltR/qp1LviOI9cRjbggf0wbluzrccAO2zY
Bu8Zo6pgX5YtqAiRa0Dqsh89spCIlsMOB7Q0WFFSQ8O37h7wnBA0me9soKKiH/M3
OqD/DlDIk0meO2PC4sZJ1wF47KikfqdcW6Eqmv2Cginnk3EINIR+MYtI/s+SIs2p
cxmcsWLqy30XkrY9t5pVktfMXbtes5D35J1hMj1gaGvUky+2bi9b1NC1Nj6PDNN0
ftOuC1sh5CGMSDWoTWIjEA+NS3H7Rl1vZQjztazDl9rM3p8QMebqNtppbZxjqvmv
3ZEavFadndxJYqRuXwbxM3jroQbhRfkdnlEE3LnGr9i5Hf01XXLo4FaQYZgmku1D
Nifdkd8SNddvLLv118Ns/ilZcnZFPa4EvCnvHmPQWVRnhsYRixMg+MR2/GGV3FgR
v4ypa7FI5b2PocdHMSFo2V1rYT/UdmbCnFbVGnoviGfZs9zJPYrdT0IT56nXa7Ut
MbJ+jMkFzIUR8Mj0iVv1rUyzfimWxqVAAtW8Px4fDARotpjeOeuUhHzZi06LaNzH
yKsp3FRfqBsLb9nkj4F08CKO/Ekw4Xb9wFT6MwsiB969g40OV9lRFLN0Lp1eY87Q
azGVFSwFkIT/4/u13KwRdrFeOQZkBxoY1C8AS7KHCskIWxQS86uoVxFH+WkPxKpT
emKh1InXZ4INCITP0OdgoFyzC4WOtchP8Yx94mZS6h0a6ZSK3pyQmKr6eKPAb1zL
TBXLbgB+lk/UgzLdipP1K1m3oC0eNQMFq5AwSc3c0SpQcP5DWcPev6kcQsh3DvLE
Txgr4QfwpyhbViuMKohXZl0/R86USZZl3WbHd9pebbWsNxfkWR/IJmaf+xz9fEWR
eMVIZ5p3Fc20eSxGLdp49tdIU6n/FVtgFHYUUC1fQkZ7w22OZcU74ZcNUUUTdJxt
SijZ4l7c9/Pwd8Bo4qW/AD6JpxMp2hZ3+ewBMB1GVhpcd3Tn3IxRXVa9ojARBqPT
25+LU5c4cbSzhuX/GZPzHWC3pgz8DsxfhO9c/80voGknQS78wqaKDwyPOnAmDLCd
SrjDWFJVwx6l5W9grU2M/EkdIGZeQ9pIrL3GwpSu1qinC/+VaKZUBZk93nsyfEts
16D32T1ZN/ELbXXEFrhWFQq4kIus5AvnmCEcfbmFABqSVpAdM8eOm14c9jwfG/vW
/3UaD3yDLMbGNaBBOGmNSSJUM024pYpGWWMPLnpj4zLcTdMoarO5yAixKwGN16RQ
9QENiHoDf6js3N+51YBCk9xHgoQRmI3If9viAZVro0wjW2CWXypB0dSNImQErtux
JHn2ttAJ6W4pmPrLyYAl/73r62ysQGLxmTb5Xsn470WnCmz9e7fksn6ChF5ZtJz9
pGR+jk9J0bk695fk8pA8cA58ts7LzRPP/ODHm/IH06bUqD+pAfpc0JQ4XuHXbK5n
nV17IWG2vJ30mOvfuoGhhtnWj4PotrMXXocvDCT4QBS7y9BrH88ka+KnzixgU1Sm
fNwzID/1tfHIHYAC7BOfuTDNfI67nkv9SimoU55ODQjLSvylve4mEZMPeOX5pf/K
/upMrnPcGf6o8i5n5RZR3WyY99DkuyseUVIrVQKMh3rphEzs2Vc4jYnbh/WkMInF
Fa2KVij6by+Ii/O2ti2WofpttX4RWseijkcetNp/nPpzqcl/KlsCS5vngCBrNui5
Rw6W4OL4phQ0mEgeRkrhi82cUBqm7e05ctauBMtbVz7B4POUlPQ6TFijF+RC0h+K
aVjmt7ijjxkN1hDGN77CnDLIIKxGNm0l6guRpqDkwXj5KwTeFTIpfQoX1/oLkHXi
G5l8QH/QDvHLT6ct2K9cz8r8fOciHq29C4PUHc5CND4noMkO1/BupL9bRSMtxJRu
gFMlyhTfbstCRG7no48YeQvIHWXsxqohSLwH8ZBe4K2KluvN3EB37noI5NV58VP5
L5XFPphkzdGVTK87/e2cc6Ja/X/19wBvCuQW6cXHvz1GXDup6APBAtm6BrZrj9XL
n9buM1t8L3ccRLTdoGAAbmz/g83VKs3Et4bFaQb+pPGzZwRKtsZ12sdVybyIA4R+
8NMLUS/Yy425GVVFD7z5Kj1UsA7KNgoWwflEK9h45c1Af7u4ijHCTkli93Rl6JqZ
zsJ8draafXQ02KeVIrfXAOw+1Twll8E9E4WwDgEpkIR5KuN+ySsYe0cnR6sLwdVh
2zVZqZIoZSnjQtJcdRYwxiQct9VBZAzDHQzQMByZJMYm8DlRyYI9Y+IXUjsREMWB
HFWw5ubgHAgnZLGJqK3HdDvb4EOGVJL1wC7rL5mwSy3O5EV9svzy6olNFURbUb0G
RMsKW0ckkoCQlbAWcfZuGGD7ma91YIDS2oDi4qSSlFoD5TCzZGTTKJRNYutsFwdn
wRqjchwX+S+asqym+8wghW2O4NYfbRp6JKRm8iwqhFybgA0tDzsrXVoxq0yfRyLS
jAef08nDzTRYT+BvjbV6z0XMYZRbWOl6caekVuqiO8BKRp94N+qwQpwZjaBdG6ES
PcT7ovWZKIO9KY7yQaZQxAhPXb8hOdAiVm4OrC6174lo4TDNVXh2E1vu1Wh2PepX
qUjXCRVEqQse4J7D54gy6HLdocA0n8ausk/yDEXaNOBz6r3jllJgJPHpeQUSrRdV
IzjFm7DzPYxaxwwX6HFRGAZJzsh+IVQqDtXha8pg1etLg/uzbtOHfkt7GxuBD+wh
2vXcjP9zGHR1CfPGvJ21IY6YqOrqSUcFF76dc0zRxVmcDt6mCDkG9ZvdP6OoJj73
0ZQ2yg2Wu27NreX9uWkKd07NmH5VyqvOAQhSenqsXoLrwFXKquSYOfAt7qec5Y8S
ioasKHImP7VLArYu7BubEY559htC5+UKXU7ldZdFxwUQArFTslup+pVcgv25XgW4
JJZdypT1Ws2HCoWAg/M/0wmgjOS0hmeFoLd8bgDPZ+DPZ8XUz7qgJDtKQRpaznwc
cahF0t0AtsOSnwmIuNoVu7pjS2sdI8wCG06pFvZKyPUUFmGtZ3V/H4amCpKR5AqZ
jU9UDGvtOxiqB8+mPBq+vn4QJTpuM6R1rDiSmGb8L3aW7g0uZunjK1pFtUL4Lk2m
daGHzuU+WPVZyGvewvrXi7MkP5m752x1tQMdFttpCkSqrz6SIlCshU6RE/zT/Ecn
uoAL+YHHpmdx4b7NJkB7yJCd6Lf6nV13nLiT6GTq26HOqGtVPPAhQBPEe7lpSf72
eNBGFjGLZWWA1vH3xRLfN1VjBh39UU7WmFfLDlK0Tl0RVcKjjzRjfdWUccdMyqwT
7gHgw/NP9IYkPJJl+/m/zz6/+Hj0NlTwv1zjMOM5xXW9SKVzZXKTe/SYu32ros2c
qMSLmasIBmP8l9byhFrQzWZy0mXOCr+08P/pAAjfyl8fwcvaH180zrXDKFqNnvWy
QHJ74Ne5Aw81b8CK7Sx60b8U+GjltXlK7MIQuM7CxWusTglECIQRcLyXnEoc/o4z
XT292fwZT01OE5EYg4TLR7C2oKJaMwqWngcZ4CT6PFTb+C+pjrmVxGxu0HFYDyRg
kof0SSVo7bEG1bFehXbC1FVpBG2UVj+bamkaytFEupvOzI9zwsPn9AgpzJSsJQTH
E4JTtkbVSWHoBjs+MEtKg2DKeW50QBdlG7N0paYlUNH67dvy9XGig911h5vc/p0H
t7yK84fiWxIhWyLP23TOFiR4zRVtPSico4/qRpEFquSIiAwBtxWsEDt66nQQww8h
JAxAIQ1At6PfMj0Xfz0F2tXGhyKhRg5+ep+7HpAanj8iG3LjRDSpoKlNcIYe7ZDm
Ln6y6zWveGJVK++QNTOOy3kp6lcRhv60mUduQDA/oL0Qrclwbh+i86u+YOYb9QYD
NgobcgNyY+XFgz4g9i0kQ38brRgEYER8+xtSSKv9jedeIBbe15l7tZGGjn06p6nk
tYp2j6xOUD4UHujNdezvAMIEVVth1rw50veAiE2meKmM1i+ttxzEBo8gyiFlHv+6
LpBCVakdB4c+nUesFY/+AU3apgWeJRUhxVgmJRACSNaSD37hdKtmRNvvtA3SQroj
uKrY/Q+rHWs2e/FRGjB4CyIVEiyZ3FPuOItoycb4VRKGjm960yBLtpbe5DLdZ+SV
pQ+i3G93KxSSBtbW6bS9kq1yn69+5qWeEHuZU+kReTmLOL2KBhS5rZB35z4EPT1j
Th5bmtxy/J46cxoV43t+TXnEMPeWYXvfu40HLwxcg+xACMb7EMbUEayXcDrpoGfk
tl37hSK4QvQEGsL159UTneaz4pSjCNU2ll53dTlSyWj2T4bKvIwHHP4/bCPXr302
j9DURI1N2Z6KuWhKI6pRNVgQAJi8AxUkLtSW8knW8i4zHLhvbO+mBfTZw+OgpMvG
Z3OI1ZwjN2XqDCEDFyNH8SIMGmz5dOrfxwFTI9IS5vXE2gj70iQ7coG2WL2dtqZQ
7i0QWbDNDH1h1rDQmZMoVbI9HjTJUnUDzu3FrIyMCW5bs3ku0stZqkbXyF4iDW0q
jxeq4NAOzt7oDe4ZWGhHeQfNSVx60nhAEt0WNY/qyCJBfvbGM2Hxd63FIJDUYn05
E2WqoWQH5Vsnxcqu9J71dvE2TPhLhik6P5EIKJ5vhKVaZ6T8rjrhhJYT5Y4Zim4a
ZUYTZPCv1qIlabGwvSheAYm3J9fOTFXVFkOpP0hxIYwI21ORslfmfEosZI5CxYI3
wmmSdzSW2dN2SpqanZ8I2hZUIkRel+aJ5kFR2I+3tWsnSILLMEJhgto8/yw092Br
k4rCxqMMlhU1z4O53a9DXvbmwhXxvV0QRQQNeTt7u3gSgctlwc3B8zyIrtJPA8aa
fhN068Re97Mda7U3eywhn/vUgA6vbirOxl8zIwMaZAPI+u/8SmkEYLOu43Q0CguW
EWWVndRSSu/lfMPAu+5QvOc4ueBNrMir//dnJnJFM6M5M/R8T+Wregiv/MgqRMoT
WVT7WjYvypeUuafZw+XcZAQSPrge1tm6wt1JQP9t/GGid2yz+FObhRZwajvdvo1t
pnQET6B+NsJtVKg7wtNNK/O+ROgYmkhOZAJLJ+1dpmoO1lBKi6GgC/RxIREpykRN
7tRpqKfyo6uroZXNzcqnXgaWII+V4D2wZBF2p0bMq9fUbxUqNCaWbnZSs6H0uYIf
rNfS0aTdDQPYmPN70lBb2XYAz6DT063/mI8sqeOMSmjMI1tl7I2B/TLzfSiGcfXX
Gf8AAwvW44/om/H4hdQkZ9+5JU8nzeum4ipVZZOPzEVahFSBUrggrTIaeiZuPiPN
/wFJ1tim/aRsViuuYjohfJxDKElnzpEL1vPwxESKLxiTl8V8+Fua5nyhBGm/RgDM
tnemmAta+WFAaIzUF+AWnTKlhfT4YEpdM2SG+wWG1QguD5A3yRSLJ9x/GN+PamDu
9vohJ7itZjx90H/StzwYmh1Ns4Dd0nxT5VIzS/Mtnyi6NKNOx5yKRfVqI6mvujIW
FloV7ilkWaguT9JAb/QWJN39YaUn5vcpkoc6eFPczfNICWuHrxNp20ypNVPSDai+
BVGTGi98S5eLfICoLcTqCUucrYrXVRpL+OmLrvbDnW0xSgTpaUvw/c2Iz4n1uNBd
b1r19589KQQ0U/MJRg6UiKx8jYLljYSGom0yLUP09QgE/x5Gu1ljk/Ok0Z5t5wRE
Cqb4gUGIz4RjJmIHRfUU27s1yGikOrZ1ZGohB8jZCKR/g534N28Wa1nP0HBxX3rU
dX8M2qlmRYvSzuPA0VE3i6Z0HhIClOVS1f/4N22rEj7/IszKKCpTCqa1a8iMlEai
DZBaSBRKdJYZnQfNkM839vfGIR1VWUcMtYwmAnDMOUeZlkhsXaqpnkh6U2lbSyYL
L0U4OIKK0CjcD/jo9VdnZLOqbxWvUax7P9s99ovRD+iFE3SXMM3ykUkaeGACHV4O
LhseYRJVdVQLRIH5eYxFyB99ex51jVTkDs1vZZoOtr7sOM/Ua6k40BUqNEYeGFTH
Ydq19pJsIziNGeYqbPxp054Mjb3ovHDc+RglSlEtM/4H+9wajAxYdS58I7VPmpYL
eHxiYqPP29E+oC3gwOvXcjkJiYxK/ShEmSvRrxh7MrMIxku7tQXgJ1L6vJwz8XGS
T8i9x9TWTxkldqxwx8M8Hq/fWF2VYo4RNv9+lSdij/znbTUQJHzZMmjBjJa1DBsy
eQoM/og6OdYdh4pDjZb3JapAFHqpEqG9r8MWK///FhOj9NKA+LxGWZk9k626OlFj
VCnjBFePlg6lfbiTeE9VBZXcp4RyidK20VMkt19t3EevGx5iLCcvba6V5NRwonV8
sdhSWd2Z0dolSMcFEj/tyo0OYe31hJsYRao1lr3aL0y1x06Po02eGA6fCdKVkzDE
5lcicdTsosA3/6rcPLCdf7qzK4bexIx8xSPclgK43/v/gyfomItcNT0jWArFu+zq
mL79dtPT6ZvNngtLKg7FUbmhLkjrCutgD4jnko0gHGQ0hDAc4nyZuBqupyNiSJwX
KzLmgmKf+ZXcw1T8gb2G1aOfcfPhqSjWT8AxxkuvGG+Y1uWdnVR8A61V5j+2Omeo
Md6Iu/RDL9imSv8zkJ4CP+MSTB43KJsi8Op67RFWvqvt/IayWlGecIqgKTiHzRRC
6v0JS/FR1GbPxaywB9BZwoyktKLAN4ULFkt9Uj7Hs0HIBslQME7q9e1dFnr7Sp5W
s5dNxE3gxWvsvhQ5PDn5/dHezSmqMEvdMcirgmmFOfEOzkM7xh1d4JZZc7aE91kp
X35zmEgNTm2mFLcCzI5O0XBwBN99vdUgaJKwX4jivsBxfWT3ze/eWSy9vk0gJJwW
cQ3jyOY224URBDuN5HPxlGaECMT5V0fkCbnEY5O2rTKfaLlWiFj55uvr/zJlt5X5
FELmpfvCZ5r4c6iKMPLFGrLEGAIiu9ZcJu+6pakkHmoifZjOYBP0nHo7LAm31f68
6tHzK9yqgud1f6a42aHtulI++dr4IoFHFpY9mnYgt1Gov1dM/IBU7y/lW/BwWj8I
fNYisOosQXHVpB5gPj3fsV7A0R5uwAd45Qtbtq9++zrTPEPGtzFmzSAT9xiMoi0g
D0h6wK4pvyKCgJiN6Su4lwM0yDKzr5ddI4sMXxR3Ki/Xpu0lkDgx6RICDI+TtnmM
m4Mm9HdolwrOeYpCy8cgq9bVtRIvvYmEoRsPovtz1qmBAA06L4x5teDcFCHruSEP
s+dTMju61q2b2vt0iZ+VYKMmftfAAWMZOLV9HA+KhVzAyKbkQcD5mBLqh+dFqGn8
cAUg1F84VcWEQlTswVH+BdxEtPqGxCH3X1uEw6Iov/nqZqs90vkwKpHS84E/INjo
z0ps7Gg17X50D7iRrCH0hXnRNBwX+x7l/el/tNwMgiwcbCKftnRbliXc4sS1E95Q
/0XAQVCyifH/+dLGGD2qwGdFLmRV4tyvEI9hpLlO5vpNIQxRdmnZJOj2fckBzV1Z
1MSFo+EyBux0oT/60+e0hE1aQV1ZytA5GMGdUtdoaVQk4mFRbLRNXLyiYIgI7yPx
bNV+1KIj7dOhASkZDMzkMPomJsAygfk+ge7YqliEnjcsIdG85dhUHGjFIN/wuyL3
ayILRBcs10Gf5ryHUjLq3XhkfNW6LqpjJZTdXWRbYHuGpgvLnQWmk5v89hOdlzRU
UAGJAFpMmUNuEAedUvkPme3Zl0HKHKHq/H+RpCXG3khcBTupzmsCpe+FFi/vKonQ
eg1oGNldvv5WsXf7wrNaxucAONvpGjX88Bgx7NlL1R3eWliNKKWRiuBgAvpZ8ZPa
Q1mGxT7UnWR5NsBbMnzvGYhA/FYa7uGebveUAZYc7ux2vtN8DhIrhGb1OpTySoCM
C/FbfJod2Tlwkco2Altt6/EvsreAKdUOorFALIliK90bU7hI1G766ZZNL5mvzk4Z
/72SPlb0NDVNBj560fxjnfkO+0P+uHhLThW3Xseyr+2+7pyvYW8RfDfuGLPquoGA
OmC/3cY3WeMJY7FfD172voaKAjcea8PWpnEf4wODljP0T1NbngQ8oxdM74pj5wvz
tvyU7u9pEq2S7pTAs9H1VWvd/KZSzNLbke9jIEXFj2UeSoZXz5VPjlazZ1G4ZusJ
Rc4/2lfnS77HwUMqxaq5Zp1LEGUQDAAEJIS1OECw05Qp1ov5e7VVg2txHNLR3Bui
AOigw4gmzvBG7+A8qBz79gY2yuyle1BAzJVzRx6gLdp+Em6lx2kFACaZJdvW6p+4
/8SQJ1mF1Dl1Bs67yAfIPnrFFMn0oBPCNfDcszayR6lXCTSxe7Uy4eto0lDXiegm
SRZe0C2B048Z6CQgooJICFecKRTwcaN6seuSnXJnbuYtoawhsedGBxNTvcaavtMm
rJ+2lMUaCjSbv2vvU38EIXKEOZK2basBdv0a/IkoJZfUKHVFuR8Okm/4cKWIcszw
cZssmebESmJwBQytSS2GgZDvDvAlUk2Su9m3aJALW8LHradHUTQYjgOtViLXNDyc
I/ute1sziSCYqUsFs4GbKjxKOAe+YTmJLJ84McJDJ8USZtbA8nLE+vesXfeRy4Gi
3wzUjyKXbmCfsQCTpgki+df+DMllAyftzJcdzUjDnqncz8vMt2gizKnDh3QWqtLZ
G7+MMbRbhKYBpUn4+kjB6UgormUYSbEN7agFmOWK6aRe+Fa4oy8tJERy27923pck
bVZ7TEMeP0eDuJlysh+4vr/rwxybMaZtUEnKBTvFPmnd2UWEzAI/SQFp3wy1VjQb
YKjYBxmujKPNXBjQfWszKh2WTsnlSE/ErgOhrdmfo5DcSl/ZnaEbVjT5uW+e1Ta2
uqsNWFGwX3y5WnuPAYLDapZVcdVP6iCMEF0Z3mdqM9R9SLN/e6HRdX39BBo3JbCX
OdswfeYWavS/75Y0ZRJFjnbpf7NlaEkhZsQbbYfzMSsRoKxSKJEjhftbLJ3v5XHO
C/0xkFz9c0OTU6dRhyrFHX5csrfNup+Yq4nf1dq2+GuODG8Kv1tPNtPAf2dijGYI
kEa3PuKHsp5PRavxdgjekGt3waoII6du3I5RLyWtLygLPRoeTrzNHEth0jX8UJEs
hjkXucbIG8kT3v+JECJmq+ARIab/7jm+eIhX2+n/34bggZp+NIS5d1FP/LoZekBH
YqjkOL1Yr+pHGTS/y7EgC4RIDetiItqxb+aMEIiTEVsyg0Jje6CVXTWAQTkDOQOr
T636PmIDcDNS9VNXZHqyGfsdsKn6+j4CTVw6TDoOqQIvs7dcP9Ml8mrppCJTmVPe
BplcoO++5h7/yzBbiUM3wPk2cr05MuW6KSAzLXkVYBEEcCp32IEWys5YVh/2vHU8
PvRTHRhhJhnJGWx07L9TGSrLXElZdqzoJxtEmwuGrYmHpXOODWYrRh/+AfkUmUnl
xV43JE/nvbalZYSYHF9MAWHIWT5hTeZZ0nVuu+jOz63mEvITd1jbgfxKVsY6lCx9
++3U+BeoxaxOZSoT1nppfocb1dE5SJNNiLHxtx9Mdv/PS3Kxd1/RePIcNT5jkvV4
E/DJiYmp4URDAe2qlBGp+jRDllKLsulYMW9lLKvIPnlPf/8pVWP58J9dLtM85JeJ
idS7A3ys1ZaW4v7Q4YmFtWV8WSg7YEYDMSGYeHh5Vrt4O0NI5q2gQ5E6C5+b8fY3
Y8bay3FovwTbn1UKzJRUYlCrzk0SsATSrZ4Mry4UUVgZ5ZRIcBj4jaPZMbD4h6E5
kK4TL3PxqSaYQwzR28lY9dLW9IHzwSEQzmWb5gIWfGw1hv+hnd9KiKlKeTYt/Z37
eoROd8xJpyilWgdYHyY5MaHYC7lyRqpsgfacH2OdKxpnxfLepEbsLfJrlX7lkSrJ
fYOLwLgAbNjX0byJ8JyX8WcthtF+BE2MoY4xSPOCgcuOHfmoip+pPAZm4xryQ3i8
IQw5Ksa8yrT39Wbnz6Lsi3BHosj1C6l5ACR3Z1Gjug2mzTPC1l+3BpQEJ7nqrRIV
X66TG4MXqmRsFDxr9la75d7QYQ4zE0C7fIiddDB8yy1IMtXwfwD+H3Z/inOLE5qu
qy16RyesFXAcffLzTToUvjlXmcjkRvViPw/Swq8IIT4jVmlt2hI9y1Dvo0FlzwMN
EhLXT6w4SXQ/yc0dahf/+vz0RUuRQECVCC8Xj0MemPEa8GFOWvgP5CeCyLGl7RyJ
2aqd4kHSRcgl+EtvaMuMJGnCBGAUDYdiF+8yzZ6PMzcl0Tck0jreS886MqYhfLuI
/kHwbd1aZQoEA16Wx6hSRI8VqURVSdZuxmL9IngNjOr0aWfwn3s+ZGsYjH1e3eTB
+yCIx8dabw8yHKxKEqG1cRLVvOE/Ln3T2D+Ptxgai0SjZI/KobMXEXpXvSef/sii
fGBE0LxFcxYxfFl0DCUqg465H2kLqX0wB9Atp+84APTk1hlR/H1l7S+LigIPn9bA
hTMWmRVdvOZgXNiojIdFxxUNjlrrAkqEGRcamTl3FP3JaRsqAT+zUkAqSl8MCIfU
oHi7xBSMYIYtVR217K9T/7tnFtxvyVZl5jo6MfHvPnJ1zW1WrUXm6b+bgpzUKHw1
Yepk6YsbqTst3kibUexjrXNsEgBY8JwC1hfNTK/0t9HN+W16Oyb64Byhpy2inQfI
zveDlkaQXUwTu/WXNUAW0jD4S1/3tuGrtNOngcru/0anUCHeQq+bAveex+mcu2H9
0KumVsurzkqjySG8axpccYpymSI9tfi+yyBE2uPTi266fP+zauXPAVitv/iLZILg
1QI0nCt2Xd0SLnQojrWLZ4kTATMdSLbO2hmB6ceuBmomtPnzFMMPOz8lFkgzPCja
pyP8zTaZP5o2SDlSXn7jKfjmV4YGMlUyHyVFswIeXU9KBC+exUBTOlt7FRWAZT8C
k88rfv6TbUKKJRbKkYxDU1uJbR4nbmOjijffQNfQN8u7vw6QF3mK+JIWo7nS0ivK
sQM2Fv1l3HjdsBCvfBmVFHo+ETWwU8ODgtRqAg/yTEVepaEP3/htc7uo/kF5Rv1Z
Fpyl0nVJRbf2TEXETA3uhbvelC6744ZmXT2EjfbRmOgzCx81JBN5eE8gT+B/ZEzm
hk/uT3IBglsioYLpqICsh1K0+lECdRMEKP1tpWu643ydP6ZFtnbQ1GFggi2semEJ
+jmdMVqws8LU5sa5ns8P2X3QJYxWFJbTFWjcyUm+FddsGeRjcV6/Pr5zu4oz4p+N
iJ/EQ//ULBmUDhGsvaU8Aa/Oa8TM2R+WszSnh/aGdogDbPl+QacbGFaBvsS7IZ9x
BKJYuSLJjiInftsOSh7TParF561oKMayOaXSw6jeWHrFDWVxrdEv1YLGDz6aEmbr
5XczlNZukJmuw1l/doJF0E02lff3/jUbmZ9xjp42GX0IVqLTw27o1p7cSp4ZOmJ8
KgrP8nJKxtaygcbIl/1oPiB8r/d9qb4+C0PYWfdY5xr7Yonm+97XmQLODW1kRDly
O2/V82AD7a/NxIF0ZIoAaRdt6Dw6SQEW7m4UjlpXRkcUTMS/norsANCn3rs5lbG1
m91nsjZPgls2NWoAa7gWlsm/MMST7fTws1ZrzKGSzF1+3yQFpJRrJOU3BvVnvq5v
b6afxMKTRGdUEqKw1TCNtPt0nZ6TbCVwowZ2e/5MwxsWkSuYAgdxSVh4SZxcwD8U
cV9DXZd1MGTiV7JWZMGhgPNVwo5LBSCZV12eWNEq1KGfEzKCNzqfEnnlQomgQYFf
ANGrKCLCjqlPGfbF108HF0RRrUKEVb6uq2xUHm7eWfy3eFoANmoP+0DvNLFjP/UK
9yDR/kte7kyWJ7xOJnIClC7mj/bzkOnQwROuE7wGFCDo7MmygwZLpQwNfB8DBxNu
YBbvRH2LlaQqVqF6QNyyPidmHQA3KCU3zdKcOb3N8P26oumDvPDVWe+g8K+wFbcq
NgNzUzJfjmQDJfgZrvIjWCJKHE9y4YuezPQSN8osEd1bSmLDHu3zon9NFkKAOApz
7O1nFWiV6/5LF4QAhN9yufO5j1ed38nyLYh7WV4IXDjNryewPZV4AfFhE+IyK4Nd
pTg8pQxxjhUaw4/qB9rKAHF64c0gk0jJQbFM2h0sXSwDHAILwbzPDfOWw6mdUazE
PvKNrKkhTHF4fPcmUoQGQUFEi0tu01LBFH+d/mBn0sZ8iKTw1PxK0FFM+qWTiz2N
2B2jTejxyA5VuiR2h/VJUqSiTIc7LQdgj5DCCNZaHH0UlGb53KEksfsRbTVcteQg
w7foQQtpepcFvhYKGvJtBzIJQXHQppFUQ4wn2YnD9vGBzTkiKIf8AOmj5aqGck3u
EYq1225pqq4DGE9GuHd6m31pV5+mkHDF9KbAe+vbCl16xSH0MyVR6OYu07y1rlfe
meEIehlaC9l5v1SxwCOm+hSTys7c3g/EtyiaT5q5feiUU6M2Niy/8HKtiWdSkSXu
mIiR5dLUHoSG416lxeWNxdMOEICA9A0RksFYsdq9nphB55qfT2WaJkWuKq8sJnLm
cEwjzpkgBtI2g2U35fhe2+0AQqxvqxC+swvqU5gv1v1TSgenGBhleXqpYxu+E8vw
li1+YoI5Vz2Omoi6hLGXt/PpUElwr1cVtOhkvgmlGUjhUGwgJbwcpeEULISNUCfr
wknWWZX8w+RFXSsPst2E7Tp/Xu1V14aU00ZMs77w1jH14end2iU0xIPqcA+BNWks
u6ysjLkMOocLxxMIl1we7pqe+iWG7jV7Wu94RL/xw2wlr8voZ4oqiCFLs1NCJPC9
nzZQN2IdQki9N9s1TMaaoz4IUGgBEfv5b0qWgX6saJjBkjI/8lM+A3qNotkO/abh
L7dnvcleNGNO1zTgAZ9AoLY16UqxTqWoR4dpBI70Tq1vzyVz+tCAQBxKov4xn5WH
eV/pW7ORYSk/qpe5YZ5fexf+LaHx2DKBkFbCFWRnAP45O7EFqnBqRuCjhJNuri2S
kWD6cWMhet2fbMLLkttdLwyzKxvzqRlfsDF75Y0gF171TRQUFjFgRtk2XHHXUoU1
3zug7anOAp5rZIwgR1en+P04FGN5M3ZWaNuwwKh3qKzcdprM1t+5e/FaaznHczSz
+bcRidRd7Dzveo219aQbczkt+AzK9r9cn0w8Clh8AXqPrqHwV6AUS1oaUiKPIG9B
mymjtz4qH88vhqqwPGOmZqdDuG22EOb+qMpqbfGrnu6u48NsigXfH0v42/usUoFE
0cW7257P0UGU1ZHt0KD1wAesuulBjliQ/uymtDFf+g1eRTQTlir83u3z2Ka4ObLm
9EyRZS/zx3M1xHAYvi+Y6NTsEhDO8sh1olliW72iQ7DinNGzmoQSTyfPdMVit0k0
weE5kGMka07WTA4RFsvk4DYR+rWdCukitBE8gPSffHiY/PqLphCNUOpk6/QahZb3
SF0M6OOV5pk9hJztp46n+3pIdNMMdbXy2pGt7D0ePidkbGINma4wtK2RM/fV7wVu
EBg7/gbz5J0C4PYQC+kDhowPulhdijR4OdafiYjbeA39V8BB5ZI78KrBPYy/1Wbm
1vpkcjcGxWU7woCNWb5SFqMVE24wcKw5WOslZdUqS55he2/zoh7yCoYsgcuddU5I
OJgBNqN5s86MYvgXkg1G4UiMFyghYZxRKS+w6+rpBwVTO2kw3rtIG2EnTNeocICO
m+akOGeyHW3dqLoN6Aw0d91fXedlxwKO60jfcE6IwkCZ6wMCaIrM73NDbig77iw1
Z7U2zgE4vsU5ATwnCzoDj2Z0nZt10N9o5FgyF/3PSzwSno4t4V63wAvNuOP1/WV4
5BR1HcI9XhgrsBsefLloM6KSTl+pXEGqfqGHAaI/Bi9vo3Z29fwF+4tmwviYqy2L
xzOtvecYoBDaMYpH3i26XGRLDjw+t7L9MUWTAV3GGGNUE0Wb4m5Kcul97sh6uVdK
6NTbLguGfT4hKLtb0XUXUrXWOQZGGpeX2eHuRFAOzX90cYV+wXrX1Lr0kqGuZS+q
X2U6Oa7XyzBXPdhAYZ1pK/tRfAd+r6CEj50puQmjIvT7hZ603PN+bEvZCySC50Ca
V6609Miwhau3q/GXHPxXTglEzNELpnsDa177MDH+4gEzcyE0vi6lx3gWVMtUkggX
6kE+ceuC9h5tvkNxppb5XfQC3fQ+QjX70Pvxn/prgQGzg+o7ROqyUbc6KRfsoz47
tp7JwecxPr35vIwuMrJdzcFJIMe3biyEHkQKXwImVPzW895JrNRadI+denZpKvzp
mbtWexcx8xm3Y6ul/4CszrZUQnYfumLLNhS/+chpSD3Rzv+bKhGK5A2mfOymC+h+
Q0/b9CNUuK5ItqFH+dQDdbEfxyczESVsFH9RiGWeRLDhrzDbJO1ezzIOUzRBJ7ss
vkh01TML3XoVdTH2Ge2PDsLEOEaUkLmIx+HYSGbgj1qp8PtBfdExHkEejkBdu7G0
c5MJm4/0Yq8pN7zYxczggNI6W1jprYASlfWHRmObdg7aE8g7FjW/fRh9PvML+SyP
NRmoXuS+3esM7iZ2eASJNCnRmHyegIzd0g1CG4niyjfsn06lon+9Ue4LJRBQ83QT
Y8Fv7/xyM0/7X5MSmhsszOH8+U5SxU2y6loA5Tb88aOiEjph4oOFqg5vBG12aEHt
KX/T5Vks0Vqy6tHjc6dK2+ABkg98MuYAtP0drrd0RDRpAOuU0Ga9GaFUPYUgSvNw
X/tzHOeR7n91nkqp5W562pLSYZcumQ85mLjUjn4dUdAfee0xv1NSMN2kSPyOyJnt
tJ4TPsSqvnlbq1mKkPHmgHXizV1cG4Nvh+RgRC7gSnvTaOwnF8G5bWOobz5NVjYd
18H7Xu+FgyA+bHRU3p+ZZzkzGlIwL7uYT1u9IF27+D+7Td5W1Ibr6j+ndNxbRbBY
3Bow3Qk0UYEmT2IySXhSLAizCaD3yKgc+TshMLRF03ygHP3lljtgVEuljvZDS96i
DCoEwlpJL4dO0oqn+FOxzNARNe9TagQDvzD6+z5hoHeYi29tLaDrzWgpW1PTdVpz
AScmrQ9EdO064Xx5hkMMLKORy+yI49nimypUhDxUh/dyM6NMxLTf457hffC1uV4J
DHo2ajy0mK/Hjru0tBmg1wHUqU6USZLaOFtqNHmn6G6D7WF65oGchdXmMlxF50cf
9tBeISNuAbIqVzozkreGudrapJ20xeJ41aQfHpWXv5L/W2Z57lG5Mkupi7ZXvlG3
e4TBknenVMhh6KDFPypGzRtLye35iSyYUty9ZUzEX8+dGXiiVwaHlJte3NBvsitn
EvfgPvdzLp6arizEirLesuUfLZrW/Q6y8Xcf5573I9s5NQIKjHV9rLh5hDMmP+gf
u2kmPEKsPyMJI5rWjDFoeCmX2ukgbQdlZRTlVGFGc54McCSEpQwr2ONFD4Afxnu8
eEi+lFooQvjS//p0QPgpamymhrWmfv27D40bL3xTrxRthNvjMrCy07VPIqsZs+ZQ
HKJ13IPasFXh1hLuhIWtOTrcNQD3LShOx/WoAaFAHM0zX78lg8X8nUBqUrWdBI71
Faw3wuE9hnvPN2ivPS6hFg1X6bI6IDLcpxwhvMfGRN0SUKWa/netpX6gt1unvYdc
q95Icnj4RvFg8j7Emj8ichV6UAbQOlJ4lB+rLNcGx1pmHBJmvoBJ6SIoLEVDEN2C
c+F72/L1fXa4WUjNMgAAm+hrj6b4Ls5GW2Okw++jGU2KkhRr8RuS4E+uPx5R+8f1
Xd4jDE16MbIxZD0Fbr9cdU0H72aHoGWVlN6laMofOUtNOBSRrdZtDQjHfB5Ovf0F
fgOgE9Ygn/ph6Qf3CXq4hgq6Lb2AgAnwzEQ8lojuM8xNpZ2D/lFvkaFKAKRerY42
43/c7ez2vbO5t3XDrGDRWPuGwCmth5oYCr6fuLbPg2/DE6QQ31sUdqe73ha5VE7g
qExpdMBnPM3mS8CHh3FuWOmEXkepi/3617u6tGKXnJPZTANubTYTlwNBqwrl1jQt
k595RmKBfov1P5Q/kysKwQiT16uLm9YBhy+6kKDgRSOFuL+O3eIur70OWHFgU1dX
sZ0hKClEd/uOcwuMRgPV41FGPPzKpq0rvfiNyXhlFFyGyk3MGlOh0yD8POc4tWNV
QXSceLsuO1WyOvEFbtc2SF359IanoKDYUNYb5YBglX8bJrKzv4Pwdl/z/HQi1EoR
pU9uSMxJd2rQOrZEJA/OFTaX2/clhJZPCc7PRdqWD2IrQxEhRvH1UacT8yOep9jV
FdborYEDmoovMXTDaVi/vujwZO7QwguAdgOBmRti4ncDQVfLx7x6iOAzEJz6/jZc
FZBQdGGNfA6F/32ssW28Uk2mt0AvBZfgwZ8ZPxwi/ZhLNsKuksSBmp892efgTIV+
+MaKN0zqkGGjczxw2X2avH1K+fJ6F8qvrVhryzDCv7rAFKqgBq3NwiWo4bG/vXJB
7n/oc8T9IqL2JSX7CmI+T6js/ZT3fyj4ePCH0CogduQ2rdiv7jtKthIT2bN5rfZt
PJB060PLisZQIk5JzXXXM6DNJcbnoCHkwtCVTwWxvdBGAeXIi3MJ8sYw0ivPD3Ki
0yhNmb1qu5lbz1K/mdKH+pFNyVgs/y7znmN7FlNbnk+fhgHXxheaGBHWY8quTH5K
sxyFh/7VJ/7s8eiosQgbOtY+F8oJsiaUBv8RC7hMdl2hrHZm+asHeSh9R2L0Mwb1
P4D4z0oQdMh6gZyj3NwbNMU3zhz1spq5OkiycBATA6kWjzgli5gsHezRno88WnQP
nlfuS/aeUl25P17BxEDKN/OvcESBZQfX26aa7wCiwwwN3UEcP48m0FwVOdqtsOcT
WkThT31r9jhClRtDiFqt9TyVcl0qyydQZ9euC2TkZZVearaGq+qjGVHd72hHBVFQ
FwybdpvEeLB96CHrCGaRnOsx13uXznURZQGYMT3JH0LED931EbttyqHBrB+xNICR
IZv9rFkLm21pfukw19POufCUAjrPl0rx9iOV+7NcJGD7ULXiFL4Aka4giK37SY8p
odmdGJw5+UEMBHBWHMp1LL9ijkeT5QCK1y9Cd31uijlRlLL0mqFQpvVtoFuwBcoM
5P65AirURbqxoBPmIytqOgIEpyFcPuGVRXRLNXnGJvwUVmw3O7RXqgB9IxAT+vZn
ps/kNdO+MMViC22QNncJOKlRvvQb05T6L+j4zpmlI0eIV4SHCFa96A2o0Vk9LJtY
5nSCx2ox8ccHWyhTe1X6a/BeMa5RxvQ/jvXsUHRUbcxA4qXAwNZTbGNyq9zJRqu+
O339tVSjJQpVsgMETPIoWHFwHLh/1o4Vp15xWJqngMZEru7Vv3VEq1hL/9vgb6aK
a0A5ZfJKCaqAW8up4Vgx/3L7pXz5jiPl6BqP/BJahxstlBIoqOtl8kCW1pf50k7V
Z97svNpNHC66yv68QISScZZb8grcOTXaCwDQzTM8og3OnXbJNwerG66CbQCnbmwI
AzOi6H5VMkMAjIlMi8+CMeElsRLXVA9vWFXCNCmGjAa3tP8SheQnUX+mOJhTmYoO
tYdp9AxS1viq2+kyWEKkgY04qvQ6NIVDfr8HrhruwVyu8YzSvxpCdhBk3eQWgg5R
c06vm0PM+ng/8SSeCQozrHJycuXJK2DsMfPtMAv14c8hZxtXyBr6msCe3DZ2rivY
92Je9gCL04za0EMY5GopItE4V+TTi3ls9HzUFYpAMgXrun0owuQifLNQQR7HsD1w
zduwB9mTckXyb1jVzbQ7gXFQZCLZ1RnJ7zylbXQ3u9gDCxangQYu3/dS82vdmLvp
b7YzK4nLOjcEBwLqCaq6z/lE/4Fwlofq3txVEnzT3qWaGRh9CepI2F0WVkxlPkkH
omPPFyrJLsvWzzoWJF1pCHbsybnCOQHyVMi4EKnT0RTNyyY3fgUGFrTx61na96b6
L42qZCQPsJU/rik7A/vJ79hzjBClcNlniaOfG0F2n61t26TcXvLxfjmJLiF7T4zq
2HjsKGjQ2xN9UDy66/dS3Tkrj+oCabb3tY9upPD7NVS3Dh3hx/3CQZ4cV3A5aOf6
BXsfjvzS2eEypsgE32k81pbqqL6LZfOmbTPBGpjVPCJINW5a300m+RDXXIdMYCdi
/2/70JUfb5PB2ium/R7CoYihNE8shgvkKU5lTxrxIn7LxtbvO4Zo27+iVQ1/ZJQX
IcRLRFxCoeN+C4ELidVXX/8YCNK67UYpd5SK/Ofsi6aSnxt6Dpsfgg3sCQ/97IuA
suOyAGfE8AUJhr+P4UtitcySSEWAdjsAiwrZ3f0uS9jxnqA50Qp57uy3TZWdSiGG
UVIlPRdB7o60QGZrLkbnlsLJkqOeUV/SjoVfP/ijsv+EuJBgoxD3Q1Ge0kAU753r
oQUu6KaOHtF2F1lx/rm0ZRCa01MjBrEgrdjWmhLNi52q7GiA8gemaJ2ES95If3oK
cOONT8jQJo5JX6w2IEip0MIxJiwQgkRp0HgR4K92yA5lpoOLFw4d+IhjS5xgeM2x
IK4sFSapLWUtnKU+JkwrP7wSEDIF1l0s7zBR6AtDB8QIFfPBzL7fiRiW6/wfj8mY
1V45k+ISaa5GZn4Va2nv4sthF6OhKOU2AkjdtW8Kp4pSakJv9AlEszJmpEUSDsyR
sCq8PdX62iR3jDmgoad6KtFsoWjKzwe/BF51PUQYi1XMkM6J6VNT66Qgnb/eHkCu
r6URFqoYGwLFmmWXq8h9SMknSir+5eNYyNw33uHVIy53z1SURe/8vsvmCKOxQqLM
gCicnBSaALyVPJH7Z6XkIe+KaDo/ccaHkBwuV71Bh2+uccj1I3j7jbzP0iV7iQdS
ajZE4VDQMc7MnkRY14muPGD+UVo5S8NIUEOrAwJ74Jg4icRRrFBgkKB4eEAVMaMh
pyFm25i7eaY1VjPMOCXydi+8L7UUXyhu8WpFYOdVH31viNzmW24rwr6Usay0MCKk
fbpqXDCuGr5wsxP85u2Imv1gjm8/hqcuZ5UyzZw3pk5Go2rKVheL0USF3JSw8Ino
BTDYWDq7+Eww6TaJoCYdpU1yELmDdQJQmKQ02H1FY9vauXD3GuDluTy+KYx34CHa
LFUzi6xqknnWe+PU25OnR8R+bumXIKBVamtnlrNWR/AYpYkYLUtAX2xRV3lYfKv1
75e9XQzSngQTbyMtU3ig1zvvPosXcCwzzvU4wGdbV9q8zv39iC2NkFz78iB96nyJ
rlUYOXjEuMIbM7q6yQcNY8LGsNG8Odb0gTUL4PjVv2ohrZWQK1nivMzESvZ0Jjqp
j5+li1LYbNhjlrIbX2ue76S86WHMgx5lBKHiniXwljgtK+akmEwQUbcPEUAYTxph
UtvNvS5unsjJ4uZ8rpmh7qx6yf3YU9PjuR2fZKIrsIiCFXh0RZYhUOURjmCjum2K
7soVDFRZQQGCH7cgzMEOaZqu+U5dlHPMLvDyVBzmjlCHb4LW2LXe8agN9AbBlNJK
XWSu26LWQXnL9FSpCFIN1+jXJM1BssU6148NJLHCOYLXzJgMydy4D1GFYm3DoSI2
3Cadxq8mOGE8MRaxsPHVs2L/aCQAnYclQMzjyFbWnX/Un6H+smXOqN9l4wELm7bV
ZM5tY8DBGth8Lq6hRwfyWsmzfYfviH4iSPBzZ1CsK0sTSApBSbTOXQo1O9s4+ALL
kOB9Xo349nYH4QtuBESMyJnXcejTDk1wlviy7TLLOG7fS8pJh1VF3DEE8l/W6RXV
1ij8XLt24XtTYGQpn82MRDytQdKKD+Xkva2mgSuCYKKP6RlDoXP3bnhgt9A1UAwz
b+G4mpJaZhv76KtwYryzj2N1dg1ODr+pp9heE1AOFvikLCHm2sFxgU/IWIfmX6gX
D6+4asC2jU3yzl6GnLIMFE9Ys+Wu4x6On1gH+bzMW8sMvh11SdXW5qfonwgCHrNW
FGTKxYJ5pecgME4tGKbXBybHjY7FBKS4zXakZQ1NY5/lkt9/5xJ55yUxO7KDtz9w
Sdfd2MR8/gEe5c462FtLA5VeVguMKF0NrOQa7vM+jWJmX6y2uVv2soGgvVHHm/h7
aBUtghthazHk+ir0G02nc7b0wITwjDxp4dLGg1a7yx0GwEtApPmJwWbixadcc4KB
t3r5NBUy1OM+tBzLlPgkqyuYYHDQZu3mj84e1MOGK83BVNBFb49sB7ubvSkUiWTg
rMV837OsLPIDlMKCY1ngLUmMs7OCdvTSoH0XrTedymqssbntv9c5W9uLcmhUTaQ+
N6KtmeavMTo2vtX3YgfYxsdCgFRVTmijQlcQGC8hxra5pUgb8jFwa5qTRAgEhFrK
e3XCnk5H0LBb8h2X3DDv2MT5dMTZNhiuCbuCpjYtnU43BkzGMrwNPOTlbkWj8mgK
oQHldc9hYo/EWXqfJbX4R1WvBoc0QroJK/tuX1QJU0DrnfjKuf9YEWQC8xro3P/s
aRn/aOsIPcRjRNV4BE2b2GZ64NVmzukY+3FPm7WiD6o9rsw5hGokaaN9M738OQfM
xUdXuUWwcc0umorQtlcwK4KZfKwMhoz2veITCeOnNCpHL5IzMumC1UDPJmOju5GJ
A/KnxE37Lv+d6KKPMmwfmuTJczCgIBAQfxkegfcQ1e3ott8BsLSi6WWdIwO+drvQ
0YDM9uMB+o4KB5/z7+OVd9eNcpwGdU9dUdhr+xm/H/qzbc/fymhxYW5748vHwvtE
JVX0aGxbYqUjcL1TvUkgk1QXyq4hLSiDzM5dSoJiAnfZSl7PrvXoowXxr2FDwnrT
aAL3iP0yyNcn7QbCHfjWeEOkDk+YPMNLEiVkXpuKmhGkh5aLKJ1RP0nSzAqmJ7+8
7Xx5c1f5rIYpL2ZafgyVidZOj3IWPcqZGmE3YnI3MsaRLlOlMTJLHeBQUjYnSVgb
xSFEy4ISpHUJtM703NvBUtxHdHm2hVaUgZYldCIZqIAz9t5MR27Tb45X7yjR4r+a
w+MPrdHKn/3nlWe032JcsFsuuAWXfVfqhxDWsNt+phTpZ06j1EcOjzFH7+ZeiSef
J0Mo5sHKXpdmK6lSvBKb8aSiM6eIMOi8kcIe5Q1VhdWCdQG/R3RCGQnngi1PQxYu
U9uR4wUd5Qjy068qmJqexU3mhaCnJKphuiAbeqx0sXxxXY+dvpmdM6VdAjKqRVst
8i9FHZ69RWAVeSJXRJwNLeXVcxuBmixC3VizShjPuxnfobyn5n/gYkHySyKlWdwn
rscYIE+qvwDEAs93xl1vSZq3Ed+QSNq4CoICIA9Jp9270g6QB7AY+DPDw1S0UrHB
TDQekP76sYhgowrhlji7i/NofeM0I65ZIip99bpjeuaBW9zqRvRYL8da+a3o/L0F
eIvbpq6C3FF0PQNcSFvBemea29rq/zpoAKL9BZU7JfhwukAGB2i6iaFonX8XNGqe
mWAJY2ZpNiE8n3vvnkwvYJdkuf4vfCzh9qHJqdiLqdmySBTYfeMJ2twplSUAW4Q2
uKv7J87ttcAWNR7XxPQg1WXXNU310hbiq97ouR0RmsI1r9STZvmRdkH7hCMF8AQk
Q7CO7/V3UoowDCowIL/HfzwJpvMIBwMtXkAek3cOcHLCzMuhWmRYPnDJqdPjZKRI
Wkfl6K68QojTdEYwD6b+HyRpm2WkbEumWN4HXfqkhUiy6aVL2Ov5Oa1TEmJGnFWH
7VFbiMLHqk5Oy3n/5sm/tbhv+k6i36orl2oNPgwwOv+8hm3SVlIis3Ba5Mtjkftr
9DvXnRCIFLT03s3bF5p6k6FLoaAdmAKuX7wjXtYIJ9ymTsD835V16UceXEBHlU3z
rZoeCpt6AX2P1yg+8r+RGHpJEFPkNYwSYsuyVFw7GgHeVFbn6y5UNfiEhk9qycHu
sCI/60FnK7VmIlryFU3K1hG9nUT3FVEmtnl+gQAo+OR6B0gNGBWOKivkfnpzAmVW
JzVP5RifeN24krK9sov4UVYEyBDjTjOzHAao4XgpB7+FcbayOAJwFVnOiKDrdbEH
F8gFAjB/kU+WahoMK2mZMbaOeS7c6BJjlgUFwvObPlkr8vjR5kFtgJlDWeSpQFEW
wrRL/Or7wK2spMR2JW07qkih5TwPbdQwE0PI/qDFLUmgENUYF7VZNvl8W/YwykMW
Qawigs3YTm78UwYJOrZRDWYbgGF5SVH11CsoohL610bFC9bio58FLOL6sdFhJK9U
0sil0VH0FPk4KE/V1/iInFlubJoSJ+r6O+q4vSFnaNMwASzaw7CADORdYYyKKvIA
aOJK9s8Plb9oJV4F0XqctPuDuOqlHkT6uL77+CTsPkdg6vNXFzM790cod06NC2Gg
pIqxv80cAsDavyY5mHw5w4Ks0hfsfqj6aXahZpwqejxTMtTIUsqE1tMIevje+480
Dr+vUAGJaF1ttKt8GYE4OR4CxCKMsARupcHUFJTljFVP56hL45qb7Bis1xBi9DS9
rQeSKy1yhL+TqklEKZLq8WafmvuNZoERlblr9/MrQu1qz+cWmbx8vj/KJJdRURMg
SryPx2QgBgRnBFD37Fv3thAZMEUmD74KW580uaAl82E5jS4BHti7zE0w2x/GdP9z
VVFktwlI/yxucvvQ4GFdrWAdZITBgPItQZ8HUwNxohsJlbrlD/Eo/+OZ4bGfHC9f
kfSgUTWAIeU9soKx2Rcyp6Yog89usqnf6HTT/0PCJTZ7Ai6oFR14uz/2kcMlXgLb
W8H++Ejxlw2l15VLIjHiV7qTcUSX02h6xOQgoxFd9LI+8qw0GutpYsAcZZw+VkNq
ANUy9BZETi7C3XnR+6FRvB3dMgZCypBEjtEBT0j5GI2m2ZKDiJ9EULdXTBAAXwSh
pzmX7LjmGEmJ3VTRWOd7cCyHsfa2hPWIif9cKzcBPvKpdxTJqjTS6ZISz/UEuCoo
dluwzZ4IjJwMjSCOwOeLWWvlY2O+te4dK8fdYUjoSfisvQp4oXftFljsIG1wgH0R
+nWgBJld1d9UD/Bf0ze8+uNB7I0f7k2i0vLhED7rMDS89BMyOKtisMMV+wZNbzhs
Oj4TphrD4S8DWfMDY9gVhrnIPUlNEcUcmPaQWuSI9jzZuF/adY7h0Z8j1RiLCdw8
BHzFebE2EuDNUgBmcseq8xdSyo5Doa1DD6WkLOgANer2qkmyOAxMT6y3t7v+kDXw
yRXy9ZU9g5RHabT2stzoUtl8jZZTClkNisRROkyWltUWsmD50l5ORsBc3aQ70GBK
aMLmh19j3H1z347pyL5gRStLU8ecsH+78z5W/F8iYhYNDfyrPMVeeFlqDR3WzUt/
E00HneqCphzdouUz9DKL5qJehtmNBDPNEQZaDyBaaFvzWzqML5EkHdEdPsnCx0DH
ikCJ4uMN0qxUIA4cZ0C6hZ7xGaGhh0Oay6vsm8VaXsBv7uI3gOpJzjqe/qjlg0yH
ksLaWeks95/hfcLcChzbaW0nXkZjPU5mhPx/TY5yDolzJydRyja5DLX2znlC70QW
199l+lU+d4hti4OFNpBPRSGviLwFEDMA/6PGaPV1R82UwG9TDn1bNPaZgpnn67Fj
F4PN4iW2iDimuMcd+CqWCa0DF+uRTHK1pphW0wSiJmiN6sUVeBRsXo4csS/ADI6u
XaKh0PdZKosisjLKzPUu7o4dt1ww55MbD7I2wmfz+CANjenZRPM26tVTO/UM3UD5
cmpUjjGzgW9860kcA4pFmIdLACV8k4kBfGsjWEOI7fKn0kbNQFYQOwiZiG7XYGZO
8fiLLm0RIkiobcXoAVgxz6bO2pnFYCLpk32xDvT16llqF9xSdX6w6Mbv1gAb2yrx
cqbGmOMOHM5QdkVrX6l6hrEpo0O2+W4/BOrNDLsydUXJC9h40EYF5lrwNBmnM9Ax
1c5GBf9oM85kQkS2IFcNSXVO4aWXmatnDVMrqnj9Tqx0O265NqA6dtnObyqV9LJz
6v1L2wy/LvzO2WZt1DUTkb8kaRIektjiGJBbA8OCI8L0recKxH5tWHRgjGBFcoSj
l7Mm00xZiVQ/sSuT8wZqL2WqmO5lUW31RrvoV2EIZWOsa//jp+u2nFKWzNFf1sCp
qn4NaGNcZ/f/aRVglMCl0AjmkTyJSg2wvpePzQdceV5mDCNyGLhRi+z15R/ghD8l
7wnGLEAU340sDKxSsWIy3LLH2jkOFm3rw2uansC5OEATCPqZaCW+pvu6Sz0IXyqh
fgaAzTBI8RwoxPbvjW6SYc+Q6iIlsbcl3c0GBktOKTkjPan45Y5/12fAlec2Zl8a
ZSbb+P1RcEH3/sQUYu/jcBSc9julReySgDzfQe5R5ytSWwZ0Pskv+o526Xi7KR1Y
iFJN65dJM0Eh3EhornLUBmjA+POQn67S9iW8Jb//b84ZQIh8WX3hzgRVhMweIFSN
fUkkt/Y+BP/Y3P5ThA136maIUu5GerqqGr64pdq0fgp8H48z2c11SGSyneq0dW3d
/MorNwBKLifCH6mLyjvFEyyXyXOLq1a1eR1Zcv1BndvxTYmKkn5u1YBy6op/a9am
NGB01q9y4LGAWmwM3CB85aKA3SdhLqRj5bP/JntKDt4IYd7uxctTSPBLJke7VCPG
+4ZkgV9rbw8WCqKx2916xhIAN9E1XYg+F74G0Lc3/ZB0SGJZEgJppHg7rRfH1cWe
Lk4gdqf9qpQn5kN1G9Ht/HLf+JAzhvmbp1TBmBne55rZOFoOvfB8/8ZO5ewG+oEy
Ns72cdWbGMsiLBwnnzUBeAaakVhjDKaU0znU+PQ+Yy21YM8ctc8YB7pfqYZpJGki
hg2p4dTMoo6n0TmllTbjwz9lWtoxmYFnfPqscDbeqqqapl+OJx+6IyDRdoMKeaAJ
FYCM4pK9X9LORqWmfAhgVIK3zW9v7cBWwuDzLsr6AgQj/DjojIbUt+bxdvSK6UNs
5l/F+1gMbK+zuxdV410XL+FKC36jxzCvZZH1PNlj/nBsT4MGjLrI11z+0FFxeyyF
8m4xd1tfY9VOwBPdOlWExSMkN7LT4iBkOVSQnBHVjQHPu43RIeM5T8WN+1yzN94o
JSab+TbxGJcnzuJRb+7Hjs86l3eQFjHN0YQ4uQnhkHetEflU9Jh8jaS2nqJ9UfAV
nsU7bN9XiMOvWxBL8OxxqfbCxmK9O9Y4PM+9vZEoarrxTQMk0ynF26ljEsAM5kP+
qWTq6imeeZhU3N4OdTSQWG1HsQDKtZ+6w/gkDFr/ba8Yr+USd1skY+/BLZ1n0aFS
6QrnSmDZU5mkJ8VzeD2ugn8My/wWInf3+mR8TAWJrBVty2y0gbG6jzlocGMfDiUK
B3USIw7SeCd+BYavc1psjsZXQxQ+stWUUBvCsTI184qP94jZiZtR8nXnnCYWrQhe
Wg8ygQJRKsCwAHRhF+mwp8eu0Ly8MCUaHv/uWilO01aXAdkDhyM8OwVHXHEA298N
HXlQJV1k/2DLu4PWSuvZl95l7RJ5TKV8JehXyWbk6ho1LJYiW7+/m/cFzRt1ezIJ
yibfudkJc95YOooanXMPIUDjKhpTFasRrF2KKK8hWd4zh8yTLSMZN996RK75Zlbk
FMKJhPJRE5bfuFIdSMTI3ny51dKPgk0C9YQk9ZvX/L+tG1dCR6Pb49ZCcDwSR5pu
2mSQjwO5YATzBeia28dcq4W8lWqmm3nTdhb2eK2cI837CttC9VTY0ERsgNASLoDf
P1P2Hle6pLR2iD/GYPeQCt5I+F2yiwZpobn48M1E4E56UR0qACXBZb2np0LYkjdv
h9IDcORs1gyYzsC+VqikiESaAqNcMbgIujoWVR9EUN6OOUfpL2j9qJrz1ung+De8
JeYFNHrfC599OVI9LmVle3kd38V47Z/VD1Gfy2ZUeeUsPviTpkEB90dyFh4zVEZ/
A493A6RsiSGf0VsqyjBuROXPlbjsTsrHjX88cwqYGm1MZt+i2sd3E1vrmgn41ysR
Zgg1T5gA0qFU07e8lg9IHpwuiT3pfIzppJkMQx/THJpO6MeBSqrn/mxLaYi0YY8z
fVyjFk27UugWrvhM+LJ6u+17UE8ZsrsKlvEKrljOMuR4Q/7ge0yLNvQyA27T7U5v
7CYrzCvl47WHtCyOa4U87QRS3M5PpBiuuH0V1+Py+ZLg7hMGRBWoQ5VZxShpnjCZ
oc/KA9rsQYFMpFde+5C6x+WJxGAeirl7+pKfCUNNiW0drkpADz/RZd6aNFcTwHez
YNrXqQqVMIBV7NzIV/cuUce6yr71Jgr2/aT/9oEWyf/+ITgLg1CqsM+6/VP8au3O
Kjas3U/CTIYzZWKx8t8F2IXjcqtT51EuWU6jvQCzOD9y33H9zj2wBvTuVW5f7dJx
qbfNF9sCEHAPC+5l0hwEQ8kCAhaS/RyGk4ExlkhjkHOTUT7ay51Aisk2PhGsc+g/
TGJ2+ksfxAgQfNlDr+BCY+Q42bZd9QZbbpEq+zno6F4x72Tp023OfPJN99IesMAA
lN3PoJtFf+DacT6BJPXZvH6ybI3nE/p4T5nCh3HrxS6bmoH2UwT9LmTmOZLbTWCu
mhALmob/Ka7tHh/VO10Pv9f54+eKRMOwg+nSRdMPdJ7ghpgFOSlWiGAlgCzFRjhz
Dk66qrXoVWkBMdFtXe1K/BR/ggYUjQm6N0USXxG9+NW6IDY3AU6r0jX448J94hxu
wokOWxE8i7VjRlug1DRir9NwA7SI0l0n+GcKBFfCxx4GNvAfjLLrCZnZfoUHdOVz
2+V8a/kNV2GMv+jjHUYX6pIDJpPLGBtJnAb+/On3MRiKMB9RzbZqPydb9IEgBdxY
eeAxjvDDz8LoMNCwSsRMvDo3uRLN2gLrBhoUqqi9HCnGOXZI05n1ykKwZrMUDcvk
BRWLwB0grAxoWrKE7R5I79PpkEWi9p/CvrbaoilEchcpqz7eYTZJaLnWznYaTW1H
MUCB30Xz6NC6TV0ys6GFHP1Qxj4v78MCi85KUc2jFbv3w9pNQ1m9scbdrsuBZTUe
8f2ebXJ+Ij/F2apZB0JqLZbhoEVzDZ5mdMkHdpgA61zHxzsOZSo6hAgxrF+9All4
zWnWXUmJpLHseEo9LsVC3kg6z/dVnqwTeI1WSvPlU6AOtw5cRqMmMR2CABrP7bpj
M52XDJOyTR5dCJKQCxZs4QGbJmrFy23N9V1uNjZvJwyGuVbcsUFPDBa47nvtnsnR
hoVzBa/lVSm+eS8O4fKZUO6CnsRw1zUQxWKjhqEY5uoGHyKjRXNAxcJN8NfFN+ey
wUIEQ0qrO7BjQmJNiikJnxS0Shbl7JhHQRytCZf2Lr6aM9CVcpjcIQ/p52hROh6h
5hV/QwnLj7LGGeoPmz5hLcsgCbPFk9Sh17Eq+01daimLSZeQWa4Mi2csHjEttQ8S
F4/je8b87Fjg34gf9BrFgtIYSJydhzth3SHrLbpe3r5gAWf3ku9ZlW1eoKSZULc2
0Z9KqMdRvZWnCr+FRqQUlLtMO85qdzqEJp03RzYUXFdnhsaCIO2eQpzfK0+Me8kB
kxwkBGhk/CLCL3PPxivSMxpNUSMI41Tv8C8fUQZSTjURphx9SvKFRSnvqZ3SLbfH
jf3/y3uERKyHT7T3njOqp5ek/LI+43aP/pPdrqJwqVG2Bqfyhcb5ApM/jjAAZAB0
6/9UW5MEP7dUGADeV40iydyOU3qBd/046yUremqEib4D3zWh2eu895rNcXxY/qxy
OTYJ/nbYGJGopl9HBWhrfJWjFn3N/Z+unYUQUG3YKPK8ysKt7dH/YIjIB+ka80GX
J1ShP6q4vWhxrpt7jdyPnZOBj9hGlKNTt5GgSo2ah7Cyz6/T+MdeRTSqYoOE+l5t
DgOZ3CprQHLR2P/NKqX/5qLJmpZK5KTzhK0j/atIasXe0w9T2VHUzsChcS1S/89L
6tgeYokrdDgYtSmQawZqEupyhqdr1muKO79Grom7ws6tiVqGCLR2foRpEZoKgalf
3wKEYciRPoUZUpQuaf+0Rm6srfLk2nscmvdlCUlpyxKfMMNw/Qn88gBou7G1UzNm
Ojg9FfmfrapqRiona2kYrpCZJc1V79vtLwh8NSRx97IllbuZ7psReLsKDkoWdMRz
0Wgsuh+gtWdu3V8iAuIte3RZlBmuitHKJ9+XyqxotgDyc51v1JG0J9irzw2lgNxT
dPbi6BYkTO9jnbmvZY9aOGdGSAByh2nKMdBSSosU02KtxVBIs7t7SuqCwbWqqH3V
qt2mVtWH/AJUNB0hYIvqceIPQpOP++mQSAf2NGI5KmVAHldVPVx3M7KnVuqI2rsr
R5orbi7jS53O/wlpEKmJFggmOn4HY3EmEZJFOnh/EGXhKJXh+MbAcqrhplJj0iyk
+B5WSYbo8JXMrvQOBqm7RxR2qNscRlKUBd5IGwcuzjjNT98JjsVDRhHQAcQUJpRB
Jvskicl2PpFHkXtkRDR75iBNHsfYRqL5dI6Vh9UtAN+ofvVEbYDFkXudQ8Sox+6L
jRRu7G3bgevFV8fC/4lXFlGc4RCSV4mydfOiG/8hplxAvMkPdfv4Wo0jr+YVvXDc
vGK2prl7oNSS7+UlHwiLeq7hMdBSsNyUgy0QsEHTdiV2BzdJ5HNm2Th1zf4I2njQ
Wap+BRrjonu73rKG4O4GA4QyzujJ9VYtBY+cnJGcLiAAre5l+Ar1+Shr3HgC6pMh
pWGKzw/Gh8H288+5hD7YzU4pzjvpoybnrm6mhUz319CASvHlt5gqXq4aM9vsa8fG
+T+xBZbXqfuOzllWALc9G5I96bZScM+fZGSrMjvNxcqoLTyaI62OWmzM3IZzBE2U
wlZKEyNZPcFRl1yxg+nC9l8EAbrzCuFzzCn3be+s3Qdy/cAHsZJQZpCoB41ic9lU
wpQ4NUv9H/9/NrR809tHQSDi4PtnDWixY8yDcXMUPW+LTPfWfBo8ZZStSNSqvyAl
Q2zo+Z/f44HFq9+HYnc7JBPmh/cIPsR+zVAGqtEopwtuoFTbOc2G88ew86XfDR9w
v6oZpbRBnTDRCQQ5nD83lrkWRtjw8MZY6Z4cosZmZnoHDcWY8VLqVp5uoMo6uA5Q
BsxwQtrN0t2hFEn7b2tEhBCG7l2ajH26rUNYuJrp2FH5/02yWqzpgmuL+dxIM+UA
NqMEwFGKwMP6584vVb1NC5jI47dU9roI+hSCPKw6Tel63PbdSiXbJgizw88Syc9k
cvztIgS1/dxMoQhJCTFVhLNRiqEOGqIcdE36Lf0SoJ2v4MEsU+S2galEXGM3L5Y3
LjSI5lqhGIh5eOHU2NNe7fzJQsOpn9IqB0yDhTrB8HUDy05PPVi6bUFMQd7pZDD7
z+M/qIMVnhSxsCGt4ZZdY7IbTwh8IUQrtsVCLlJGjuLMfn0y6eCrA+0amjYNOctk
KebZ3epfPXbZZTNQ4kiTrxt0O0IVmEO/fnqXk2bOJMz51Zsi4A2SEubU33IaEmsq
wtKLMwMLN1Od5sHXMJ5KcRLOV+0wi1wRAOqKjHHB9lLFrspkdphXWd7moV3bNylq
Cs/8dZEH2v1OzGTwPQhRspzOnejOu0zf7z0QvEDpvVgr7fTvehblFAxeEVYLPF3n
nD6JHFy8dhad1D5ne/mPSMRZ5vGuufaAEVJXo0tt0DzgdhwlXDwY6MZV4Z+pL+bL
piTiPDDJS6cleF2iyaheYDNf8dpV2g5TKbCs+YFcwhEkkgFJKI64emas1v5RUdBy
mqm9GIGuPscwJDyY6ZvX+gGDCkmFM62M5I6GKKEFaI4BaGjtQ0tfo7te1xx5LwqG
jfyNbLpEJ9zHe40MqulyREKVM+0034T+R8OBj3fqwUZeWgnCDh0zlBlebm8m3ghO
tRsUhZvyvgogTgTNGkXdD78nUnY0CCnbYBWMLD59yhqv3Ol10yAGBfK8cMwPKFrh
HyqfGBQRVpZWqtbJIsKEsf43I8ZC9PYRMfPCe58j8F4BcbbwNSZwu+mtlxJT0ORi
p6OtBtgaG3pTCfj0Rxl/942OG8oUcSctGvh9NYivsVjCZ7aIm4QpdxpdJCLY/43w
obvxPvtz0lC/m1c/pGxdbRcTklqC7dfJJVsHO8MZhGcnzQo1MA//5WS4zVjBu9/O
4JTNviq1AgugrDk8d1vQMoEBY2/wSfLUUbrl68z2MVLfgU14r2tWT85GKRKrKnEi
9nSrKZH1ukHKYsCFGYW96ZXkjHpS37ur8rZl5qfn+1xh1uq7cxMUtPMQapeQHC6l
8TYwk+dza+QBmXfwqZxZBvVu3IPUg06ukIjJsNToS4Lo6Zob3s1EGo0BWFQ6J9Ns
fPytNo+AdzHhw9rubeFdXSjEJXwwVzXOfDdSCP9ggnJgz2fT67cmXdOk/Z0hzAlz
f+OGZLWeXXlYlsiw9amYktAtzsMP1OgIasHfe/Ndqpt6h8oR5WDkwpzhCbJfhG/N
TKPkc+kyU6pHcxRQnSsBdymslx4u8khHG5RjCjk1pqJj8uRryY8mB8oqgUN8q04H
0v780RE6z1v+6p1bBILU/vd0dnkHAt7hnP7PEjQ+vSOf9Vb9fjjbnGHyrzWXjZna
muPMfKWJ4WARKRBo2jYdZkENb7JuDxMZJBpohoL0Ltv7uZaV3arKVmXd5DfJkAgj
mjxvqLCglluatvXyIUPXOH7SRYJ12CTMlFzA07AC8nNPg6XRvvL3k8p1orDTFdmu
cAST5fhPpU/ZuWwe7MR/wI3ozqZYEEfheOin7TuC68LI7AVO1XBddbNbws6XxvRa
op65rvJJkERCQvMGYxtBPiN7zZtci7bgEljUJmQpnAJRUez3pql4b0p/zGDqS9GK
bkQkysdbV/25GO6oDJ8OfvHNjPWukGdqC017KspqwZKeTyxMzc2v1Y1T/wsd1t5W
NX6/BM6qul+mq6RIbixouyyzdYzNY6pW5L40vK3WEGbEpBV/jWSCUdN/ZQSqLBBC
okwH9B9ElatUanxUoy3Le/vPOEbwXTtJe+HZ9QxvvM3E1/h/VLLrPUa2PFXepFer
52xYg97t+EhzDoiSEdzFZHE6kav60pDxWlFHCt2IEc8cdmkf3WSr0pPsz8MMYbBY
jAV0ygJCzBbRHO5lQinR8vM6orzrhKZwIM8/yVVhKAq4WJBAIpyZ2qf3xytQfk1c
ois0EUgzO2ndKvAIYb3dINI2AO8t7KSPsFDGOyAmFS8Y9U1/22YWkb//E8/MTPDC
Aa9vUpWh2BZ06qEi1XGbUlz/vVdAwKppamBy0r63yep5tHQGzrXpT6cFfMXpPfAx
qV9/S8GGXmlTKrHzFJE0ib8e/7hybirIM5fR3T0Ia9q+o5kAiT7z/w14k8MjLuje
JKgsX+BdHbkHk/UFMtRiU/28SOqxN4+CvLENQpv3KocfW2gnDxAYObgHR+loNoG4
tvozMYbcWf5cHS6f9dnEC2JUidgcyjfszhdsSVsTccWJvZhwL0rJmaD9fJ695Aqa
MQXZ1KWh4nDz45QlkTpqzl3d8Ag5lxmZ5VL0T+jTMRtDK5y/RJPD3sKv7V82jJsT
4UnNdPBJrgDuysuZBbY5YoYtUaVq4oxnFdhg9gJJTDxbacgK8p8pg/Q9iSB4RbZh
ma0R5Ngn+cY9IsNNGy5UG7dJN+QnZ7M1tdcwaQLp4cnXP80RGXCjP7cWI9WJtQzo
8w41R5IUiQjpdLfdmRIogsi7ZITGeafOsImCZqtsyPcaotV9Bx737CmdjCYu6GZb
IxD3DRApI3kgLvNVCv7txuZX7eAzl2D08UBDEDO2PK+IhAx8fzznvc+3Rnnvu93T
nkPR+eMrNAnzUBhO8783D3XXsoq+l7CKT3YoAuza8PuhpSZ4twm/b9IPCX8Aa8KS
dkFJkkhPvrp1Z623z9nDRoWWfQvIetXHRZLRiPED6lM+k177svKCc/93Komxmu3A
l+aIFFxHgSdiAensgMHRd8c/1atvUQn3+BYsvZfusjFrXLoEUyi69Mz3lAE8OPbN
SAIupwfIAAa1hPOTxq8DDlpWmxKJzMsKPmmw0X6+8B054ey9FOKGfv/t7qQJhdpW
RP+/1XwIQhIh3Gd6fvvq3daZufdgxa977WX0JaS2HBSCUTd0qOOKg4uQf47RY7Bj
8wMNFVftNpFjFtheD3+83Gk9XB00u/NcPmXOvbyctzkVQMdGeAot0b1AuobDFcwK
VR/8N2a3JoU0JvXQRtn3DQf8TyZ4ivpDFPitV8cf76y0BAhUKzJmaubwmgnzD5E0
2PMGJ2s40tIv5o0vzN7b2Ula3jEKmgYhFIlk4ClLmL2HwWcBpj4aH3s+bVTcdET3
ekk77a5su7x4+T/205Plq176TB1wRkc0SsWnYRvoxfCHwte5/l2Eqg5rciAn+2CG
mKMy5K1xETrQYA4pJGUsDxcDFMIYHwl3w2hNlXxkfvbUr5zdfKVqEWf46bytXQdc
FYB0dMjyIy/eDY1Snwdrf9AMEFpggng87BacEHuLAyi057ctW1RVun6wtyPQe8K6
X/GXLiTX4k6mQFLAZVeqvuZ4vGQt/0A20gM+28im7901ooeDezQlJsusSUheffXg
bBOaYtqGz9aURxAj2Czj71fWXjwIFghO2hfhSGN9D7tIvJ4Mdr0FIUIcLdezCShS
6zOTcNWcV1u35ndPDGjWhVNlLnJ7TQmhm9Llyt304S+sxd2002TXpOZfiLfkBmzZ
To+cj/V72h6gLnH3e9WHjp8lLMPfA/7XjRV/BmOmbjKZOeS7Ua/YZkNMjHGGIY8j
MXcM7xbUT1mRQPd5GeQQ0amkQXFdktZdVAJi0H8z0kOdkGHa1kKZ2eRAUalKMzRV
klShBytzz/gAgccZyiADrK/eQoq3YX1qWU/CFBwu6tcUPC5vkaeeAPkelmjFVM8a
LIvcTQm5yaQxC/MNQueT7UcPDMR377nfcfCCvazx3N93eDkSIZfL/11y00Lcf05F
Ta98bR5hV95xS7l8NCPTOYIKpi3MJP6aY0wqYQUiJQ56reFuJTjmRbnDYcdqDxV7
vWSZtI1HeITMXlr0U/yKE9tnm7jzn+xHKAnLf538AO16X0Y7l6mP36ZGXfnXWETI
BPAsx/pRUBOo1q7jRhfH3wJa4ffIEEM3NFSqseq6AV3jUS4Yzq2gll+W//t9GRsQ
j/O+UIg6hlDYetc9brw2Rx/b/ViFI6nV8JXbYfqaFne7CVmMVuJ9goHjXBozkZJW
IY/Z4F8b1IbkrUUmi7ctsu5NAZkAmaFRIZMhDyjWVXHF8P0DIuy9JvuYX4va7NXS
gVgGwuhaXyw8nhwX4RKUSRwUI5mAb4WBWCDMipNsgolIGDLpnRXxzIp1lV89KYee
7k1H86hBcI161vtQHgLYnrt7ygj86cRiFKfxT1BzAbiUKz78DXjgGaIOj35+L+jG
5ZASe0SnYhey7SyzZYhz/bANXs3sFDyTfN4I+0GiFUvfXx8Vdc6w1P+2KGO2O03C
m+hf8lMJzTb4iYIxLLxHs9VZxy75WtHqJ2pWvJWspVaHdZkscH5LvXhgy04UTVYA
8ZXrZ/wPlZOfpwhKofarLUKjPBl5JppvFhKVr7XzpoDJD6EIVHmE8MQiA7oEE0Hy
k3Xw/OE620T2NripUnmPt3iPOwKjC8/gGGlbVDOH7VRqUMSq+QzKJtoPFBfWCOjW
zTGQBKLUtQqfbUSzoNFjAT6/ugtaklAEDpRbGnTp0xzE5buiqjgjdcw0ULmIkNgx
C7n7TMg5sCejFe+M3nu1/5OCnA8X4zSrfhyOUk+NFLP3nmr32gurqntWIBzT/7lG
/ZmKQX695hxCATIjpP1FjVP4uoDn4khzu34bT4/ATfgKyxJNYKi9s+VTNweoKOMA
GqLtrtf1zUkyblC/E/KVqrEpbfik24M6pew335utpQ8nojSM9+FklxuvGH53i+qR
VnbSFPbK9oB+RkKpRR9Jkl1AqFgJqNtbSQ/3C2oFnW7UXd/jAhHVhZcQdxpFITY5
81cGEvlq273B3gy93bFDRIF3F1s7KbP/Ie6fV08p/NgMcujPRNK19l2WVgISaesv
nrmaEeXQEGoBnZmBoZGez0U3dqDlBEjmrCTgt4TZNZE1XixGT/CKzfIg8JyQfq8H
8iofeIhIF1/VbTcykrlrpWghoP6qDeKlZgk6iPdcRx5QSHrsFBbiXg+vjTed+JQS
hMJFbMxzvtTp8tZpJF4gJl/XSpJd1ctU05c0u/Y73CcNN0Rx7rFTDfetJOV/1pKf
7LXRBkLWELFbwN2X2f0WsHOP+2N/Iza5ag+01DuI33VuNIFJYkDfZ399mpT6EIxm
UxJhzBGMzU7FbOxG0vhlRRUV5YmMwcoH4nghI1or4JRvxaqSP32Ly5YzFZjgG0uE
V7EF6LGWN7w5Zu6xYuQYUs0KTmDzYj1BRCi8Hz1ie7U4mpaaSOk+Emt79pgZ7WEe
6lwJTi55eQmPlj5y8C6UoQ3eBzevu1UwSemMU6wVXO29u19931tqebtX/i51w8Zh
A3JDGijZV3jfviEGIM2I+Xcjm81hX6hmyA9k447S6a9CVBdq1snWAhMrUm50r6xI
rhT0aljYmCFj5L6epNs33VQBQjXLBR/tyY7dMPbhWEubxYfLP8BSVlWG++eERjcT
mwdlZTKXlZ5PPWYQggaElZ7I4B0ECN0I4jEZ7FQGtqATxLmwxIMd2Bzo/i+aVwEv
1zqfQojSaC4CcCWcozRvOMTslPeJ9vxUZKvAoognWLnPeVJ8b4OJYTkLap9jwq72
OVrmnuHSqDStIdQcv0v/ciasXD5WtYha3YBo2CguWcPCrLoeEHAFfu9EhTlYbmpW
T4I/DVThOLXdTfoE16JMgG9AWaqNpxqcvs+/fK+Oz7kqm3GRwtn/tcEahq/dUeTr
5gIh84PYY333EzYpu9ev/R65miz2Gtr3HBvoZ8fdgMY/r+SSjgHRSIEgYvBdjrzd
vbJlkJDk+2bKoqj6eIN+0FE3z5BV6NIHrSxEa/jEtS8VBquZlHH/fKRAewwTr07s
FjxAirdC8pieWEeFabBEdr++GiHKEGtnfrJnO8pHcwpW+RbrJASDdbaY6VpM7PMA
J68++pnoyxmDmgYRL8Bj47KBQNVEglAVpPbHP7z+z9rQqy3qlnWvAK3bY+hSsdTv
/fAaPAPBWGxEeW4mFM6txmeMQx3BofzFBTE8FJHCcDdZg4PzlAUHcDnNFARCIKHh
qbt+Ix2ii+w4J6G4EC+gpSb3u5f7iclTeUH8shgVJrAJ1Z3S8VggxbmPKy6Yey0s
XFBxDncnlBwMXs4K6CySgyVJW25fvVwg/1gjeSz6xHlF5EfnsUgx4HZMAG/7AcnD
PknyFv6ymWKnOy6wX+rsAHR3s8LoimaR2J+wQ7Dxn0QYOR/sr6PSTFYZhOO4Kyoy
s/roIXMW7fci/MF4JGB5nZjexQBhQcE58xMHuYjLA4jPFW9yjmDTR4ipCOBJq/X2
t6rhF4B5fHUVQ7Z44HbyKNkKvlV1rAaZs+NO/jiA7hzDmxoN/V2UOkBkX4oNh9zB
EOiUr9IvK+HdgmI2zfDXNz8fOlkXEXw+jyK+jpbN3fUdLhMV/VGMqbDQ4xvS72Hu
cF9wkdUQ4zJtxkqH4QrPCdqCWe8aRH1fMR3dC+thX7wiCjbUfgkJjRJFIXfh7i+L
xh69qdg1lap4wPjtXppO2abkICSbvUaxX85vJK4eE9V6BKw4heEQv+9HKq1MmRjG
Z4XYj69cYdE4d84Enwa3zUEgiq8zcINISLQeHlooogVPRWr9luqWSyRccmPRULDK
/mnc6stQqFbL0fqET5I44+gxy+m70rpjU7Dlmo2QxsDVFFCv+XHuUh0GOZ+FtdKu
22/CCnJbFUovdkZeqv8FWUrdB6IYrCzxf5esIplGCjqBmIVQh5DrfWdYgu+61zxs
9xyAHIdv6RBrpbXaWVhaDpYobJCF1bFHfG9RSVA2J2rJQ2pJ6q70+ZMsufkHI8nU
eq8d8bA3ma5U4D2nWh8xTVVGT12zyXmEuKaeYsKg9daUoCcyuv+aDmr5E35+fXKS
szdc7v90JhxlWvAiVUWFoWrnynfUydVF/p9pcd1/29PI/O2hXCRB/a4LZvpurITr
Tw8RvOWNEop6iq8tUlzbIozy/F0slfOF+0vJ5bj61g5Hj0pCB14/HDeNmgK+SAch
holcr/fQkgGrtDCptngEq0bKfkAamiJ97MGiEJPAHDBhyg9UK7GSAmrqTlpXlXmO
JUCkSZw71xEuAPokaV5rrNlP4kyXmIfGDg30rSzqFPO8D/ZOQv44QKr6LYR2fGT/
zVKnmKHDvSrC9xzVI4+mUxMDL8+tXsCKiU78S7Q94UMH9BiDuaCJxs8f+7OF9qFH
31spAZyts9Hip8xuE/sCmyHuyamh8miLorhzxPzBaDUAjbXMiEyXm7AgNW17fLtR
g4iHgOZ/fGjok0SYbSUN5yuHHXc9FmfvzVbDSUcWT70N86hEXk2oVTmZ5SMfKJmY
jl9eGfimE1rsy017WR52AW1gmjtBkE6ba/PPr2WhD6TGHe46xxtvn6dcdkX52f+8
yoJTYKApxBptgcapgvMAjcw6hrzAmkl0DHa0b20H85XIRLelvw9z5AhgG0uyN9ht
Miy3Ov81GaHQw0qNVf4mOCi9ocP+eBGpQxUCm0zqeIHK9JfEeiMO6bnW6vf7he5R
0cLqK3RuZJsiVSUoyOBPvb0Mk3WQOEF8Tj1oeMRzJsLCPjb81THR82soeiATwL50
kRw2Icm5IleFwQlkUqsehkN3Hfdu551OqSNBooZlydI79vjm8qdVC27p7MIAobiC
9JKRYD1oKrkyfGzX4o1IUIUgjZUDQcxM/9HgI++wMyBpZoQqo9owxLWV54vgqP90
G7xy9gYxZ/nQ4/YEhMpObNrUTb53q+KCyY/A63iB+g9aDsn3B8atjxmlyDCQRI89
8AMC2ENAbrXSLIPw9v75QG0GA/eLf2+UUkmvRk2H4Z4kHGYRJTrqhjnDCq5NAR2j
5HyzLEs0LdZZAnF/PUAQxHLUsoomGWW6mMQJZgHRoImxotAd6LaVBywKfDwSf1W7
YZFotHpc0JXRHZnPQfwmIPRE2xyOfKGuoh/+zXRShINDGsGiXMFrLoYsKcFkKrBT
6jFDlRUN1/wW9C4Ex2jnsa3CU89qle/oImo7Wb2Kila5vBpPhuXdZyVsrnyFbX3o
0rWvR+1PdCgdDDOZORl9TyXkYOiXqTFesr7/2U1MASBgEtAWm1lA4oOQxbaOvF+3
8Qpexnw3c+OjUQYFJFb6s+PUAgAPxa1nvoK7n8XsiG3FxFhsXzbNEnKSH2kzsiJO
YtnBIsedwvCtpwo3N5YMrdAkz5B0kgznLKBtsDugOGHHJH8M/F0kOSNudR7jYShl
ijxGNgqxLjFE2375+CmiVdRQSiAU4T3aL8clW1PdQEtGvtioQTTg0f4EkuMznjB1
9V3xr73zL5iFS4s5fiPrHQDg5zqWQYx1PA5Vdn4gxFoxJtSH0X9x6NgxIP4XHWPd
jbpCfdVhwLwYkCKku/9JS29M9M+BJEOurFHkuSNO5It6CLHXqEaRv5v6ZExqddB+
qZzyrNcABCVZa5TWdS6HB6e5W/J89rS59oydltQgfGVzLervcnfQQpOQ5tw5KkGc
uywYGmvSOKF4eqsXXIaxNIK0t63bUR45nsInbGlXQgVZPr+RGFkdXxQu9pYpiAEg
NF4rtKJYfdEP10jlhT1CyHnvyhv27d9adC8NpjT/M+kOGmPj2FJhMnOlFKcxt2zL
2vvO4HurkPZpqSlEGt8P+sob1MYzNVeA0RnSO2/bJZ6w+5Gy11byG/wWfesIzjMj
yoCL0TfYnNxKgpZDbtzqe0EcsxA9qn1xExpZVwuivmb7OBdNkc4CJYEahsCiZFhN
88jS91wvTr1kEJ0y8Y5Mejx2Mpx/su3qVPzo9dRa5Jx10nONGc47zvIstOUZ9kED
lwgcQtE+Wi2bEAwo6dLWgnAZS3naiJ29oqelOPkawKaFULuyHEJpMXGT19My9o+5
7VWREhVIcC0r4XKiNPx4m0Q0O3jQzQArnK7d82+sUWBxicSz5TqtZwuYUi1Z1l+4
QoXs149G9MvxQfDDERGoNH/BYm09XNCt+565tLNLtamGfkuJObPREb/YiCFPs6r2
wTVafzqqrEty+CfdJ5+EvI857ecb/kz0BnOFW5RK16Wg5+UJ6Q0bXjmZO8KuKTqV
hJkW7Zot3nFfqxjm3dRUamm5zYLVViXC2Pp+9PHDeYhS3TLo3WkFH+Qzmaf2dybu
bo2/6R1PXybh1pxh79wKBZ/aZs8qaKzJjEWhVOi4YiExJ9kiOr+IaUFq5r8bN6AK
HXTlZxgtGGX8BHTXALXtfQcOyAEqVHmJaAbvPTzMdf6LJmdMvq0FTzjUyox5mmq2
s7NSkDloNK58UgDe2h5jl1eRK/X0/tMtfnD2uXk8+s4N1cqvNtdkq+at1CqfP5HH
9DzZ4Sa7dZ5t6Ha5hIBer7noBGo3LIWmLi8vryI5jU7uGKqU5ImpCAf861eBd3j3
bOhOQFGBxmeofUoUcnwq0gUJMs0NRkq+44coRDObrEwTqWPnoPkAGQhE3Qp7L+/R
o3hWPoYaTko2gm0Osln6Kjsl3aboikWy8PVjNQJMrindUvvidYL0PzUvj7noLcM/
Wa/84X/uRoNFQxbWY9Y4jfelBoajRupTAM+uJ2uLqwVrkkJxgf/sstHJdyx6nhZC
1FFa0PR418vlIA5sMfYLXTf4jd4AxfMlbl8WoUcoMMNJ2I7K7QtfkqsBIRJchKsy
IF8s2mG83HLjokkB7Pv6wl/RNlXNTYX0U+y6OPjUIrurDPJKsutBmnGBxIV/D/39
OfXIH/enW8hgOz+LQCXGY4Tb06pN8I6irqeUbDesxWV9ejyMbuZ7ZXzCtHHrqk0O
VxrzpYHx2i+JiH15MNFeoPLsjNE345C6Fu6+PzJG2QxbJZYpgwUUZOaZD5WR9Nho
GWJxonlVEWFGe7bn8Cw1aDIQz6EeWDm2u+kLIzIwzearxV4ZZ2CInx8ATt4kJptZ
XjV4WDBkU98LieTae93ZgSN6dA8/ZC0+7Z5GBO1OYqYtQBAPVqwDBMrQwqWMRmM7
jV66sOLGFvhIlnOxxqhnWhPPXdEoXGqP7BSZnvyct32KaF4Q3apMGJbn4k/BYGeL
42cxLL4B9LM2gKh30VZBh0tFPTFDvgXDaOH5rLOE2bunOEX/KBMcBt7BylneCD6G
HTQ8NGcXFC3SNoCHeIGise2dkVmCDgQnQ9KCIcKFEO3hMd9/qxfyfdFceavDBlHm
+RYj1tHuu17fXNaEGgOuKDnNwfYCgWUfiYKrQ7oey6p4RYPJPUL+0d8coKBXIyUM
bu3f1xUR2GWiZtiO5Tivq9WucZAxVPnNsy1eKD2GYABKuN9/xxgCQgRtX/WPZSu9
+ttc/sHGf90eL82Rnat3tiQe75xsuhBJ0/QIyvUxX2p16xN0moUwfd58E9Z6V4v7
K+R8N4Rhq5KqEUN0eQVQbhHFtsepk+dpPzpIsIDdIT1ZYJNF1jTEVeetw1pGiTyQ
X9mQu4Jt7k/rEN1NvWafDh/1JR9C7Q/8vWbLBm91PzOxCycGvEVqBZwQeEN/FurL
xECwo7cLSyoXkop9nIiUwqN0dpL4qJ+OzvZ6j1IyMj9AUoJDBN0KmJ9kTMOFgTZT
FExz0MuXhwv+WKbJPFbJXBPGBgf4cJc3ZqKVyosGZueXsJhyRCn9G2LtSCknQZP1
wC26fqAkYW7gCMOTZoP4EN2ICbqOPIXAVE+wXncu9O7KC6a38BzJ2373tVl9rWht
g5Q6Z+HAp5fSoIXzNqiGC7M+4ESO0+wKgAXrOJKt/cV9v69oSel/3h2/OArPiiWP
SOmHKzkHaUCUNllaW+EkatbvGZ762n9sf8x0zLQkYJ6uyRZJ8+QRcW1xmSrA8lnq
HqY3K5/kvPD2X9FeMnKtqGRKTgsAhm/CkrdV6DN8gPtpfA7iuo/kYUq1IreVfdMW
VJCaHEIMt0zqSzwjR7pdoFmqVx1wPJKp6oRlr+TnyOJMZWVEeg/vvZdxqcTWsYKn
v9p8sa8yQGXsA4VH0Yh0VyrChO/hgXFFuEQTPfAdzdAWiPmvmORYrtLMnzscz44Y
HyFOg+ispg0ur/jM6dK0LqVqPUq/NeTAwcw+zLWViN8UFbSVZo75dhPg0dME+83x
yjY2nTZRePUeLZSaqlcuuhmBg25dqsSyL+1olf9bvNDxXOqnzM1PXRFqtTuLQK+o
uOfGY9Bk6jqLSqzbechz6NCYcobyZYF+pG1Odgq749uKzvzrK58PNE7oU96R2WN3
pzJgt4eaL094NnJHjR6+hUXFO+bXy2fIHOkG0E2rN+U6vDymUcWXFproE4sTjOEt
QQeXFXSLvCSOAI2QS3w6K0yfgtEL+6gvkomWKbPxzV6gyqp0t9i0NaEx9HY/2P/u
Pk9yMotWTF23zWlt0a1betxFLRPd30yOz51L4AmQIA610sYw/BZD/0mHIa3cdm5/
kkNTMY5kLSmH0m1wEIt18hUQoyAbytaSqBdFwWmPE+ND/lcEO9RJq8Ao454140Tn
fem5mDPw62ROQmQv7SfIQV9zfuVK61sxjpz899fmIzl+8TKsF1EvXZ9S6Wp2XZqS
HD2gyGmE7oVVN1qHAiSyShM2V29cxmTbjdj22K6JM6vejC/YK9Hq60lDo2mhWUTS
qm0mFIltY4lMFVnwjHI5PE1q6mDZ95YXzeXyzFOGxzf2bqMR79gh3eqLU23/vPu2
iYwkVuBz0Jupo4mMDG2qZRYh9XsRJiYCXiqVLqabRyF8EDk3L3zQ+znXiJm2DYVZ
2roQMtV+SP3MCES4ehJn9sV1fxlaJT4l1o7Y0gytj7pcB15j2vI5DxRyiKM9kqfP
llBiimRV8vpie42WHbQ36NO3jO01dcXBLso+MQXWkVv4fsO8IazDlDMTEaR0GoPf
J0aqY6y8r5v/ehlhRGHgFeHLL0pXN2ogS5MiqsRT+DVLcDlMEWetGRcSRnfMqKqu
mXfW8IocGTYqCwQRqERqZMOEGmxr5nn5FxKKP8rp7RVQnW/nxwUDqTPr8fq60QJ+
Sjpdl1LXqdOg1sYtJtpIVEhjK5m5ndORTHYUL7iLgaLbv8ZdzWM1vsR0xvlIKF/s
UbwYyw6C6XmnSjHJMaUIaeI6SUhaGW81h4My0ZHztFZu2s5xlX/8tZeGUNjJOS+E
f7Aj57V38hzWPrO3gMK8mm5atkokOXTrnYy5YhSQl4VQZzpQxN5l7BvfJTiARaIr
PhGEV6C4Kpml1p0EPL5SPuzEPhE5uUb5Gap3MAYVFoJ+SCuN5d3b0OXQHq+4rDV7
GDYMM87VYG+1IpFilUe3uaz1+fOJUMpyYT4aWjWPGGxc3I46Gj4WHrHedKyydhFi
CKJebqNsUjg4eWQPAuxes+F4t34of1r0cJVfcLoB0VMel3zo9b3CPjPqBvKT+9oc
eLYmp9mhh0iK8lZdMLeElvex+JLNNJvtOHDZMMP3ZuB9OAMv27Wf4j1LKtvI/u2a
B2GcNzK5G8Li8+or6H3KIkk9lVLi23O/ksEqCw6eDWkkEcTeFTgUVOI822/O17/2
PG+ICZPhfgSfoRQuOqwguvrEV4FHDp7t5hjRqmT3Cl42ZRnOjasOI+osNvzEbQkU
Z1Ly7Xb2CM6MUG2FM0Yljv6NIDCBSpr3tXFq+7FQO8IvmjKbQgLGpiiKzNuE8XVF
lx1d7YwAUAmor61gVt2Da/WTzpbzKUzpGkeZjE/uVCpPQvb0l4HVJD01IrquiMTQ
j2ewOL696fISaeki/mKpVPp4mWtFqThxhidXAgIcA2CvD7WvfXSO+5KFnPxUYp5U
lDBbP0KZGTYD03Foasg97m38+1QDpdReD54N0SP8muII+TYlfpmeY/6XGDb4SStX
JZkaCkfyVm2bgDosYtuZ9CXVQKXjg3i/etO9DtaX6QbpjqB2iHwKy9ByBrV57lL8
WSadXhvpBv0zk8t0Wg3OalECYvho840r9WX74L9/L9VhBFf3f90p41jBIwzKxTca
J7Mi5r9FXvLajB0v/3XBNvs/ZxW7NO8hfw7Sky5kgW2xWV4e13NNADW7pUn8nltg
/WjKaiVNtRa3ZJnvWEkEXRF/oPg5FFe6/uuNvZbhE0Y0YaVnWmXHGLIEu3lc8Z+t
XfwvftILHMUm+YYyvCRMBAkK1gIB9s3PJ4WO1Sk8yxiFNe1hmiP3yrUC/fz3O/zA
T3uCcOY3VdTPmeZM2e9r5CeRwdg5xpSc9xMbiNaBvldQMurY+pMwSqlW4JhWj4bf
OgOHbNbQ4QbBv4ZzX28mOa4Ky8QJk7YYbaHsowJ0B7sS3cOTpIVsgCKH+EvPrUD4
8PZFQA9G0xkQXq3xxl38EnmmvT1iYLiGrBTxHafLGRjKtOgclclw/E5bncC9Vdf8
f9dUQj0lrd+avwyqkW3oAszMg+AY40z/mPo7QcfJJFNbOri7wJs/h+LngqFx1C5l
DxuYlQHb71MTr7aAedUm34exBQiLUSlPKEW3oqJjeGm1xtEHkY+ztnqj8ogd/fxm
Mud8eQGGQl0XlAqfw+kV+POKfMCX8e8c0Wds4wbDRBpdCH8fRx2fyzygDka0m+v3
siRyenWuQxR3aHBnrnX1KAk476Sx6EuWgzBwfASXWSO7mwzNJhlpDSEfMsCEnyTd
Gu8i5PjKlGmt2YSDKN4sJv981EQBhi2WMKxGLJIJVYGmnjw/MHHDghb+u3hUuMVj
fcsYohUNfZQDr7Ck00znSYY8SRZZWL4c49yWUdt4HC73uXu3odeNQb6rD85cwViF
koaP34LM3rq0psZzY+1JybyEd/yMQ8LKvcFgnpcEdWLG5qk+fAC02sBlMVdS5Qk8
i9M9iU5fO7bOBoK5ThsXzloRH6JUWe21h2g633UZpEILNI/cFeyR7plAtI7RoqeH
turZwueHXRyAT1DODUfkiVtv8lly+QxPMUFvpMh2alSoWg1mfJ8qTUntxd9/xSYP
qLh6vQJ19hJoZ51eVVkafWoyuPqSXXbzXY1lulJncK2J8CtKU3ZkHxahbs18XTZ+
oSrUvzHPUo5pjA+DVaLmCxmamtf0OVC/LbRlPFxFQy1afzhcnKALOPZSUM5XQZPq
wtqnXe7WiP4JhdW9tyKK44z6AHcSQNIG7XN66aaCfKoJZXsV5DsCGBSRlBDmr32t
0+9kS+htuY0L8Lc3TnOUby6UZZgo8Q31LzLdKThurfIkW+z8KbSh9PCbIzR/gL21
vKOZOatcs5eRlpYROIokQ0Qn2SFEclPvB8G32lUR2o1Uk+3uN9a9vAmfHHP5QYzD
5BKyoyoIOE5lfafgJkznAsDYAiGLMq89PcPVk6AXauHN/yqM3zgpuUcHoIx+WyQ3
yOPUA8M+/GvyHa6qEL1xz2nWyYivgCU54S5dq9PCQqsjsmtWdZYIuVkDarm5n1GQ
P6ibmWvNL8PawcTTgYqoix4cff6SRZoYJLafYaQTr1tUdoRopGu9x+8UkJm+XcDi
7gZBOBRgxtClMqCtvZoMFpK8hIvCj6fuXbxXIkdeCSbPWgjz1vZD8K9Du3GGr6hT
0O2KRWk5k6mnreGhnzP6nTreery3CQu9/1YakCrYAY3gp1ldOkpqbHbu0xd473hs
Jrg9vAoT0lK6zQ0SvEmvglAlu2grIhPdtWMNCXoACXtix0X1LppR6NLPQJnuV556
htsKXf3f7Ahb4yYAcB/2A0os4XSvCk685SvJFY4TAocAt2yRQPY2cgQ5zDu1S0pk
Sc3hCh6GdYzWk7w55KgA/DYNkCMMPfLXIOUtRHQS1/o0zfssrgQDLhvBRg/BEMDI
1aidg0lRc77C3Kwb99xvhKtwSQlXuEcB93PFx1yTxiLOOgwVNnqPVbpN7EqP3UTl
OyATXYwomiValFdTzK/QUeS89mFFu05dGeACb6uA+zkE6jnUznkefy+Lt+s7/Aij
dnrN2zsAHgYj4UxJl5Ilkr2pwHp9l+X24TPObuqKIMkuTCgCQSNRDOIU9Sz//1L0
WeK4VPcq+ohabQX/4490MDxQ/22hc9HdV9PmvUlEyCtvgXhIFe5rFijwHeYZ/I0u
9zQW5AbcsgpMLpq8eI1s5WgUR6Du5dbIKhyzWI2YLLMs0icmzfQpNcos3ZTZzhJK
u2mUVSD2wVEX0/xLgHbQXooYRpfy4XDZuZ7amdx0+fqmVr9H4kNDwahlc70pLOk2
np2XxtMHMWeonXj4MrPfmKfvxTZH9kSvQu5KeZ+esVXTchIlqPX4YaGxseK+i6dQ
q8gsTtIphcGt5QgXrwwmzyPCxfnASQT2xPFqAF9fL7C3BfUBXAwIkva42Xpd3QL9
j5/jA1oOzwDZjrM3H0Qdje+FBWu8e0GbMNIvClLYHMNOOUd4HIbqZE7zEyr5zCJI
Fdfog442c511cFO2liUsN5P/NS5qFIqsLOOPJhzKYIZXD5ELqM6wJj2d3855VcI/
pDdhgFuYBpIfJEs3+zgx2MmuuKvKpQWIDLi5cUgwNIQwYTE+w6hWE+0b8FGysTA3
Y8sBhAxlb2EJxMPI2gSWdVa3t31c4ZFXEz+Br/kUs/9NKMdRotbalbuqQTpvNe/c
QFr4gYfEtEI8nKeO3M2htwBObXDabq5oSMGi/ATqjGtK3hpH9czGn8h/M7VYLZO2
A+B61lz+U/72OOy+6X/GAar2hDad2HS1LjixIC82KBQWLf1HcmzHUCbQ901reeuN
WlsyXApXkp2oTTGmojgt9E0XtQM4U0wAvV8xB6XD3Rf/YE/XzjhrZmmeijGbF/d3
NvS7rwl3lx8xJaUGuia2M9szmrVrNixqmlKG+R6d5qjSVDqv2i42sm9W+SHVhPKN
SDy1BQeVzZvK22zvtDJ+maZtozN3JA64Arcd7GlhT6EE/seADX/XGrWBsZxjMpsc
URmakF3e3ygK4+HaWYO2nI4SzP+bx1Orsr+iZ63RN13x1lmBYtaMro33QA5bp7oi
3C8k1T6BmTQSs4LkSHR8xhYiruGwwwBNAnG82l3x5bSxKgDnzZQp4CP8qWCl2N+n
VuRHs4KEJ2M011LWWxoF9uUjo14MNIZkCqF7HuZE67XcrGr+k3gjMy2gzk82C8Qh
+DT0pt9XMcZzxzyW+8mGrtYokBYmMxv/+qw84IDfIiTSmhV75SEH/yMDVjMYCtrt
IolPuMkLm00JhX0W3E6AfNnMWOf6MoXEFgmG9KQN2DAGm5UQu37oSkAw0imdfB2A
2MgG+t9XxXWoEzNaVPCYdHa8OODqHec7z/nRwqBduNt51lo81j5qnn2zXSJLhuLg
ORP1LAKEAp5q65dLYHTVsutJhlL83FyJKUCWSypmOErXIwmq8SrfHRdNBJUXg5PP
ot3dGi3KtU7nKz+gAqPm8o91bIHZc8CO3ntAN4asSH50kEPry20fQF4e5FwG5pwi
6lIOnTbqNxE/sk1orn/xXou7oz6bPonyqrYzZf/Aosqt+00Yf7PaC/kxcxQZb/i0
W/XjRNXVbLDuhbM6I6XFTRiEiWUQzfSRmy9dm3etUoADfxGp6/SV4zkfogIxSvJ0
I3jMWGeF6pl10bzMEDmHWDgqz0G7e3vNijm13/IB4yJsPS1h50Fq5FLOQLJfaWw6
qnD2QO1E9KVcIS9P2nYNTLDKpiR+7fcqV5upRBpAg8aLgRJJAAbqVVsQDodz3jRt
QUDiys48slm1uPXJgWKRjki7yAeaAJ9tFKERbPajv4ZL/owa2li+aC0HeFaT05Bb
HjbVj829TI8P3Os4XryRcV9bAtc46WmBKpDgnFW7RnHYzOPfi8sQ3x+Tl9OQnO8z
7rh8+Li/QfNiJtL5IJEX/iwLQ2zqD82kSIZ80dbp4ZbxrYf/eedmZEfjela9PAIS
9b3Rz9rKv6ej2cwbJsH695xKnSKrz9ipQsLX644faV/kNr7iT5m0VOokcd2zF1af
yPIXhEJvjmpDEINGnIYqFyc7UMsuudjZU7Miir8x9XibPqfrtPHjNjkSZLHG74dJ
X/GCAk80hlxhNsOeUV1Ac8I5h3BmIBjj/DN1FQmbALZQHSluQoNRWCFaOtf9AkHt
ksl6Y/5g5xv5RfL0Xoa2KzGTbO04xzAi5rwE1PvXgzdg+Xqir48q4eEijZYNC5j4
/EomNaC7xi3IoHumXL0skWp9G55817kuvyx88wBS7bOvbGl2/S8G6cdT9jAHv6HU
XOiZ6b1K7bNZv31Iuowp6luf3+N1+4hX9KjcSo1ElxtPB+GrishwJ9GxwLyKrcU4
dZuJ/VGCjwwbbQRjRrGub7tfvxq4WAtisxgWTlOP9IIt+YESxMF1bYwtUhaeUc7S
EjAMKKfX+ygL0CUNMClsaCSpiCXaZcXXUh/X0VIDV8zKt1Qb6J2QdcddhxNPT/Mn
VLbhBqqrWiuUMIxbIDnx56lsA/7KudMd9OLCHxlqKbxIpS5dhkPKnZEKgP8hn7YL
Q4E/CqI0/pj48GRaN+KnlklAiMRMQkeSURpinrEii+LqWUMMlkSCK5zVboGGaAtJ
tw2LL8L7dlzxq+6fChRPxpHUwlhWSgd3ufKBAGCGv1UTvgT5pmr/YU3f8Zr3BSCu
rrwN0uHIb38y8oywNIfzpdytqrWP+i6fLAirRzAI4y4k25M99KraAlZvq9LxbswJ
fKoI3mqRAYgEi2ewBjJ6HxGGwrvY8ENWZ/220TH7mWA0XnwQeaXV2KW2OmpGtJuv
EqIe6BFCiVQtiGggzTjhHwd5EjbvRpGnGG4R7pte1QMz3LNX+UCUdpzp8PXF98Jb
QK6itNP3o7hxPCKY1vjGq8qHiEkDxAwoqS3WibU8AwBbRxA3Gc7mVOaD7R2r2iGY
2gdKGB9UTpGWNwJPgvKKLXk9ZPm3TTQCLwME88i1EyJSRiJDuxgv8PAUy9SgYNjZ
6MRCY0O7zxRwrOtIzR359ttPMafPuC1kCI+TJ1XLm76yk0BWhB03KoodCxweXAGp
qgHGgy9KY/TU+omKO0anlnoMi0+p1X7VbBVkhFA113SX9mW0mMFI2PO1Mvn+byud
k6s+23hZ148QK+TY9J6XOIrMWbCBbamDS5z8YmPv/eY+jwgT3L9056HRV/ZyB7Xd
57yNy4XwIi99Q9iTuoUJGRy1bhjisdaDctjqwzYl3cD2B4f5ap/T/O2yy/b8IW0A
GPKq8tIkPqGhb7ePoWyiLpxoXVBw6MjGsY9SX+Tic+5sNWiscyl/E1OnrnAub6qM
oIHvjc6zCv5+gQPSZ8nmHZnWfU7un0hzj+QwBOFpnwu8+Dwz2iurHiOuHiZfH8Fl
2eXCj57YObf1fk0yOYF6VX6RO06cYkv7G7s/yiBvKW5vJ4CWqyAqiHPiyNzbg5iT
OYF9m1OtInCggbnLmzN0RiMmsW06gpBzEUuOWkjjBTr8u4ySOWxx1vN2ugxV6Lew
y6js3mlvjVYxKzzsOfAKLmOp2l5e2scj8KXm7pLVocrC9sDX7zKznYB9sqrz+xvz
2w5v+cgCpZUMCtStapEZ6OnvM2xFGBRPsOdgsB61+bJxRkAJPeRqo4T4hvnpzvNu
ImXlPpDa280NqAtZHpHOSsn9NgqKxe5KsrsYWBhZQOWGQF6gGZvj9RzNvjSFkBVP
gbIWU3VfMSjbuNf4uS06950MKa8yOPYTitgcCgzW/x1ndoDyHlSZsbTsf0vvkAaj
oOtExrXjc9dkFQmPNE9DUK9Hotshsaaw/PfJFAUpA5pJUAV5/Ry+YTny4De8xfKK
wVnDsGhbxP+ZcyE2/4h8Ra9ruO2vUJ7V9JKRNqKkd+lnQ2aCJZDUHN5rkD/iiLnp
av1jqwubkxcMhNtL7jGZBvxifnXVgenchMP5p3f3XT+CcxCgZAtcFOAMed4gjjeA
+0fuOJjwCcalrsOaabPwskEnehrdw2z3nMlMBgRPJ/kbPAIPsg0NQKcB7DeX66lH
DVJcxNqXc8KUvb3MCtKq2xCyZCIJxhzCYBwq7pMEwFa5Af55byVuOytM/QQGBK2a
V16UvGv2WgE8xAqfed+1RGidN4o2+ZAvfK9LVxoRjK3qlsgySi2x0F7s/nnMiVIB
p1IlAO79iYaWtlXUTn26k/zU9VxwJ+cATR4OeCu0A4IYHzeZA/kyRSyB5jlNnozK
UgD8brmzvL0xDkFvUGztRvW9/+pBmQVRlJrJUTswvvIlGp2brfTQKkV9dgkuhMJK
bRhsCmtIwJq5nAW+jt64RW0g7qkaaXQC3hNFOyV4dyjnBDJAVMM/uda9eMX82eH5
VfK0D2nVu8NfIPHA2kxLGK7Cz4HqTaZeqAYevCwI0DaWUa0KhJNwIEJ4EEY1sBPE
WAx/9c+hWeWF5qPxcIZERHeW9bMbWKvg0WpvBs7FcjLvauSRys3HICkI7Rg6rODl
Vgyd+j6MX0Zdr5QRoH0Net8ZlCB3m8LsbLd1WtAwfV/8yCglvaKZDvbaR9K1SKDn
DEXTD3oR1qFrq4GWajD5T3i2Tfq5Ux4Vo124RwvazKqAW5zGk39n7QNOkNbGplUB
NLsvSet6kre28VRDVGzNkO4VnbrUW/NDk9TftKfHoGWUVCfA1QnKOIeufZ9YXet1
pbUAIXyaRzpE2fKGHoe4zUTvGhM5db6jlW/Fzk1ZhjYygW7Ga0I1loSP9pfDIe7Y
bdiYTblAyFLXqYtQ7lo+CvG+aSWZLEJw9sYvAS7i/tULEOJQUuiTeJs+D5uLPGWi
nbR77acW+vPzc5T42r8R/oI0FzgyN43Rwh6SGrWGJ8ioBc/To889qIkAUtJkstlH
0eaXwsYz6MfJA7+rkywA5vsI5PDPHzsDFhOtqD61kY6IUPsQ3QJTvBExmd8jml5m
jN2YTv8yzIFWaae0wszfUYBEyXSGsNQ/xuyaqakjxuoWfgXfdxsVYdLYK1AeGA+h
C+vyYLAjedSI7RjLp5F6SZCUn52+Hdm9TwXP0X7TqAUFOJhSKyb13pq/2PCfzSWb
dgEz/8RHpqOdy+O7Y9L/wX/MNcgO1i/gwOtHXmhIS5yL2bVFwWQbwDjf023sFKFV
ubOPvNK3xEBYKbYTBK9zSDFx8/Xg+PwIVOU0ZUu04Lsfa08KZWsJd2Lw6Njw/zY9
ahDHynvYgQEoyLTtRf/8xDbuxXMG3lmhy6xAT+0KbrYVqW0WOiWWp8H2rNhMVYjP
/gQf6YP47m7saHXz3mQ0gAgg45XXZraycg7VeJgjs+bZH+DynOksV2QgqJraCtPn
0EE7Y71oVpjALbuzGaGEAKTDtTEo/B+uhimu4yuA87uURZ4zVHCqX8sICjo8M/Bs
G1OvCPlMV4IPonmAD5yDKC+HssSVwaSjLcNMjPgl3FGOCLO0oQg/k8BGZ4d1Ugj7
EFW3h3okFyafOK0+lJruU8cccgtHdN53yGntWUZ1J+5yi0FmEyLDCLDFeI5DyYAl
eiCqqyXcONNFxKuzCtLt7Qgl7Gyktb8CT9IDdZRdbPUfUdvjhU7WyfhqBoCgfHmA
moi+ugp/Jfslzxy0pMGokY0QyVx0DmkQkDetIvfwNajLCeqmvdX9o7p3Yop8Yd/K
mLNcnoCkoT+WCuwWMPMOj7xEkLWiqgsdjTDa3uKsLvg0fRBxAvjPt8eFLWwCZLol
QO/lce+6Dx361fXYFGLU6BhO2vu9rbsX6i+/SPdgku3VPr85hN7gRhIRjdOAVyh+
nVPlIrvPJj7zlmezygJVtYh0VgihUmOvanek+niGWYEFANkm0aBaSt5bhfYCTYk6
c8KAHq0Et8cEIwLUbfIJSjOfGEIJwOgLyjDeCOxqjtl64LkJF6xbMtTZpk/AfYjD
qf51JgwGMV87uxnYDl/MsIZrPTIPCMFM24LXDrj0sRYLr9+UfLt+3N+BTVMqTAuB
JXWucPrRLJs5dIYRIIjXFaeW9xlNPBUvA+p+BzPIK2/kvfMGLgSto9QPEk5zkqWH
XrlBCcjVsnvo6gpF0MPqwsYFIVmrnQMmDq40HxsJL5t1ehuSyBpW+17RvUKbOk2J
wStuDhxA9pD2avu+No0uWKz8KutYZysW5BFHgVFzR1Iy0WW6bEnv6mlbq68Aen4r
a4RuZObyhbh9kTMGL5iqsPbjMJMrRiYaqL2aFTGVuZwT9J3Fni3+CJ3RYqfXdzeD
kyn9TqZIoUS4vV+dioWhnBkesyfnV2jZwbQ9AYOdL9y3YJX7eEkF/m6x3jXxALNi
GTFG02MBiP9tWotvslbTRNVGNNZBcXLxC36YxUvfi68Y/sV8vc2QpxtZ/vCotFiR
cTPfQM0su6+8apvG4aESb0DIH+5s4rriIZuSEhfSlyaTjPHwXhTVBj7GF4JjR0xf
mx5yWXH9xoW4286HwpvHdSlBUBEvYMtnGL7o4w2nWb/smARUOedsy03WwCS/bToW
m0+oIhDCl/2N6Gc3BKbIH/t1L7xErKophNAu8ZsspjNu9al+1ThdGI1gbTnM0jxm
k1y7eQsW3dTKvp4BKii3u7/HDB+KmWcPHY/O5WpUNen253SwgSo19fs9hrzbjjh9
7fGFpECKSb92NVhSxwJTL+cXZceWgREvXA9FTj/8zoRjQCVn6ISHcRXSls0FpQoW
LAQSEZNUcISLJ7PaQypVFsl7sQv4oIdR164UnLh0PqPoqgLn1GJaaBpe92Z6cCEX
KRYqbxapWmUnaPqovtn5GFQnXOUX+CBC2xnonHsJoEAldVWuSjLWA9pahMwYctHy
TNcJkyq7OxnGyZ+fsWeKiFZ2c68Bx3d3yynTMW6MPbOyoCPYP3BnIj+4BqNuzzT0
ubPkzBus1x9FALzjJxwnXbo+9L8a+b+x5vk6VUtykGW8TtI6n8mXyd6vPjbQcl/h
cp6TCKgXRGfv5R+qj5XwasR6wdSlfG9IguPrfihp4Ebr+lMMY82qYfCH+1IWltlL
CrATxN9/5/DeavVIRbc2Dd2tJ1wD97w1SoF7K/vG3ZdPYRttnD57eK3ubKfAmCtE
75Wg7l0CPoxzTdzUM67dFRy7tW4SNdlrbdg1nBiVfuIMM/2en9dDUZg5tddUZ5NT
lb928W9NgWiswYItKd9g21FmaAFPt6czhrVNAVhUFrGsdQZy2SpQBz7RdGjkposF
BGkstc4Ud61chog84ls4taydKAwp4C+6hsxMs+R7bVEjvY+diWSFXky5atPOdSy8
lgSOH+eE4PVcQ4sfWHcsIRWEjYxfg2vhdV4jqWUSv83oLCuAO1/PoxAq1EO4F4eW
s69DL5e90G+SSisY8vY7ZeSStlFjOvXu+A8j9M9yDjB6GUzbGlPSKKUfSywIrEm2
/1P08VJwyswaABOOG5BQYQPoKE4IKqQISQjUfxbubYX7eZTehZ9NJ+IOQqKeNY4o
H0Ky5wzwAE5cFqcYVI6CxRIwOyIjebpEMddxHE+2ExBxukT2IRviXmZoGovjfCrn
Usd4WS9SpP/U5gRYACV/m8KE4A9qfBAWh9ijcGJnVvFwH19/Q9+fvcGxMgSMZoZg
x4gnK5RxJbeNFIVo+gBFbZ/LsKET08cG2bFEdZmrq+feDJkG4spwrDZ0OTnQwym/
0MJxosKg/yIe7vXhJLgqODf370pDwKBNJagFiMhh/V0eHZMDZ5QdiQVnHfKzWxIh
1k7UDQSxQApUiHOcaqhhuTsCQl+kTZGV4j4foEn3wse78rhNrDkpvxxUpyBYOfN+
vxEVqKSI6HRLCUEPADl60bzshFt0Y/pBmrZeSKUjQv1QS3lUMxL08zgLs2Kd7ZkJ
uPCzOW9KylGiErztWq3ojVkksYHlxasUPH79f7V7asEN7AtkcoO4mckkuPAGyJs/
DdlPuU4DmVwM6vc5zMzTtT3QJC7NKWKaxdNo95wboWqqa9CejN+BwEyvp5cC6Zw3
Gxh9KL1IEQu1YKtwq21TWm3zKOyPjADWDSj9jpbxpRdsaOb3KCQZCnOcT+S19d2i
f9XYGyHia47NiXgOxTVwdgFk6LqKt5lMovU702S5VMrm7tGmefzjxm/r6FgyNFYi
3LdQ5CFrcyCQeuUT1hvXg0NXMtKXgSCZQ+qmByqiintNpaTp/GzfM84toOfilDrg
DbXQqiFrakLCZ+fodNB2Ig0Cf39Q8XVnjsynSZD7dVGE5aySwdasYe00huv7Ul/x
7EXWmRiYAlup8ZvdAitsCkKhBPK5YO/ztNm3ZsfS6cwOzHWudDYzrhOyVGtalTYC
FnczE5seu1bhA0rY1by40qd54U7NjnlMo7OmOoQznUgpRzdR7MZ3lXiO2lCJtRYy
H/VCkSl496W2yJaZUOQJ5Ah6OS6kBUuKpd75+5wK3+z75dbW3vmQFa/RvDLn0P7p
GDvqP++QUzYQz32pPsBpmTg4BouABKbrdsTKMfboWxzGyRHSwbcWYi3nvECy/bxX
WHCUZqOFf1Q2Q+VhRPcaohXL4ZmCZ72MC3uV4oj58f810xF9YLlZlw4XV5Ejn3LZ
OBvL18PIJg9Ay9KGW+Ga1zC3Dq3voAdhGWZP8t6zPzun4EypUqc5ytqyk54n5q/e
r4jVdgd/4AKKpOpj3ktyFb8AQH9ZKBQ5LEmuYcfM6kPZUXYNJtJ86Xuf+xSiaxin
DHRclrBA9zgdBF/Y/N5ZN/0w2N/wTmcYnOHfKBNJO1wW9m2XJ9GhR7ALJKJ2PwAF
J1pXNsbDs7Rqa79vIhcF6dfwXyYSe7kN20ffhQ7HAPBX4kDghXWljEkmLIVUFzA5
o1AEUpW8SCi1S6g6eFkNhyNlgY1ES07GwKT8a8RweInz0jJhi5m6Lu3M8ma1B8nE
4vZwxejZ0Uwmi5hFT+Q90iT+DicdbZfCJrngsQsBJkL4f+TOrOA4RzFFQdzlLQxV
72+ku7fAW8QAf06Qjz6Y3DZ9yLiS4TRu2CsjNz0QBBhuP6zM25EMs3H52/Gle3r3
x/uaW5t//FVoEPvJfXRLNlM5gbgmray3PMPvURJEYMW5dt3aRfS99VthqEynmBhw
T723HopvBch3xCiAKHsTewx2iSGChz6Hx/LJDGp8hvrK4cDCQ8bdsXhSo60FVyl2
kxMouORyzEye8Q3MnBzXoOegWYXBWFQqL4ay8h8txDLsF3g/2v8zd8EV1qHQOKrf
8AO06jWoF4EiF8pKQ8dFdFBcpDYoRjWtKrJ3ye2X9GUf62kgw98wVroC9oUfYen4
VY2lv2Ba8or5OeehCPYpPfj9/XWSr3KTTNkbQYXNVDFrynbYLWOrc4N33mfXCtYo
Wv5Zr2KIu/kbGmAIQpvCSvYnKRiq9fdAI132/YyxG31K2BV8Orz5yxz9BmsRQJDC
2mb1QnEC48P6gpKqkIcCw2RO3/X3x0wSwtrIk2yZgS6tfQD2gPBzf/9rSp30Wujy
eg+xcC+qPl+OdCmOKejmdxM56sx3joyj5gkFjT6YV8T1tPD7KzE0ajGyHX92IBlv
8aUa18eFoD/yFpjc1YXJIhCLEKw7OlRN7gBbQxoOG1AzeiapuXnEi1d6SznUVpkF
JuNQD4sXLXaimD1Ib+E+g1Gec86QM67FbQ48egOkIWTxVqExGKYbXV/V0mME6W3d
/xtgxOs5yPoPITRJZWdijxp2gJmM+jdok0gat4yimgHCSS29yXrKZ0W1oeArek7a
r9cuzeK9TXAzKnRyk8/1wTlx6pgyEdd9QvYypgK5xTUIgYwzx6DSyWuhw5qr2CYR
2JZRj896/YpJ+onL0khtJCrt/Z4aNzvaumNO79ISz2vHSkTXwZwLHJWIxDZvJdTO
+W+lXuIRdJDRXXS6zDqxn+/h40ZVEE5EgjloBHzNyGO6CwJonkJT/R8OZISAvA1h
5bZ6UpLUaNqnpxb/HdG8iTwl4sCR02ioI1eHI7C7228LnOqHoBdiBkLbahN5wRiu
Lg8X1vwyyCig1lw3sBdxaxigIFBKwLT+9HafdRnyJBMB+3pU2raf0PvcARvLYZcu
4yHt5S3Yn56YuAZEnrxi2vpRL9tbfWwU5UdEoWV0KLdl5Bcz9mSmw85WArUzM3Ho
shIt1PYbOHVzlgnFZ7HFSFV3nWt7ABxnaqL4YaADfzwkYbKkcHjGrQKx7u8SFL9/
rYBLVyd2im0Ah0Nf6c3arPuC3Us6Ic+cg49B4DVIdW+B5NQ8jMD0u0gQ0auWEVHj
k/8Kxj7079JtXgcdSP/w1GPkL42zNvKOu/6stSiHqP4ijJodgRVZcTEVLqdl9NTC
xsAWU5GEJG/3O/oSVTBSokx3DzAe7MwuEJYFBb9AxYEtfhz+H9GZ3hJpcQrcqVaJ
HQmUk9vPl6jV3+0KXnOJv0YTPEq6ZAFTRtQyKIsBWh+TimR0q0N4qMS1IPcr7Zab
y9Ls7j6vabJJaoidl9hyIFu88+CCes3k6JU8dima2TG1QHs6TmIwWG8YN/mbUeGD
fZNtisYx6GILgWExcP02uk0pi7Mp3D3YYpJjrFYEOa9oH0xkJtte1ZmmgZeI6O+N
kjb+rO5pb/H64Sp6A9ZX43ZDvpF2zasVzlEBXJwIkj3Q6miYLFpculeN6lXyx2GG
+o4nSylh3tLEr2XLajvFhpiWKblVpDdkZf/qwYymCZI/8BPwxMDZjQ7/lG54eNjj
YO2jYuAdAIHyfD4DghW48r4hSFUnO8+tEqqls+yiVhjZujlKDuifYZibeE3T7wjc
L0NwSOCLJyLQqBgu1vxYcqbXQjycA9j3Ip7aZGr4kcbl2QaBK56qeTueRHYgs7xV
SUhzV08lqgR0dktVVolQW5+IBu/tG1LncBU+1dKhxxd0LpKIO/SdcbfJsgrH/gH6
Hw9Iqeo+3W56aaCzuWCinm0sFP8ZguoRX8RGDN7vRM5xp83WRKZtsoadLAoK2+57
A/x9/0pcjzwP9ASI08dprQxhTKSMrKBzZfo2omR3H/p762rw9PH9HVvc+yFlpF9R
Ce7McVQFJQ2BSzg4TQLV3+eoeOzmhQpoSyNT1hAS9TNf/09Kn+tpd5Solpw1z1YG
uddUu7PMUTe6M2b6ZzdvI0mS0eyT6AJFxEnqC1fDAKQiJm6ZHrDx1bU8xQ7bsgt5
JdzwwxXM/rKD+38sNg5iHsxz5DHsvdmAIPLdI8f51NrFwXZwB+vFuRXH/DWX04ND
OZwUuxXBolQuSOvzxNWjJfNf4+HpIkLD6bZWCLMRnJDRCKWZ0YW3y+hE6LeiAVqM
GyBrSYUMrg1JjAqsbYasfEQN7vHd/gUDd+hfVQ9ojrW/uLDk9d2p1Kh0ajE2PWtE
u6ych1FBpYtPePYgR8b3nHKHeYmS34jI+C1XJwa2oXdXusZWpONN5WXUtjd++Ns4
iyD2iWFG7mYrKU1G8NzYE5ZuD+WVTsUF44Wlhoq2KY3sjK8ySeGB6V5PWFY+XVO8
Bgug35+CoTDFCxcskKnIPALpkIwSYHG5cgMIoKI+qpngXDjyW2kyBhr19kKas6D1
FT5I+arqFAIjWgBR96e6Jd5kvp90c1bvPnbgZkbfmLNjC1/i7T4nPvdj9pCnBVMp
U0Snq62bF1lGQ9BJkQqgiaADohXrEzygvl3daKNSk2/NFaBc7oW6rxAmhOckOhj7
6dCqfoa6TilnQnq2RyZWmvneBNijnQhTeBgGSne1A5D2Egsi7uTdIIY8zH3faawr
NyKHnt7LB7OFAmgO7s7gzQJVAlpUIUWI/4Nwl6Y8UQ199x9OlTboQ/76zoIVsrcE
59tgyNuSpke71Y+1mC2cmrNKRnNGWLCJeNsTJi9pw3m9j5FMQu7N6fYn/fO6Cjn5
c2/SL5Vx54pSfEECZ7cgCOTNWQ64zt6t1WG/KtRcdV1RQFLUs5Sa+7DExrODSjsc
eA44Dsa8dfe3RHHtu2d+Z3Cqu2uzL32t3x9z9Er5+X9aZjQH/hzmvzzbbbUNxEe+
eEuWpefSJUqBElM71wKQlzzQiI63Erwhjt7TYH5OAPd/zf9AYcdMzpKK7qoJfiND
+2sptHnK36xXBdjqBJRMJUHmYHrHa/MhXMip5J0U/EPs6RAS6YWhlOkF5ZK6nWlJ
QbzC0JrwRUGhyROr6vsvsd/uh2nBuw1e4f6fWV7O9jWNYW2Ia8GzJv3DhQc4wDtI
dzEWCzv6cEH/niW2of/Ytk7o62JRBLmQDzIbu5ou+PStee1qnKW8YQuFrPMuYjCq
QPfbDz0RcE+aV4NC6FAstGmTBijBBkHvHcztDJkFqfu0mBqgKDGdr3a7MlaUmW8A
Y07XeqFLH/H4Gxiv6Hy/1ZaiZORY930ik2CUKRxadxE3n+AxGW58Kg1B5MePNgcK
Q7RJabRTt02v/lbDGPVW/vlZr3a2eoZe2tVhBDij4iFijQR0A49wruAom5+9OTA4
SoCxfA//rQzWVgyug7gj6iX2hRJuJLKZh64nkifiMvR8MqVnrgLnA493FMiJHG9C
CT/x06eSDyXHIBexi+07Wm+DQ4UASsJSxBXR8JJsMGSf7VOZXfMbLDDRL1c+TWTn
aQ973x+fZpAdhITjXa5bsU99j89YIrEuyW+Kf3/rVFXCYk6szZ0yKD6/nhRym4TM
sbO4uljNXX7TWWIORmmGPu1HZ9H6K1LBxHPX//RMo1mTnnJRTl0C3RNT/6d7xQ0j
cp/I6vmxXdnZ03fdbBg8qiEP9I3MJEMXAAsrGBkkWrjUZxM4PeRcBXmszgU/LuP0
NfD390zXfIh5QRtivbm+ul6xB1wbUJOLJ1uNgKwoeQK02KemARvj0+SxO32rP5zw
uK432O1yGgr3iuZScfdnCyVvpsD2i2SZW3YnAQHZJrX33zx1WWKybY3MM0QWEr0C
sjX2AyLGA0mnRZZ4BPa0vdy07HNQ3fvc82y52R+kJHjA56mNNTJAXm9LR5bgVLDb
XTgS8R2TazXtY+44g30VwWESnXUQw4jwMNg3F7QwFjdqUusyJDPiPTmttNiU9whc
fkiGxnLXE1FeTBClzjSsI6dlBH224InogAMBLvwX7BetrQoEXNqodAng74E6sr7l
+zwIYjcvCZ1E1RTE3GmyyM5CMS8uRfO7VJU+YRiqlf/4srS0xuWKcqviBZmYIWWm
ROzbDadOodI3633ZsP94wbYveJfyuJjVuHIpvuacMAxnIkgqtlDzVCWE0XJT/TNT
V560W/tvn2GjDOZsWtTJN/6hhAMkQS/yDbD/mDEbZ9zk+KyMmrYAv/+B+RhlRDXe
w4RnsAT9pQNM93AU8FYqASZU/xdmNGU/L7qmJob2cPKUkp8u+OWKx5Vb1r0lEcWH
/4trFF4UgvJKXe/CV90Zx5jeK00rGipaTZEbSLRjXdZjStCgBO8R0nO5CRAg3psb
3EIZJdNORpxN17LMyzeSmhSmASt6NlyZF3pE9cTPFlfk3oKoj1AAUiYoKoWuhfF4
YfpPdocNMWAW4dXpUUJ9c2I4CrO1XH5yCloT1Y+Aoaiu3oDQhAoeYpvb4pSOKsAX
AoimzYP0dZrQv3jS/CS1UPmYNVuKNqTwRuGkQfuErp/fYF488y4MFYir6usDql3K
JIksCLI+h5Vsj+rg5JcMgiJ2MYWYwqIewA1xqjvkl54gZkMGcSLdgvVAG/Bif4qk
2XqvPZlUDGFRl4SEJ/8H2gK6neYzIYBB2gCRiiwecrdAy4KHnlAlGw+WsNBW5CG5
y+pTLbzb9jUTUUMJo5TrRNSV1lLy9mYrbsV0aRo3v9bJOT14m4temMo6dcVelB/b
aLUhAb9RvDS4WIpWCJAJqWC4XoEvAOLjbKWOcCzpfSd4ZeG5Vq1zA11pTlAHLt3G
SJips2gN60XWCpR++ONIs4N3tq0H4OAuzYhrAILOJut6Oq4wG7ZHrmidajF32uFF
FkoIsVBsqKhD1GR3Tg3ndA4R6ZGfBOF9yl2fIvKBMqbcVEYtuyvlW7mHN2770wBR
azzEp53yB5zptjMXxkg1ep0iz3mhRcyJwMoEVBHnweoinnjDA4kRa7kqGdxm/yWr
vANVitsaPC5U7FxpylWN2hp0GdT3e7UVuyHNIA0DV4dOLTKbfptSD6MiltNpfwfx
tzquCiX1zmWV1mYC2mKPSTOMP4Q5tmLzA1wiEQd/okcUmp4mkIZa4asvjB32Eqf6
icUeLFtB0Xfhlr8ZE7783FlAs357XKQm9Bk0GmvlcwOHlpCiVG7pNQslhMjx8bJJ
qFopgb+VgrfPNUMDqq8d7dZqTl1mjQNf/G/wVkyMkUNT/7Y0CSSm2lrDkbmWQJL3
MJmcPw17cG5KU/tNFqJOJZIO3Qd3vQr8D6+48wpTU4nDrBoIV0WjGM3Psl1ebvwI
oy0T0mSyItyUsos0yi0QGVUcSPwWCtmadtyDaCc/n86myuAWC5wbjtOL4m7Np8T8
HV2OjYZa91rp9M0+CaErAeONdjUaH9R5sZ3IU6jN5YV6k+SF4hXtpCnt8up0olcs
nBU/vdof+IOFrER/7S8CxP6+Vfd7e2fDdhd7XA5PmS/ko5W9LEgi2SsMqtR7gK/T
mgt3BDwF8Fn3f/TaJ05wXoJKZlLF0BUNwaWMFnM0CLU5UgOkdHhJvM1xrya2Jitd
V0dutwDbC4VkzjF6+5gi94YEps4GZWU9YGTl2FD8uOroiNHL/WMZrxskFSyU87XR
FwYPPFVhoPS8lNpXMaRmEqFft6kDBQnR2wm+2muWvCJxhxK1EjZrvHhLRPpbhX42
a3InX5kzwrjVFibKg2OcukbIo9q0Ty+A3T8vO/qCSJqxNvG0Dphe2y8RHd5K6lOX
yu2WAJI0P++g/fypF/0yrO86mnOdY9ngH3oWhS8JV6ltjJLic1+bwPo+UncgqKJQ
pzyZTTVFeXLZSfzP9aSwzFVcEvJBug3wA4kIRd2upwPVF5mB7z3WaPtFCi6a2cOI
VYhWmG6p2zXEkyzsUegV+Rn4SzBiS+OSSsD2MYP1nOpfk1k4tRxg04Lif4YFWDqo
TPrphPJHCLgBT0UKGqvq6hCRFw6kdZEP81VGtOjajMoNrLDMRKUaEtpk/B9NMJIw
qRvds2LRLf7/i1uGpVpmyUr79Z/+StghSL4G2yPP32dSBbR1eDZXr6M/A1zFYIK3
mMNzohV2opDJE58/oAMBDVkesSGoBOzX7E0rtsm0I3oe1HaJs37mHClE2olGWD7T
zlU8FfJq6zhHE0Bks/74edSsbaofMCu0gKJQXngp3zW2pgJRdC5hBaRFTmAYA2qI
H50xE0ww1mVrVjiHIDtXssghlRCjcEmCEpFkTcfMhZ8e1DpjC/0zctqhy/hKXUpJ
BV2TrtZUhPNM+kdRfQYFNuyX8iq3nl+CpYUlmEIXr0kjkkDcgzwUD4Zpr5HSBP9J
KlR8Rxfa9oomccA9jkrY8xt4HLIxihF+i45zb+X9UMsl0mIXV/HOIMges/LbGLMR
dcrTwbMmMfRsPhFBeWD7MSriu4/UbWtAOHmHdJPSy8RwDmCL0SSx36cWEcS8B2iH
+knycTSEZGWJUiX66DefVzQsPvHIfLu8Tc7h2g0sOisWPheq4wqPwkc3myi/11pr
H7nFFGqIl0MjO6fg4VKulrD+sbSQD930UOPSLOvpasXpsIDASFjGFpvoX9cN/+1b
wlcrQU6zKmbzG2edWW6vA+EJycWfXAzFaKEklMrNPKVpwzeYE1vgqgYsGGATNol2
jDIkGjP//SruGv5GtY8wc3ZdRUpsbKgveqImE2LYgJ7lCfGfd7Q0jjDugcv34NF/
mo2Qx1f83TiT0SxI0NOWY2LNNGfPPsDKDno5zTfRwkYHG8YfJa9bXgMVx/40MEzR
mVXvRXrFGzunNfouSJT2M1FkrXhc9D7VHrHX+H8kV7nWFmhQZ1RM1PqQYv3DrWtD
r4Ikjfg8fpogQFFotvOTe224DumE+KooptJ0ke7DEUpH8mdbeaR46NZ3Yx/Sa/+J
Jfy6xy0CYmjuwGcVOkGTXX7RKy5N0ex3m4VqsPBIQ1ejOjUkOGx8Sm2kfWmNY7mL
jP6o2lQXtC48kxa87ZsrQnLQ3KjecgXs3W8U2Y1Ihz7Gf0MxQXvc/hbD2RiwNbpu
cLww9bx3JCauQEw6Ux6c/Yv9SPcrycJg4ndbF9tE7nKA58nchxb+hhFaHH5fTn9l
FrGEXbcle2JVBI50m+HUc7nUCulJHkPkfPbpT4Arq9iQ87IP5MSudtFjO1NzwCl7
NaDFVnqDGLWEcgzAZVym2vDsR9zL79gq5KrTDH4V5SR5PA0ZT/zBwM+GD1OEdg+0
6OUgtFEBY9RvdHrT9Y4UTqBzYktEUcJjm9itKNX59jNC0Ojh7WEkwo8tc+P1B96f
x+BoMEjN6ARPRBrsNZkARL6J6VZg4d2NjgfUN0njYMoFE1gdiUdvd3Ed96u95Tep
bEtw9awM/duwzf9DVfJ9+eY0JOl35xh92QQcdIWgPxcZGGRuUulvLBgyWkeMx9U2
71Ziaapt6O4I7SJeWZ7PofL73uMCk8XPFG244eubfKrlK4i6Qe7U3CHCgoB6/6wt
J+yxUvJ5zUK5J+yntt04ZTLHkRWqBQoeKp+7vRfPzNTwqr8V7Mnrp0BFF7SgjySf
wPIIoeGAINPLKq89iFFRkvPTKmJASX6hDQGNNlO6kHU0AZ6VYaBsAn4aE4LUXDSi
SaecKZkXYU0GQWWWtV9lKIGgI9Xa9bL+86beAQU8jH5H1JbBrDErySlAgC5uaw8C
RKJz5lNQO1POXRqnybLAcyE+jEp+BYUFG8as6Y4TXI7geEaqpJvplIAHrpmTGqmf
pNSMj33fwoF34upreWsOJEBDD3Hr+y+1GVW/8VLqAh/jK4/TBlSXboBv02qrDiUa
OZLad7LiMfLeumLbsuOoAjLLsfNsKEB/FGyA8ZKpaaRlIs2jYPNT6zXZPQsfQBXA
ILG6e4e/H4TjuFJrt+TOxtTvEpyx/Xbdm+ePNlPugN2SIQ/FTR8ghiZvC1Rt4NFS
jVoZFEQZH6rT863KR+MVY0o8ELRMimdGBuoC+p30vdIttY3wyMDXDZtg+tmUN7md
HTAM9u0N953u6lpZkTCWkkkq8IYmkis+JL9TdNBlGWnepnh08AXARdU0ETtUF4t3
YiMYshC5kKs95e/ixTo+1q2Nnb4NLVTf5gUu7Z8tmBoB3aVoGIvc86hmg8qYBGw3
D1szOAavpVOEEYZyZdfHvZQHYqxFDfG8/bdyvxsRYBAoVgBlBiDzIh8HXJKD1HhL
oT17xn5HRs8KSlZg5l/Lpg4hHU4kTtpyQTad2WkN8n8wua4nJKQVbJGR+EECozAk
rh+YJsBQquUSSwEA/Hzv6CvFV2ceq7V4mHhdIhqRn38+MDxRpMjBVETcAfJQWJIc
+1jkyFBRCVyQx4cpkmyBM1M8wuwfBGo2I/smq8mKFU/Q0kDKrAdu7w4OrS4dtnLo
TFl3UPE7eayJIspkxVI1wxh32S0qe9HtXHZUjMCEj4oHe8exhn0bC1MU4S64CwCl
YDsnJol76/GskQj1GFlE8rPjOkpJRmn8hWiPs1CpuudG12r32B2Zz9aMxvO0V3Jk
ZPBuTP+a/6FagjRZt+84ht0Tp6KSxwelFpGVNexoT9qM7w7dNiLEvgrBBxnM1BJ2
N1VgyRv6m8JVmUVPp1vMnkKjQa83aZxFI1RCb6u6ynjIfpeU4JcpItuihsYYoYit
o0ASrv+lC+GnhdZZIxRLdTlfZjBHU74ZkZFURhjn3WtuoBZQnpZT+Lq21dhh/7Sv
mqRJGlO3bIhrMtHO9X4XFTrbI+IJ/ZMY99CoriFmYZFkmSg0KVdUDGW8sxL2Xn7t
zfEF9SO7DigToQFFlj8Pso8sgY7eZfAzkJB7RCyA0BLkf9CDCaTJSQIQx7NjgpkI
7HkukupRnmM7JItgCDfDCol4Sl+ymkGOLgy53gl9ZigB63H7cM3cmN3jeOSIrwHb
uh9Sy3c/3MK/1g84HQbSBoq965ueDQLThwrHh9NjwnK/Up8IJWun67eCEJV4xHdK
Sk/XDBH7Lj2ZlXetqhXXKjJS1rlRHqeuoC7MJbRD7RFHfZWcFbqZqbklB06aTHQQ
l+Cdh889NFeuKVe7Hnnkzy/VIvQmRus5B+wtLPVYH6PLbwE6IapT6zJgjUbGI5B5
8ejRkcXXecf/0KXaFVygQ4hMWxXt0VQqgPEPesOCcX3iVR+B/7unk6hPUe+IzZA+
7oI+uV1qR4i2E7LFF73wWF7Ry3TyRt1WgDNPpeXyKMfv4jQW9tFg9ARBQYNMxhvM
CURb4KGeUKUT+Pp92fStzU4W7URlXYAtQCWaMjzQXMpPwrFTtwyzNB3jx9RWfwyo
SeYVkfEbbGTXyw2cH+pKgUTylSltm1quUMKmNvNyA/O5KAkC0/LDojVIy2k7Fzih
t4n4YQ36zZJyYqyggL/i86ZaIGogsW3v8l/xVh3KO0ZRLIyYzwRPFRPUUhfwKrty
Ot3aR1sCbZP61NVb7Y8zFyXhLenxcNCLDqpnAvhizH/FgEYiQ2o2hEkhoUunxgJ7
vEld39GVd/I2xb6k/V+59r8103p1JOnLLoLkW2UTs2uHDHcg/VJRuMUbs3BDtdwJ
AmA/MM1KVpUAEOt48PTEtBfxiSUqvTjlwzvsbhNXC+nkp5fOWcRn2UIY5Ec1TONk
aPWOeX5faoSj6cgqf3W4JF7MNQJ/9jdit8vcT+srYAfWEQSyDm/FlO8VNEn6zi/A
QhiyIS8Ihr6zQtMBAX0E/u4bk9ojmuvTtiSTkBCMNg5OojSaU/XEZTtsDsZM0hA0
BGC7tFunGYNS4C3mvhJ9k0ZWqVlRPhREILE8tj/Q8o9sZIx8OH9nZPm3x9orYEkL
HCAkJst8+w8VliLzcP8VkUcXyk5oCBBU35Cm7ITC/GFvX1l5jEkIW9QvrsQBsshT
x1P1Y5zL2DIDEsTi2wJXcZhz+pXIOaXJ9HktSAsLglLQUIIIdgJYujAzd7HqMbV6
k10Z+SGvpEgMxV8n2rjLPWOPeZx0SNZVT+Y/eWmuFtveKpnyvB2PfbjcrL70I/xj
lKPaI+9GfPCpNI/SBjmx6TxvkSCUNk1nNe6MqfUv1By6Kf4cLKT/b7tkj8t05CHa
8FmiZdEZp55OjsTC2KBsAIH5DV4f2tAWD/msU1dVVKA5ZTlnTjzk3y78UL3p4p9a
etsHAKydymoqFw+8IX7VKUmSvVCECmBGV5aZHFN+bGCVKXm4GBM9KaF2kvLU47qf
LIHcnpubWNC4b63nce9GtAel3X/pCE04AtzgQr1Bcu457r7L4vfDexW9LuZ5iI2w
/CpE7HWGz3x3mdSGEG6fNdOtzKgBlB/hamAjkqDQMONgXk1KD37de+D2koS60NTi
tW16dSGIm6yPJomfflMZrgY8UG7cpgz4HMaTCi90nV/CZ/MODIlEHZsNnOsQgazC
EOQ8kW0LWJzsyj2kQZ9kE/yQBuchQkmP3+O9hqjLrmU4mr7T1tZ9Vc67C4BxjQH8
mB0FQbfc7EB0aIfiyvjLUJRhvh/ZzvneYRk/ELn9oFoLVxPu2lvgKbytRTDU941Q
n0MMMRbbp3ETxTTONgqiP7rMdDcHZ7qB3MafjB4g53V1u/9WGrPSnPSqDiTg+O0S
I7CLdP6Cbu1ejZlUZFM6Zjgwjzv543CsmTtOHQngA+L4DdoYKbps0KvLqS6r0WVH
byRJGmzFVoS1IwEcp5Kq8RzO3QZrZWBg327CL+iOqGLO+w0jRah8Yv5CdgHUosf/
QWLWO7geJzgF8w9w+Ku4RVs1F5p8miELTvkshTZAO6Qvdquchtdg9dFeXbgd3dt2
hY85DmLzk2IoNt4IaLT5/e/RjjbM/iq320CofJldXg5dZJKxMpdwff9Uy3cz2HZY
7+bF02VN76aXS7A04h9nPzPD4D1bZUev8obgWXBh/OCRuBvukCr2w7xrLc54znaj
OPoGWTCRVPZjIeC8OURaZL0LPNmgNZcSSiyznSmeCay8luLvybFSW4KYWSIYznxN
N6mf9rIoW+BoBk1DQHnky+6CahuhfM6sJcrMJdWUTZ3C++IhroWHeQIBA8711xdV
rVvU8HdHy79wvsNPEOOJBFxZLDZzdAuLahq6HiV0OHMlmzwP5oBOVBv8pWQmJEc3
7kHiWdHCsiFPBm5NXb6IXjRSzqsjKW6+Z5HRffNNLSzUglwnYntys9VbXeesy17L
uMRUqH+1L3cR7dDx74OF+HWRrKkFOEt7kxtsjAk8FxgNvtFfMAQLiIEyDjOP9mLh
CXmtV22mKbfIlZdo7hYqygS2On1vjQ8deL58NCGGnojWmUsLaJe195lLDtg2vpW4
KyzmNacmn+hp/NCnqFw5F7bAg0LdC1xpHu4ASOP0zE08eR0Slrk6U1gp89PL3qtt
r9ap8qCpzxZmbUbRusFVlXdtnfmg4f3FF2kNdAO+2Rm4YPUlGvNjw/39es906idE
fO9eVDaPhe5zoLrb6tuWZNa8Ck6WmZjvcTJfhN8AZcXedl2SJh9FFCSiSN8mDHWI
FORP4HdD29SNqKlQk63uA8x2QsFJSmrQH6yvM7NLju4q6VqPeJr4qm9U9aFjbMom
+h7S0B7LZ6lhGzCixW6cFCmIZ/jfZGzI24tHvxRdcVcg97qrrQIprvuQXh2WC/ZW
QIey0fBNwiBougINHGWu6asAi42hHGA8iks2/cqbpxJZIqX0kUD7SPVnEct5hG15
4wludvSTcz9lfYaoS4y1U/EgtcvwvDBhNslfaP9ejD8g1/x14oJJvqEHnbBaQZQP
2nFfdN5/gVCgCmGSkxunJOXlClDQSASp1wOhDt3QkmFlyb+P921q52GZLxHiqvvZ
yqE5IC8Qcp6PW5Ki3P9jsv6iGrj4U2IOA6CexqCHRqu48tP+mhToCOoL5oQpcAhv
1gHu6SH6p/cb+MRvA6SzoZ+egPYQshgPj1C52bnVbF/psKY3NQXI4BmcjOi0nlcs
uKzxRtAqF7LlSV/w4vvNJvtxfmO9LS8wSa+X3ajrnExh0uGeN/dqdqlfdfUGcEjm
ZbjnU0OPghqKBeEmDyeNM8pNAs89m1D3Ctq/hBbOKk/G5ci6cQU8dNuAVtsU4Q3W
O+3XPdEb9fi8xF1Km03MsY6+hT5rCkLsmlLL1Rs7GReu/igpFL8QSO8p46/7CNtB
AXf7d45DXa486+DODDSpcZeTVfw3nCK2aghyFs5H1sB1KlIgXsupNaoc8mU2iVbo
/CYeLC8D+2Tahr53Lz4+DPPAexSSTF/ut9VKdDGpZUQQOC4s0I4SkfZIij0s1OoH
kfvhOyGd1G6cA75R1UvMOIyLZPKXCzKLg8u0S3ogX6r8qygfEH9Yio2IDDV9mOR4
v9iLEP04Ag62eqUEt8ih2xJWxVd7VP5XCSEzKGKpPgDgUbGtZsZbecERmmQUnv58
obTVfu6letjP0PbjGlfkppkhNYnhRSCsfXp1IKBMzEfE8bF9gxZNjfARI6b1iHJR
QmW/XYomeBphE0HTWHOb7LUhSh8YIIvHpMJX92GsiWR9qieiAuSWFg7F+htOMr5G
mL8vFZmzYCJLzYWxglmPrxhaskFBSLRPtuQ1XRB/1kdNWfwMrxw+vuIXFl2BDCRd
kW/7/MYML/GghcuWQg/V5CLiUFi6E6KquH8ut537Aoi8oHwo9luYC6Eygu8uX115
msToagfnG6UGnx3DbajBOFyext4pPo5X9i5w2tGqcZoXU+6iXgSsI3YeEL0GRE+r
Jt6tlhAZjo7165BkyMsqOBn6G96fzPQ/XKBCy5JFBYAFlhjXTvDKXJXAkXS6ccDf
KF0UNygoeqUvTU1scM9kUteFqjT6aGQJix8UEHGXWitnGcnLHBRSKdze3vwwJGoS
BogJnkWfbqMJnr3JqJ2Ph1LBVPcylL311wKM4Eq+VJpEOOf5vYTasslxG0Qpsr5Y
srL6xxzI8BfUPGLAPMzGHnB6/QnK9eR+up66KT1z14cXGwEpYQykAQ7hrhdhbcKw
dArizas8xGowiBQOZFUVmzIcinjpSNN9PPSF36tg+MHWeAbXcbT+9PbZqQxo14y0
tr44nGZtiksJoE66vhV00FriFvrWiI3/NF0FAgsM6tlQIDQPkn6Y9OHUf6IQK8JM
FiZCrVloS9O5SOKcj0VQZIjHnxhII9IapdEFPA2NmMOnW3+aHl2wOxrMawuun/MY
UzzBID/+Gy6qgJVVVu0CFn/QeRFJ8sjEA0gnbIjgaWHlSuSFfR1juwLC+AfZCRQO
Vv59dtgfdCzeXa02kxXtwwy9HTZYJXH07Mp5geRjIXLFFbqIktQd9b2dxUBlkjtp
Y6y9fbhOT88s0hZ13g+DRBdYQo2SrWFXGi45XXIn5m7wXwmiFt43CX8IkNtHJ229
kS2/8Ca2/H55+bYeyR1kEM1fch5qNhdQF1DVNF6m80YLDDZTYdU3R84X2HyJMpIa
ypMN9YKYuFkLA9c6dD19O3rT55Ol7juvVT1MDNlOmNqVhfRZ4AYeNV5eg70segis
d7jPJ/Mp8uO4vyDnYrjHA2upWOd73Y3w4xU0MJKMTrWi3L10yHUtvadm7eeCtz5f
BROxq6gbCPmkQNg9NYvGc5a3FkEkCjue8LbmS9fOu9s0p2eOAHUAI4FrS5aDoTlZ
60k9YicSvqBEXcYT/co4EcE5F+CSN4HqMw+RDotzgDJ7TJNDrelirPupXm6lLjPt
njRpWyY7pnqbe5s8ub+O1+2U0P1rpdq+cMQPKGCPGBT6OuYsJpsc6qm/kwxkjj3S
DJII6jVu7928cR619H9RUIJ8/+eNeZk58wsPt+K7nH42JQMjR0Tl8/LJ0GLusvx+
ogDhaRQLIMzE0e+h/Hyps3gZCkTqTxYQSyurVnnPYkB5iUBbXdcIRw77Ef6uyRV3
m/ej6NzALsU8hVkf5RSm/DFOd0pccCiyPxJFfd1FAnyc6045d+3fp60wFhwOLJG6
DEHdaWnfUFgKU2oqJQ7M9kC66HCzhERw2NADpeFMSfezx8Z60Hpa2GrtdmrxG1dj
u/GYj2+GZ7lz1pZTDp/Xxj7Kh+fI0UIpFruknyJyfZKGvP4140Ta/yPMVIqpm5Mx
NPRukF8JnvMPuZroKPmw3XnUb6oCK1mM46MhX1zyHeMYZ0EV2sRl2ceogWvzkjyi
j7uelnjKrxkKxoi590PhGv7bti65dkqjQnetSXTXoWY7fu+FytXL28u0yy7KaplE
b+l0vyWaiD//MqWIjXEQeC4QE1qKN49AeUuHDJIyaXbNRCfBAbAFz97AfS3kuIJ1
oykgKYzawsA+CkrIqN5LJxI/q4T4IMO9YapE7A+qPrLwXeTEDNaKmRqHmeEY+FV0
2g2J869XILudDK7xsh+REkOZi5ToKi/7fYx2DSlthYbc7PYFR7tzXMw2aW/wtftI
J8vnFAhJh2Ff6cAu8LiTIehei21yFyx2XZjT19kVXDUMQAlyHe4EdbcoV3kv6fQr
r9ITwpi419Y/nht5ZyWs4wiBPQ+DM9N2V+MuzsSi1gTgH4H0Vlhf/wLlflzlo2rN
djkHhw5o6QaRrgK5wix/jDtis/Ltf5HI1bL+4es9yIEsLJO34HIttWdQEK/Rgy8R
BkZH5shZBwMcCRC9375L/kDTvTAsU1flsj+h/Jmef+lVUG4f1fjDsnvV7giSrEZl
0ASDACIeZ13dt0R6zVOOIYCW+WcZxxDXWLQUAOv92lwcaxJBXdyT+C32vU8/C5qx
f64WNizyz3HxrxdCREw5SIbm6PSQ1ehtseo15u5TQPHhHdgnPRPKgYnz0s/FBSTn
ILecrnsgr2puM5dvT0OqKiKlTIhttAua7WDxyWS28XiTuJo5ekOexv0DH1rfGnR2
GL5ghrOLt9605BbRTWrXkDCgsgxtVIAfW/NxQMDRbJ7ryVIsZD4tYEnwwp3qgvt3
sLIBa0j8uWXL2oEnIS8aklftXYM24L9P22carlXy7myI4+uuAyQ+VsRvR5ryolcZ
bp9t8wfs3xi7oFrLbvNEEy2x+XdhEGsgJyIkLjCCcYSdrXRF+HP6TlUS9b29IKXV
lX40o+lvONBkKHYRp9vpKV9x0y41PbrJTjtCA8VKZ2j76Yp9dwni77+bdzEVZIiQ
yw7uhqBjmpenZEhWBgaYLpkb8eW/S9D8Wgp7fzYbJZLHJgwym0XSyLeDmQuyapi9
o3TD83M4uX6iLUrkPVY9QKXSIkvw6fs/khzEeEEoOrtXqp1xbK6im4CbZVoxqR1O
r/LDB7Lu4fVRvafzyG1GJfARpT5lVgSr7z8X+0f1eqHuDyQiXBy+fHOh/xfge8XU
NeTRcAzM6f/VNSaBhaIKh45N9Cd852I64b9lOMVdGAcdlndrJmj5I087cts/DdbM
EFZkiUSDW+w9bIk04NhVakK5BdhBVvCtjU5EA445YE3VghKPqpkf9wT/0F4Fv+Ly
lUHMMvivPnLlNEbA36EpHOY25Xn78CHMHifLoo3XN1nb+FuHkBr6eLbPtH1BJHro
jIb6UpGQJO1yFm/O8ttGsrtwwdUgBmzXRbXE6+1mspTrZGj0dwEzXCs/oGocK0Xq
cDecqn4gQNXIJi64wh7otgNq+XC3IMIl1ouLI8s2pwz9T+71+YGROJuB8/N6K13Y
rIbLOxroVcA8TlDDFPfEwbDnpo+gkrPa/+zk7VXJeM8kfsKru7f7keHIOV36kLTR
Fd8B6b1Wf2cFPE6banHTsIbOODWj/lsOgR1TJhp6ZS0XenE4tHSvN8sXmr8lVjZY
epIonL03zvOSpy7u5at69JXzEfERgKL0tQUsSTeYPir8lHvYZCdlmqC6fPiz+Zw/
otL+L3psQT8j//9XqYanOIkSF5lzn3TPgY2cPogAWUPT1tc6mxmmXQo4ZC0b5fjN
9AMGwUIoM2zYXsbsAa5NYLWHJB5qyfWJtjBk6Ol7EUqG/gKV+wRjezS0SMsvt6/y
3Op2J6FfQTXpGDJGoqY9c18c7DlX9oUQthJ6en4qDtqclg2F7ijDt8gknCDAdUyA
ai3z3qMOCuWLnsDYNwCxGvnLVO861nDhuZNcNKlVAWrd9/5/vQAlbVtzHR0yXpzN
LOP6zZozmhrkKidlHUov+3Mop2DUrNF1jKB9kIyojpNYnFKSuzfIBwoUYN1Jw4el
irZ4viCbEr5sDAUtRrDhFq2maIzFhYYJ8HTLtV3eMTt8QhlrKKzWIxCNkV+KPf97
6c3Zi0RpNJKEVFmASM52rJJ9XaF2QcaifiI47mXHRG9axb739Am/hzSqET2ZgzgR
qacXXeTZEDtqdie7esC77yOzqyNOKbLSPAE0roFWLJ+HsJDVaZZ42Ox216FeFhwz
eT42tCBb/UgUbA4LqSR7ebhTzsEhEw42qNf8jgxZ1sycUAup8xumI1xVzh8qTvh8
pkiJA5WsWmchZIv5bALS7Fn9WroNRvVgMu8g+fQrI2rIKZADKOamFaort1nMwZ+v
cHNfUCTE1iRUzkhTotHPzh8hOYtSdT4Djbc6PUloynmoi/DH1dyLG5EVunv9ex9Z
h8iJnCeRihUdhe4JYl+YrMzU0CeCshFNOhWze1OX9MkUDP/GDlsUR+YgksE/fN6f
Ol6pW9jiNa611SmwEmMzGFzd/yiVaJoQdcHR3rLFjtzYB27kBlSmQbjC24uHydTW
gOrNLAIek+aXA1qLDce3ziqTRX1nzrvLMIhJeZHKbXE7XvMmVB8m3GHg/2/j5aq/
2mTNJxbdfbRDg55xSFAkFNA6MJ5jrtSNUpQrffSr4eHnz96ZqjsTHHFS+DAo2P+X
jPg80FJq0m/kku6EKnmuy6DwkmNu0Heqil9J63GPt/Y05R3xcfe+D5BdbR1261xz
knClmKJwYH3m3koWup1PAax+ncUui0umz2unxElQGK/i1N2CVDvA2BiSgzDzQ9zK
3h9s+oy6xb6S7JYIzLpePEaJmxGo79ifopjNx9g9S9kq9JAP4JqvMZPNVRxsKfqT
YxiB1hg4GXy9nPrcx9xCmK8twAL9Xw+efhGBsHrgYCUpJDZ/4honhofcJZqsRiSi
8mH4fGHbZhsbcgU3O88AqpeRXzNRDo4fH7g6w+t4G01baVg0P+BOMGsKpB2Ewu7P
AMXVXBB97l4yjmPIsjex3Rgl440QdWv7moceWNURY4H4VxnQZlviPwHjT2MCp/Mo
XVWzWuATjTgblgdJv7X1fTZ1aDUcaDLm8jNPltkHHOwSpCC3dF0eVpBJwIqZ7Tpg
0/NypAGfTiFm/OvB7NmQjuao5X6Yc9Bwo/TIOQAnZq8UgASRPzAgfnvp6L6GUYBk
c0EwF8HRvS9aK9pqey3npGEpmzYihdcHE4niH7qKrXmyJ+pioMCHXbNDbFm6cnbt
SFgnl+Zs0MIxdxAT4heeP+wdFg/mwXok1NMoo7CyFo0N/3kGxMeZ9Y/XWxPZKR3E
9r2c94szUUpanxkfkPnPfD7WVGzg3bRV+3u4dPI5nioQa+4p5u0twyeC3nz+4B8E
y0rxIQ0Ml6SKa53uAnc0pW+tc5ZHdHPhDLvIddkkpz9pwe0syrpwxdHG1J2zdNj4
E5MP9dKYJaopUdL9wCipeTKoBgzN6LWa+lli0d1BZbl89J+XjDfCjmTT9HZ60UgI
g3VNIz/kMgIIs7KEAtYw/CoF+C8bpswCnWFE6SYy1HXQm+zjyh4ym2WOfx88rYcw
tovGoVlBsRl6MJAl7usrAxdBLXrwrE/VMlkpJURWbw+lEwGk51S2IPGnf7aWBGd6
7uKMcfdgEJALNh9zTLrLwD1eNT0z1ok16O8/zDNSf+MB7F6AOVppIzf5HgoyYtfX
/vXFw3GfLFWVwFoaID8cPT+ph/H93XTNiQ7RGauck8F5fd6DT2DGdC6zoIYkgpYJ
N1rflHdHbO1mIj3MrVFrC648qnnlpEH6EHKXF6isqdKL+R9A4n8hlWZN5IVes9k0
d00rmUlF7kYeqQJQI67FqzSRsGxlatR4yI+JpUWvhnSm+Z60Tqveis6eYSGFAq0y
vwhccDMcHqh0Ij9O+viGz5oEMdSMftCB9r4hHAM7p30EkwwhuTd1QjU+qrciRUy+
HYdLW+CfnD0WMwsgJeW+jV/D15d/Oemb2/pkBzaMvspDf2TxFqDELnnL/46mwrmJ
//0aQt86p0SO0lnRPvuUggorlgfVmbXepXBhDi+jQldTKDxaJzXYPyraSnT5++xc
lPPkVezFVxsmw81nHlbJcDdTHNhVvZZ3D76V9c/WYhFuh4bTWvAYPJ9/qGl8Z8dq
5v3mnLrO0I2nPQ7nI9lDMXu/GxRh/P+xpLDO56a2aUIAllNxiHoNizxy2EBwsb21
7OTqEC72uu7oPgaA2KkDY0IR/9sPgok7o/DYuk7jCa/B2XLmoUauKsYwm4ffJWHV
Lyv8p454BmAkui+ef6lZBppt3DW+eB/zANPq06gz9KtOa/1wsw9hphkTvIhoO+3O
9Mc9cyxsNgjhuKYLWGVi8o+o96ivSVROVTQ6bg1gvbDRlkOJWPqBIUtJ2zx/kojJ
P4tRzPAQqCwQ+qItgftQ7vCcv+kvEPJJq2Mw8mWrTQvphaymZ26k6hNFhS69VYMz
3ZYEnsTYJvRA3ZVsvWWi1c7FLX6ioKXMCaBCiMD9O7kA5+HwK80wEO3x+/UMkawc
ST+F4vIaizRBnIP+g5lYBmHmviz9KMg4fWNhksMSE/cAzSx1ewS7GxVEL071xlah
hkM7w02N+491a9dq/cNRlj1R+xMiErovXmP1VXSERYdKdmpM7OC1YNwjJxOYe2F5
Wodel1G1bo8EjemvAvnSwJhP21HoWUvr16wxbClPriY2EzdUb5lj8p/Qx1JWOj4k
UVjY/E1CdhLiCelLQ27A4zeL0EMP+9p2/uRYoPcSlP76yaOxns0xqU11OqUh2t29
HLZFatQYvh0FdkHNPfGHZfkjIw8SjEQj+w7Skha3j2qtXhDMMULQX9aKhl01HuSE
sFJWgaOvwm6a19xwI5kO54FmtnVIB0t9skfG40pVJ8Qt4IxoSfij02esTHtpplJe
qeEbwytClx4U37ybWgrkVbHB1hxXddN6+yBWAHucntcQ+v7g4K4HjfzRS+b7VK39
BdqyWja4YjWtppsm0p/Cy0PsxKNM0o7fY37Zb8s7eAQ3E/ysk/ExpBWEcVAfPGjR
XK5Q9/u3GcvYcHH6B5UGWky8pX6k2KHjizfMDaSFKVqBatf167737ZXfmaoqHFKO
3wPE9SH3o10tHUqkA4OInj/3+JRd/LDxxa7V8UVi4ft1WI9Pa369XsvHbCuurbiL
Vyuv8JEsns3+QGJq9FE4mEXkzGzX0k43OyUgFRNoCwzBX3dWMl7Dij5aA3EfA1/l
CiFJkkcC5N5CZOGZIElcpPCyb9CzWhNq/xmBU9B9/KH9CAFqwsaY/NvXugMhO1xR
G8caFVj+xEYsiuET2A22sm4WkuU0gtR9h3diCgChPXCl6NiY4UOJSmbucZo3/xau
uXV8Qo5pG6HdHiyi+uHDq0A4tLSGxxmDFACPd7XMX+Hh/K/lbtfKESBZbTtqOvAT
ANDNEEtDNqhOmmuevdhY1aCGE9njHk/Gotf+g4Q2zWA8YQsIFVupl9yxQUCF/6TX
wdzQ1THN0DhzI8DMAZNOmVqD6m/nx+hviZOEd5QqUfo8K8RBSfZC+k5/CzmLYhue
H9hTVH+f4h6O1yxQAfyIMkEHfGz6tzHjOgjqhWHO3qHcEiZwQwqSPRn5mpn8YQ9/
iYUgqsODOGtvmeeDZuZFdsUnxdZVLrtAzv5Ik9rBdj5dNZ+pzAIssDutGsQnO7LC
VU0TMKZ8roTtVUJ1gBvFuX4/DIvVDbwosZ9/XGc5oLfJ80pipo1zTDFN95F606nu
mm24vJ7zNxysGazSZTq4wLTwXLvOwrgIpr19SpKbP+WmwiD2clVsYgxmPnq4JTtg
hkf2yBX/f25c5sCneFZf4m9uQR8CEwf/EZgZIwlbAwmym8hE6JvCIAoJ3cYrkYbk
fLiG9RQ0LPBeZ/lSJgNc4S49C1DFuuDZKnLZgUfNZGRAXjzUutPeU8qMBCa7EBob
mo9BLV3xuRtOetPpXoszKEnBMIbyL6vY+BS0UgkIYz1GTT2rKPKTR6evkelaJu6B
RTcssZMXGgIaA5fisQC3yh4CO9lHJhv0PoqtQUVH/UmlW3mIx1X9Qa1Rf2jFB4cy
AU0zftgQx9udutWTwHjkZeTdrOG8sPiTM+CU/W4RmVW8utkFIBJAzJ1uAghaAiXb
PHzVGHMB5K4DQcAA1zhowg5PP1XNTZSWuzqfuD7Js5CH7L9a/hov6A0eWzTDuUuw
FQyVa2i6+e90FiXjN0zpqAC+ep1S5BSdh73Dz2gaBPs48tRj1CsWg64hHGMgqZLP
MPPllfwju3F3kY3QMG/IPjgP3mT58lPhVwd4Tgl60gCcb4nuxytKPMk1wZeAGCBD
ibA9RFtgw0fD+izBTmZBAVXlxw7GLVDQWdsDrI6hp1vZMVmcjVNpLLXLHy9yB21z
fHeOJffADJH2ZhWEC+UaNsokciHx4Lyr8ypTDrSm5tVMPl/mvGAF4S7F6TdeB2qY
OFiJMUV0hCDPanXwwNvn2HXRIxUBJ4p8PX8JwD2Q3rsj+WAVwtxZXMd5+tmXOa6K
KqcEz73wbdDqlQfhDVUS1DAdq9z957UIX1qAw2XYc5MxT8VwrPQ4/k83/ksnPMs2
nfBsEFBsxewBUNLn5nVd5HvKF2WZD1AslhgsB3sn4qUFQA3TARZJhocaeSgWDD14
BovOC+aQm//HkjPgEtohbkOH2XcTw+ZUkKKTDAei7oghGWUg3xgdNwoEHfkrw+OF
xTdfBJ1fmYUaMrwU3eYi9cXZs1fRWLaoyRt3il52t5sStmNRLb4+Iar3GOgB09bL
lEupXCp0fR33pY4md9L8z1Qr3igegq+tKeyTeKeLe2qQJCI1bwdE72exJ/zPsr02
LMqoIIQFshRausBNSM4hMBcll3Tu/hXxdSxLaUlKcQt8MXezVJwbN8apmq5Hd8nr
XAuTSSkWtyzStAd1oD0xf6yQgLgqI3gJo4lsSO2UKEeOz3206CeLnLc7/7QUVwMW
x7c8oLW1dpT7Z28Ab6jfvodTJSMKVi1oBOnBSXAtaxwpMPbrHA3pV4wg0tUrh582
08AUCtiTayf8OkjrdHwUT3xhvnWicZXLSHIXG4fVfmaLhmeSWS9XIlmq6eIEpu8F
P9OQOmZUJSTqn6ur59IfBe32JApnS5Sn678EWwqYd2yOj0Vmjswh0SvquP04zFd7
q8Ag+yYD4bbCPs23cmdJSakfRi+MQeFt9+KSatMPt/+0QgcmmbFdS24Z7Q03ZTPS
4vB4APpM8527JvlahvCDJOQvajdVmZsD1fAn1bRU197IAt53pjykroOEAsh0z/zA
VuXES3/yZ8TOgnthfzCrB8ig2noJ5Be+xd/KEFYmyTSxOJCiqljE+XAtFhVlMAWC
nZVcVkyqnrAccX0Nb77JUmTHK9gdoqXZkHHagUoSHoBFzY8FxQzz1mUZtomrGPRW
VsIDXYdLqmEmBVpP95sDztmHyD64heyEINnDxCqesdzm8JY8E0ERYIHqLtKYaV2b
tqFb0rMNQAx6qSlfFYd7VcPi2gkC7z0JFA7lvq18K1MfEu/xaQC1Fr2rhVDaUoqL
P+drveWUKdEIFVW+r0dYFD+rO+suY/4ALY9PIGXUsR7Sr3ZKcFs1TWeDkil7Q5MC
wQ2fYcrFLoAOLihmp0zZD3mD7dQonmqhgpTEu8zMSWU0P2bR3cVo3eFA7UtlKjub
oOCjjJH33Qk8KCYpL2Qj6AEinB0aKvSiHq5q9pviCBd12jUx3K28zDVi8VQQ8C1c
ekhAKhBGZUXv0WdVQImSrFifF2tOYQOMc1e4Ji4/l90xaxwmmRjVMfYmeRrPQ4Gg
D3Cdx/uexL4Xr7+f7kzvrO8N3AzUQArkjSbASCGI2fF19N9+M49o+Z1iWTJpl1Fe
UK4UEIEpd5YJviA+sQBhYHUSKkzIbFjzFLhZpsn1Ah5Hry+oskmr3szFj43BJjl5
wb7TW72XCt+eC5nN43bHNnaW80mkTdJko4AlvbySxOyql+3uUnZk3IUUh5o+w+lH
hoFIoIOecZ+E7lNqf3NL6WImsRm9pOKYlvEUTbSO+EXkXs3UQZz35b58iJlAMrkb
nLwC4jHImQEk4o7qVm3SVQmk8rYCR5y51SoJF5rhbdnWIrFYznAjIhOYIX095j5v
0/sHp//bsQNqOAOUx5uBzJmslpIqpc6URFWyL+tQ6ZGsfibcLNgUIFyfm3d73r2G
L+8gyfJdEYl9drWc+EdYZKh32fa61ryLAvet35hJOvyH61cYPX20iymD4NSTyB31
3/6IJBGo7HdjNo58xRfz1RGPOcG4+Z7Y30s8koMQx3XFUwOYjenivkyzUUK6ewQj
+/e60pdHxLJeLC42MavHcK5vT1BsOfZgNtTv1oneFcKy/yxhiVvJU1gcPLYucz34
/S/QkodHDat22J0VzJ0bBx7lUMKXgEcQ0XO1MnpYoAZq8Smlos6W7g2URH1OrodB
i2Xc2DCzo7140xy9tUxm7JFfTuJCDOE4E/74sJf2KhQmnhd3ab3LG6co3qUHqLiD
vyt++aYZ4DVFJP8T0fkq+H5WEGNZPxDTy3dNCO/Hy/wD8z98PQzXok9yIZPj8hIn
k71ENOLwZ/8ro3U/8BleVhhZ5P6GteqFzQ9ICQzmqX9b/TlJ2llnyJEVI4rzBMWi
G0TzY3DEObQpH8pF0CnCFKI6wGHdsCSvgIQ9KlhFnNeAdPeOQSZQd5MX6aOs5muQ
lCHq07DWDLMkTCymOSFLP7UjrwJiBC1RsrUAsv/1uhbtZ84IV1Br0vd20ugkUojL
rnsZDz8M+U58c7gyKDyYUQsAyH/7d8tGgXho7ngjOco6N19ifNNjQkg5PO1cxnfG
zeWoVsiRGpT35/gu+yKQfK5T+xQ5TefKe6wpERdjl2UWY2yLdvUX6GG+xCE8ntea
IxV2d6+mDEHDckU2oVegwU44t/mOja44KKlB2FWP/QrUmHMeFWbdlrODVlCkNImv
2iXRQ9Z8Svxu7Ad/AcuJp6zPpP9udd2wfXlrtnFLvy+DFcej9g2sbqf2/HU4ORRt
uKB/PCOkqEPP6A8g4XAPuo2XB5eco0FEoHfKximodMLU/qVgfD/K23+cRvFzbRkf
g2oULHVJFp9JgL+67Y8aZ8UGgq9qIFpoomeW7jt6gLI13fLD5vXIxCH6T+Dhnwjy
7HPQ6f6nM4oMFd3a+ammo588zneZXBfUritamSYFsLtb40cExB3KAs2lI657SeyM
PEQI0KiVp2WLIbWbupHuE+YN1pAJIdyQU8L8gJAG5iRumPICPbmKgbFQXoPyN/GS
x979pPed4g98E/nBNuHcARnrQqRLwiUu72VMsyrLJJhc/+pxRY+drHlox3Xf9TBQ
u0FIMU17eEFBG66j0RY5jOt41u607bde5owGN8xzA2LztGUD9uP1QVS2FEB8ZHY0
73GGVtGLgRb7guzBVs1LKMPzDr+EpYPF8umeR9Bk8BT7X3jRu2ZlzVb65+uNny8Z
TB6DRuzVunr4L3vv4mSqnhK3KTF5x7iDmWrEor7334L+RU/1l+Mth0NPed5l2Sap
fmxM5p3hANeQteEz1jiF8l7svSYombKVP+WXf4XnANK1NU1CupPVY6q9jREXHdDi
zQOfqBOC7SZti6MlipYjAJgHwTgIotR6X7fhSeCTTxLFrDrBIj4B89IZrlxOb9u8
LJRdPCv92MA+h0PplSHt6Gej1wn223JGLvutDCMErQ5pwZWR1tVisk8XnzCJADLj
AH3MHyvDuqFK4C+UiMEyKDLmPGs/bfgqh5/zGKuk748vwrVHv1SBTii6nhh27N8a
BT0KMBZX83GB0ErpWkLjJEjPw+b/9ZkSyVDfeMkczW6jkXQ7UuVP6vCBpgal/raE
SEqasUHldzS52OKLEOtBEPmu0lZLdYkWXE8aoLCISCe0VbKe5Gr88n8FnGXiKEFD
AEwc0ON4hOE2lqjQs8rHo7KdwZedyFs/l9T2NigQH9k3BTl/IA6+UI2eU15gAvYX
L9mRbiYgad9OnPbnjN8hjXMsyQsuP6jzZV0xQTn36SkQSvClrJ3GALaK5Q292qZ8
NS3eLJoZvUWa3qD/xHIeNfPHPYBjyWMIyyeoaK4lZI+TibAD9HE7bUYJ9DqE6EqL
2O10taF+DIWyCOD5BfDqS+5K6abUV9tOGG7RBDt7zKhzzm1vOILH7ruszrl0rwHy
lpBmVPlhf/SblBkVf0DpjZvWeuk0PMkhyP3zox6i/ojIsrQT4U9ljnS/zNuQWrM8
YvBWRpxnt635aQpHU0BT23KuzSh3yuTG3gf7jLdA5uTtOxHy1AjSOObpXJhJNleO
bpF8MfDKHWoGNoY20nxFgRJ5yYB+7DOGXd2+4pcFj/RhHGqH8uo1s0CUYrflVwC1
OiDjsSWARS8nlFoChHX61t3k++Sb8KdXxXqQ0LPLak+6JwPSukE5YKEcUfYtI1nZ
hkxLnpXPt8kR4wGzRtCJBB4RtqnX6jrfwEQlDBcCG+5zeMke633ufBczkmT6NYWj
zt+xiR1/9vAneX6hltK/c5ei29oAp4vkcdna5QsLYinoXQGhEOsyJd/gIW4MWaYA
0ddiUzPeDRyqyTAO7SNnQea+zHdScZc/D+E9QNqhxPklVB2MLMXAM6DqGhRlTeed
DUdxhWQlfss5W7renZJS0N+5GhqCVktneTcydwMa+z97oW5AfWYBF5eqRlHxBFZ7
U9xdpJBkKD7vLRvAbveRGZVcJ5MZmpNbCFhjzGXuDFUwlvoNcebvYJ8IYoPn6e9M
aAVHBJtQCx0Kq3aBEb4FlHKLySNKCHuSmTcCWurwaUXf+8wkVMIOvL5LxM1lc6Gk
7RBTL3XUAjwzmfQ7QQoo4oFT/dQBn5MeaV6j7R3frmOkbs1HZziuBWXmYphzk3WT
KbhDIVWzOWQMTX5pjon5c0bjVsP06/87Zjdsd6nqIf49E7hnR0aE00WY7xY5LvNb
c57t4W9vkMgfJMzYAQ5gg+jJISLX0tf5YoHt76lRU9N+ry2gYUS6WxzgL5/aa5Fu
OjZFwB8wKBuakfrpfEwGdTtxTw3UpWOJlargKa99J9IptHk5OvdaDkRUasUsMg/y
CBpBft6eCIA86ZldehOVXlZf5ihLb6p9rANW3qhUyhJHlTQNSswGybRUGZaUk/rc
s0/SDz+ALR9DePoVLsGZ71N7zEi82o6NJnDHghziQOppmeZkuGgBgtcYWDLjH6e/
ZPFXs2u5UJan6NGi2TNsQgtwE5WPFa0VhdlvW8ByOQckYntEflvEG1jCA8U+16tU
WBM1udtgWcnvpxUJb9yvTBdt+DBfYJBaS8FXYXdMgePyYJxmUbsmW8Dsrsd3vGde
x7xKWc3i5p12qmyZ0jUhgDkFAlOSijUjZ/vjpjjqBi98wUI2clJOws62fj1btXlJ
c5/gGzMzGy9SjEqT9q9XBffUTdyZCGgYPUUMGX5hbEUxH//cRpfq9OyyEyzGEaVh
pvKazYfVNjD8L5f6fxqWfwGB+HaexW/zUvtYrM1uJZm0h0MBl0t65HMzLoySvbhi
OslPstqFCwu9j9evM0iyxIBp9QDaAfCgGrUBiOlbIru2zONvgwFwj4itF46O35Cn
bnoJJ97wz8GeRAt3ktf0JOmzd8boKpgjRZ3IOpyuhTxjgAvnNPo1wZA/T4tnUI37
ro2D0xdLZbsAmxaYv4SNmzxsUs16YmtITtCwKeUnstzhtZGCxC7nGRXKUaCNAUss
ONUYh96n4vL/o9Jn27+gUVgayWT3PFkc1k76o9KnrqheBfsU+Oe/5AIEk3AMT9T/
EWwBoem4+LHpGGY/ke9UFq4TWfq6kyxKudE+JVmo0C8pgGyO1ZadQnpQBQBgdnVe
3GfrJKI9geERZ4FERUn2iTU82ZV9Xdqik9zEkAMSfEkrQBBVUeutrJH0uOgMExDM
bN6oI/h40MTixMTKdsWg8L8FiRPtnMXPEOud2PnsrGiwzVwI6hJnOC8H5IMu9Wy+
jd/IvXzjD0Qoit4BaKCPynOxCaRAqy5tih4GjCWTMlPK4VR0TRCPL726v9xPEN5p
2ekrp8nJU9qw5PfYRA4vwE0EChjzd3kHG2jfUqlzm8cjpqO23JuXO/TW+WHFKxVj
bqM7aZ+SdOe1n8QrQ9AzSKWtrSWIsGoScNqjXiqDG00ss9n9+bE0f8EYFbWybtLE
r8N7YrKngtsZa+X6E+eaD3t/h3sCgeP+yb4LIppvUGEIZ6I2+R9+ST6UQ87diTj9
ZVJbF6tesQnLkory/teW568smqYXmLABY86tW03z1D9oSbWayqQdIQ/QNFj22llS
odagEomMf6gjp7j6dGTym/8oIHz8mB5+Xv+iJ9cn/B5Dr0p+ESVUz1sah9/0SN5s
XJF32rgnlvQ4MXY0RwKVT43COsISm1HFI4nhreFmqSuNj9+8h4qtMrzSv3DDuMqt
5Aa2/A1UJNiKGrFTkQy14NrSkJtD7vJSoXRDqqV4sw6MOBoCwn8rU2nk8/D999is
OygloTuC11lLc2WFkdaw4Sutc8RLDBUXPYL2xM/8hqGsjqnQPJGxeZYW7trZrPHX
HspwSO3H+blpRLK0PvyLChRgfp538+USOqTPZXyrTQSIdFVVOfnXi3XaYJ/XN32L
ZYcDLAkxS3W270ul45wGgJrath0mkfzXg/nQyfNQZbZpLW+qICFz8Q1hQ9yNuGSp
934VScvn/dONaqZo5ca/JHwYADWjiZefIIq3hBKwD0KBkiubUktCxwAuyMGIsmvY
P6oeqYQgVage/aMuHcSV8irfrerRlv3P7UcocJIrkWiV0v3D2qmv2gO/2vwNBc7x
aUTeVj9of1mq6I+P5WfRE3qM5uHT+lZDfAmThTNxuWuDPvqnUGD76fZDa6R8buNo
2SnjtE/KFpe97U1lMNPrjVT1TNUXye9DYh1hXCBcqM5Vh3gN8f6dT8bfyVy1SWvF
RCbidUMUpLjS1dVybYqQoHiY8JKaOHvxp8N9qug/AZAqVgwawINeLn7DvqGRTLHN
VQy35ByH0LbQ+DEAuevWz7KTWdWxLnlR63bn54op4rgb/+bV92Pev4C4qrJv6/To
gz8KPVvOVAe2xofCLe1/h6GFGx0wfuBK6I+ntyvWWfbYGnFF3c/nWxhlVHnCSKHw
9qK5v8b00tNcFsjk0M5RGIXXR7YFDWgsmSGM4Q8E0jCmlIreuOrvSkCc7KNdTe4w
0YIXPUDV8dKOe/1LkWRH60lyYBzl8mSEcYeHWNrICnbhiKAlXtNXwVWQceZeDAqz
BXtD42kRxQUzhIq1ANZEJewXnZJ7XOfY8hXwpdo6wLk0pNc7vzRh+0YGvPNBkd8+
CWlq6m5rfMxrjZa3RuYy5p5vymXdar+zmZPBWPuHtC/OVOnqYNMQlXGm1bXvBgOr
Q6hJ2NbfxaM7M0xjIcollogPZtFIB1cEefeP3gSde90ibxB/5oAnWL2Igf7/OU/U
RHhzUuO6H4CjcP4DIU1DPcdsRILh9evW/BwSkFq7J/h8VUFbNJxr+1M/r/M9X5RU
n+VzMCytf9EmFbSde5ghJiZdQcfmjG2phRsTqlJdEB+A3U1Ews/NwSqSfgiBCbjY
NUXGbE9y+kZoQ3x7jCXLBcQQ1fRNqypvq0+SE9TnE5J0ghpOB2HJOijleO9IZoIB
EMRsNk7NLo72KgCdxt/v57o7uBCk9gWpnEKCDvThy5J5XqDsKGOg7P3Wi5nfcysc
zOk+HO8sXEC0kC0xG/NESgvIz/oZzKdHGtNAZJqE/LKasMkamhmOMHgNuuEnE16e
9mN6KD7/gNX9fevo7KxzkR/xXr2o3nzuplhrZskmfMgtKbI5fty2Zwpxo7FAtqyF
F3RQfQchCBcdpgpX/XsQ0DrPwl5xxhk+ihGIYxUTfA5ZSVwM2ov8YWFZMzn2K0Jl
jc12eaVhEL04HV+bXah1JjyOiYk5MmJL3OlHNdBStSiGxY54Wsaq9Ar6zSsDM4AO
iZp5hWhn16ReIPHVloGjVZ4yJEXSyKBIOAJ8KFq5OX81/2Vfd47FahA4Qt8O30/B
8pX/jtW9+iIOxTU2sJRZZrGPR8+QoaQSUhpC+rDyubKg/CVxSbYDKelI3TAm3HaQ
GiTEXO9i6IPsSzDnwK3qKhi0hT2INnwMrbrhYdG3hA/a8KAYer4NfzyzW9y+Q5dt
otAU25qiiVV/51zn7U8HQNoi/XhG0sedxsOn6yOWjR1yU9kpwWE2lhSTmF5krO77
lT9uObneXprfbTbszNnEQg0FD2lYSxX4gtOZ2+eJ3/KuNS47Ye7UaFEJkIGGPzKh
0Z9RXNgtc2ATn3cPr5jzgkK2iwZJqcF/tCFWgfpY7Ff5dsFcu4hRTwcPHa6QKYe9
G+4Iq275rSrSSSFsnXhtF5dgzBgA6c0KKN2GEWyyp8O188Iczo5E6tbxPiVxtA9i
mSdAGfUY4TMcbbBq8yec9NCqYSyEXtG21YZvgKmtGAN0EW518yTHFvjcQ3ve0QSr
38onQu8gnLCkwp7ydrh39RkRmrNP8XIcHVHi47b8WNQ+v0KANOzKZNG41/3sLrE/
uFuts/2FWbQl+5MBXKdpVyGd/uCr9qKOT5ZHoBsHf6TcwG5ztyRNQcOqLDx28AA9
ohupOMKGrcVDcjcjuEa4JcByGM9bBTEwvURjojgdTPDD3so0+a0F7dH+biipWDX3
GwOYApfVEHuIEVe5W6cgXZI85bWgdDcrEMDxxGpfIrzTcZHa/3D/nucPLG3Xik9W
Pw232mlcDtkO9p14NXKbfpOG7+E91koa/czApTiZzjK2O2lumv1Sl+gGUIwCvBcq
ItSPL6W/MK1MSEdYvAqEpqKNjxo/DLp60//sYPrpm3CuxoI05NNDlbLOjB0E8z32
AAHRa3sohZBk1tfgIbmMxTWL7nAb9jFDr300NCRFT3pLjcwtjvoXUAEOY2FsZCNm
sbehm2E6N6+MlINAYtGA+lDL9ENVovqvw3YQibNYdEvsRREhkPdIRpNMO/teze8a
6tZvjAgE7ZpQmDmJjRU5vAOYJf9s+Z5AShzmARJBCpdJlEf0TEVqnph1QBW5LwyZ
r8LM3g2lAYWdkE8LQkrtTerHCh5gXqIpNiQx/EWthKor9Tp1Gh/a7sQUOkRj8Eg9
uaYMYztLHZnqatt9lztEyjRfmVAHNL3AFm198o7/M5i1xb6T0p0F4nbm7f4gLA11
aUBIBtnHaNPtBIdmuTtvjD3oR1DXUNnYKIkwhkxyLKUUcuQexgatKWShRgn3WfPR
KgAG02gdl0pO0vlzKXJO5dcmLRdi/NDbcNLqqETK/IFWB8dXBtQ3uIJIUbUn7as/
V7kiq2QD6ee8V0vrYKu3uqgKIQN274Cy9OQAd00A8B8igQbNlfG5/IHxo9sdfcjX
mWmvV1loU/261efco8+ibExWyHcvYGiIwA0zU5YeV2PGh7q88bFIQ8Nn/GiMZNyE
PhjXcEHPKBhdEdkPie4ig+/0hL7b7QtBvZmQ7GMu9BMSxNvrsb7Hk4w4g10rfpJG
/sFykam5QwHIZwO4Jo01QuNR63h+Aj0D74ryMADqdAhonkYMz6iOewuVQM9RHZFO
jwSsQntTdH56CQKwY9/HZtvnfpdAeJsFV8LDXhXUe8LYf6cnC2nsznFMKOpqHaME
ZcPxn249uYsQOcsYr9FEce/P5t8wxvW6cVKz12MGnPX7zydDN0fzCgpmOoIRTZ/n
sOBPwlRSD0vP0a7mTr84XIoKw/IB/DQHHqPAqD71Pj2a/YLR4NCAGDMsMnEipL5E
gSPFLnF++VU4VRnLXmO+1mezZYa/+7fmkD041kaWjJjdnNlYBP4bKGctF/2+8lZR
T+kTJpI/jCu/aecDJeo8v51EiSP3NUMrKyjgSXNfS3ZhlwrQw5Uk5x8HEnIYVssk
JQLH8wSyBmvCcRDAFEgrm1hmxd/1UkoDGivHq1O2XLuKtw5YHmk+PmYTglSE+LZx
jQNaL3QA5yh6zHEYbFo+qRQkkshmTBIY5dA4CqL6m13uWd6n0C5R77sXS5lwKXgY
HiO8DxY0eV5F9zN0qvFEmPI4MmZbBc/a2gLZz3f0iHVzWT4xZ5Cgy0fQWTdw2dFn
MGYDvCuVVNsa1nK/h8TCBH0ptW2r5AHZb/0E2LpQR03/EIyYJUouObkQPqtMjEQD
H5opUsH/oDuk9maaRZrM9jivKC5v8N5+SL4ZmP6DwUcx81xcmcIB2Lbt/Q9Tzlpu
fGhEp/mxkwZJkWhMRQYqw2mwARlEI/wcv/RfeRVGSdJHnhmiSHRNQa44NDufpzEp
HrZ//fO/KbPcN3kTHFIlc9E6+zIW2WhjJRln4ooiTKwJMhaSrrJCRCemzqYE29Ly
tlk8V7KiIy6TVtEh5yeXRHrtLFaCisgG85U8leYB9ISeyQJeUdeXyKAbDYVUwvBV
7AgqX3FF2fsP+2vFIpL4v03S+7X3F47mNwNBvPxYChiFchlKzvTTlD306mEKUk5w
Wg2FBx1L5VsH4aYodhaeNiCWiHUhuOvS3lIehyQ8cMuTNKOQRKVxTKDlcby+Ig98
lyFuTGLZrukQkyupVUHQcQMBH+4RIypsAVk4IEQQ16sB+8BFGOZk88TyEx/58V3f
ZLTSnhazoUFBVN/5cx+kw0Nqx8CIPDRL4Z5axePNGaCiJuZvAG6MeA9T7BufXceX
YBfBabNwYR+cyjuUQ/1EydPqagV9EegCQBmtUWD1cfnJSn7evva548NUy0BVoASH
WMQG/kVIoQjypeIlpl4LFkliEmB7O/CIowxtyEa7Cd1KCVnIHRdzT/aAIJtBkMqV
yB9nu63/gZUnvWCVnmnPz2ZOyyaLdjuy3c4AvTLTyu2P7TbyDTlUAkLsEMS3tNbT
kG/oD756q3fGFtb5LmMQ+5WZzJpmHn5fp3PmJyZKuMhF5cHtu/4Q/BMf/48F5TCx
ABNgEpZUBblV/wruSBu1gKrWNM9N14UBjnuhTE1gc6rXLFpvoyFAiCKjqP6kHUMP
WuR2K4NczC2ERhqDUKA4ITUoeKlb7kpyjEF6vC2yVW0ZPSSjw1IsG3yIDFGIkZ6D
GkmN/WwAUhXxH0gnKHzw91pvYwBxO3yL7HGVV6p8FrnYJRCFbPozACtLUGpFLNoy
cPaoJLtc+yneB4pERoDkb7BZTrRx9BKGHCn+sGqSgwFPDB/lbgrpL22o36dEBL4q
nHZMC0SsmGL/070CTkUWRUKnCy3BuNx2z5CzO8phFwmX+sxWWB3Pe8nu3cGau2bX
b0pS2c1Chij/wPNjK1sMTuA5eF2VonKimwLiCRkufHsQOaEeKKaXA2Xgg7OFs9JD
W6sbmwaImyZ47qj6hhshn92rILNDBD53RtEzH/AduQxPc6LGU1QGHbtTEB8La5G1
xZ/oiSyPAu1UdIyisO1QtinLuoBslR+eWLDGCZtQ5l2gy8hsC3mu7HyAThJlBiqX
gLthVCqd5mYoCP3iJgvC08PSG8vapUW+MogYALdMRNfcAMxq7A/S0wde8stCQF3k
ysCL0YFTaWLjmAGq19Wr8OfZf6kkPvhxMXZhbfQ7GtnuYVGgcLdcSP+6K8zq8Oto
K+rocL3H1WRiqWxJuRUSo5zof5bv/0i++mSdif3s8CNWIE2DHK7tNNYzG1CFS1+i
QHajSHyGPCtxlnTm/V6IvOZMX2kqAahuUhQ0jcVSIgxHGbTqRoSmwyXEGWyUY+gT
YQrDySALi3uqSIkkIa9fAaTuq8qhOzGRDrhOldX6O5WFJUi/0ed2QG3Wtk9HL3ve
imtzRPy+rO03koUKfGmyW5iNb6RJIng5NA655L1/fvx+IsBf9u1Mi1gXyH+doSFs
BstEWwgzq8A38/wRksPnzn0prPPasldOTYGcRIkckY+vELHFZyzXW0EJKMt3VUBj
Z+GE1BZqyrHvFahJmlu04FfeiWsds4H3TyGkwripvXpCyzGeIdBFCtLVcALikOAg
X+bboIBUhRBOkgH4TIuKvLSaL2lzSvbwG1YyqpGwPTqloD7dTLL82R31KVIAJkvt
W2/bKq3zccS+X2RwktP35hKUr5Z6l5yOq2h3HIqpL3dQ92xAopALWZqoAncuQqm6
fH9OYdkoGKh+zF6Snx3FvLu9WgG91HjDFBN8R07g8GWDhdMNIgE28HhTJBwOKQtw
7DkapWBywj6C+Mxab5jV7zJQ2VeytDMSBVHBx1Q+GqUN/1INOtHEpdTZ1tJgMrLH
pmBAz+XetGQd82RfxhtU+tTSW/X+rY8kKSdF0unnb9Z9zWl4s4D5Eq/HkAst1jqV
MUl0m8CKnMyQDjgmOIk+GhzXm+VNhM2Za/2htc6A8yofJ5DaFEaHbAtDtdF93PuC
WuQEKidgxyw05AYgxR3LjjrpeALGKOa1BOQQs9e2vKu2KPaAiTxgJ8dgdX7U6nQm
OjnYu41ZNoiQ6pVwKG4S72s9ZBqGSvC5ekW2DDeF5tYT/vLyD5kEKtGXhhRCSGGC
03f/nD0QyN6A70FxM4PdYj0QS8lUVYjX0iQL8aM98ibMi1E3P7mr89CnOEnHH7K8
u51fDpY6jeLkyMWjzTTW+S+3WHuoka0Wzc2PolctP3hH6w7kPZHF8ydk30vIMNre
JPA7qAxO69pkMWs89W89wKt7vxXrgLIvxWF1y4FVF1EpbQK5jot6TTXduIKSifcE
eGgKLMsp8IprIjuJMRSZG32NmmLMNgQl14Fdxwx80+udy3qfVWJi52lIrlsWaWnk
MGxAqBDV3rlKw5rXAHufck9T0U0MrjDz2AlmGoVDbS7PiABzf5RcScGd2CZEwDel
+mY8zGC/YTGipnLMyFx21a7cf6ro/TjyyHJQ6/Oyf5+PggzY2NPjOJPn97daOEJe
Ui2voHCshSmqxlZJXHKX3FQSLgd8+nvgVAW76qDS+C9j5A0BVXQf+NBk5ONodVKX
GOgaH3Oqo81K2oTsBt4mziWWaWXiHnjUbR7jnjyI+iHw+Q8S/SEc/wBFKuCCTKaG
IkQkoKk6/VwfBudSeEZK5IjYFparDmyCMQVMjUv/3W5+4HmYIndo5ZIev2g1JxHZ
5bm+33vstdm0rLKmen5bTVfwGct0DA9U+tJr8AJaIoom3dGR+zkurxYzwJbwzbgv
aK2BEULTtfm/xWECZPZJf/UcFUoQpuy9a3n4V7uCNuo5MRuulr19WmGAy/hNQsK0
A2K8zhNdulw6SSbwpjdDreVg8F71kEYbHqxzhIOTpngZVfQIAnKB+rCxZGj4uP+H
A74oCbic/5New4kWogcoUEKuAS4sc6AESR7jjGjoTy5aJ8DLgNRpPumqdk7RBbkq
ZiwLN7F0pgNnQZMfqPi8bzE2rV0dGvLGoGuxmny797eoK6r3QfEOZVQ0da4BLLCw
iFBTfqfgYyb+SpFQMv5SzfnmWQl5PFYWgD2j/ItXzKBJFjGVPX5CocudRdsq/mO0
YCLK3mU+9/68HvO6a9UfSqmhXEnZvqItbPSScGrtT7pRmKnL6z33wK1uD//dUG+I
neeRowGXeHOZO1+xIHZ0htFd37vS+nv7KjumHdRV/D3/5dpBrgevJnfIpIvF+XQT
yHDgesMKqr8T8sGv8bPwJwn6hW54SV7Wj63Y+PcPap7lsyiDYvJQkro2G/AZn6J/
Y7Qg3VZwNlasi5DGUOpMI3CdD7asnXJsSB5IzHQOg5pAjkgliMl/2ogV3cFmLXaS
Uy/mmVDhd37DAZo0B2dHpPsS95mFmrGK9m8jej8ewnS6qej0LVjw0nTHyzSl+ZB8
k6+psfCE0d5hF2fR8g4p4LNWvYYkANYPyWZ4qyUEwYLi8a/F7rxpCVOcDZjtTbG6
fBhe3IIyz6JjPkm4EM4X47bueY2+hshkDOASkeKHsWYpCxCSues/bi4tl74y+mmr
udlHb/vb9UV+qrUdL31W3GC+fHJ/6So+IdumKcXXjiCan2+uwKktgNIDrJDWy4Kp
xsq+E2cG5u65QnHcNRx3BomAMYHbINrDtACprpMCuE+ZV11xYNxdbQWxzlRstJ1D
Kpv6sliEzW083AxBJEoGdtBIucupcJ95YxFF/YJ83Rfx5PlbMlCYEXeShX3tsdPN
d/g0YqpmZfuyd0yqL/vhUiu3Yr+/FUhcGGYo5WEJV1EF5zpuQ6LybY1g4VCNDJvF
CidOv2xXJvPTeIL03DmEclQGzX6rDfWz9Iqykxi3V63u3L1SzVWWrryOZHE8/zPl
TiZmwe70c44AHAnG/l7YGsHtyo1AR5bNth7Ba0+kWCD9AXgCzpbfOBzLgl+PzgBC
SrH1iSrhZwESnl24uFEIdq3f1UUKS7RD4hL6lFH0peyMkQroBDGLEEQOLlzP9aWF
3jEYIBZcyGO+z0P+2z2irnyBl49MAj9FbqWl8hY6QAcvN/pOcMKfUTTwdP+aa7ce
/hYfKSH0Ngu9BmY1dY3PzZ6IrdzSmbfnsamx+YuU7efcajd3npgJjmx8Ko3h16ar
jSVQ+jsogEDmPJfGsh4BCVJzUHwOFiTdmP1bJTtG3bOQpjv5JybEog1zz+Cb3UcS
Ed+/LvKnHhfkn/J6qKgQMw9RbCjLQf/Fo90SfQ7NOeoFJ/rLNSqtW0YLjEgWpmEZ
WbsApFC9ALhz6ATeX/Yl2UJv24M1aZYM1w2Y9UIqAMJLWWe0fba+nE3rzXvENuHF
1bqbc8AhCzVcAaaiPb5KOLlWnFnIa5buGLgB74z1QVCTX5SsxrH7a7vQ1zZe3sxu
hv/vu1/lo60aNpLonWPs2mrhYlVftDH7EfWz5OVIcBiE9Jp0JpuvlCzOxL1G2J7n
KKtT9BmraC/6sHs1oLIXMtHFpypf2RXtbAcIMX0Y4eoNFGLJJIKqxH4yAHE9jf/T
lsfEIZ3tvhB3uoE6UhhXA6LJbUYfKF77bGbntCbu1THWGUbCtD/1EYnyytppZkw5
emSL5m38tlF7Xj5pmK1gNd0Ik2RN/Lz5sQ+pzsRYbWTav4AkZWi83f2q61bQivoy
oi1D6xArtaHlhbhUnQW4r4IbQNHvK+VXQJ9aSV660FhzYtJAXSZ+aTT6OkJUNKcM
QQC2fLKY8PTXuUMMhgSHI4u7CJGqTTjh5mHaYfQ/JbKNZ4JUCZYbMJ+Y3RMRwxdc
a7x3Nrv+xjO0mab6XKgDCETmodTiRzYuQW5YO/UtcmvGydTv0yVi1ydEBX/1ulbC
gLV2IbCTC6ZUBceZMHRkZ0HgVfBAfuvU/YdOcwHhAlOAfmtlVYQ9xcp9gnWC+0MN
qgCaB3VfuXL424TzB381QAA1jXMxhXyj8AE85AUHKNhD4uJ4mHSTppwBWSryG9r1
ZAPrTRDRpbfKSDQjuYxl+QN3d8e3u2K34m30KGJiR8KB0O3CUg5yxanRnkRSTTrB
ITKYFWHGgzUDW+v7AjBT4q1Pbjj4lMcxHsA49YS1KpHhLCiukTE93SJZj9yhnmlq
z+OgWlXsgDOT6HOLBxvcOm1aNKGs+DnVWFtN4wGZLojygLeVwLB20IEJw+5yOofa
KTbnHT0vfr81fzo8TUrc0BcWk8y0B9j4bYFuytuyXqMbFw3dp2xDwLohG4jfuPor
locETdxDdXjzfPGfE+9BkzSCJlc7g+C1IN7vKbOfbvQgm0IKKm+F+ywALJ2lQIwv
CDUoF+QRnOP4AOqjoFFtjDdhPbyO5OAdOEjQS6OhCZITuzWDyBsT/iZim+2ezWTo
TjrkZxHJaNBIWrVeFAK+jE3Tsle8bUTwFd1LUEiRUuLINCxllpkU55DbNWx7X1gM
H6bI9T3nOiPPthcbVu48IoCbZlZoYwk0b+jEoS/Qy9FNaDd2pLQ/4RvsbWmZVe8Q
9SqU6RaJyNdExXgeZvPwygSVJrmvISbvfJ1QIXBEZqLKBRuRfpN/iE/ORAaOlqPR
FI3lnweRPKLzKiOFZM0gDo1ojqcV3OgOXtj3144JbPCcf4rx8D+adj6onnRAOjDV
IfLVk0HL2BZsHAauv+ZriLBLgSTFidj/JqkGtJOHH1kzhl2nHf/GVxbk1QbZNjD7
udr3PBpOs5QDzqN2xid+DjKj9DMSEXuprkrUqlGp/7wDc6MF5cHizRoHCq3MdV9w
aklExtE230ARaULvetHFtZ2MOrQe7ih6Ycwbo1TFQbQX0SYTk2ixJwq4wrOXQI0F
Jh8L61GVzmlQKCYEfg3ADL/JSw0RjcPRHJlReLmUsk8B3hFhnXRpqfq28Wfr+Ggl
jCq+SzCQ7/EaYM1HoFLmB+UbylciEeDFzz28HErEz+nFZP8VuMqPATCjX5Eyp+VL
wM/I30h1i6mFQZ2b+xnrT7v5XgIk4Ap0uFqC+H/pul0WK5h4qwBTH8wtco1uFNin
j8T0SThtEGmUnYFZmCSGwqHH2/jxmetgvF9mWYIzsYfz7SZJmvsYsTfl9BExAti5
LKRyGAq0AVAKP4+8WIDH8PQapgAyBZ6TMiHcGdIRNsezFG3Ha5rufDbL1OaYczji
t9BjtfjtGvdePGicDvg+1fi6jiZu+HpWEHVNwgSWQLp7h+z7CAyT9pwg6mOdRu8Q
LHLh/X/rw9aw8ku3ncuyM/Uj2eR43pEhgC425VvQx2zLvb7mXXWDiZioce19mbH3
S2KC/JtM3W5jgDLzdl0LhxFVWpIiYD5rXpumDo++W/CtxE8qmLGnjtNN63RWXtu8
A1fdtOHJmDeuqjlmSK2z2tvLxBC58nN3FbMiZPMvWDkNAjOozYuH3RCVaiRKMv/a
/F3XAZwZ+otB270jcT3Y0Jmzngr3j4kHKrPJATaGSTa2D77J/T7z2cvDJleSv2Nl
fMmO/uXw8latkgnNHAQsq8dPmuvnhcB3Kucdoueeyjcq2TZ/s2x2R1bZxhPHmzDc
teCLpzI3XZSlcJj0eYBbqWJnAerKkv4TBaQltAHTcjC4EnxPGw/zib5Pl9FKCDNc
zqbfFg015eC21wOig2YAIJR0UqfGSp1wtdu87Hz+cUBpv49GpjjBFSRInp6j9ml1
MyIQNhtBB9KocdOdQSmvqr6d9LYdgAGKcnWRL+z15Ywe0J7OKX9QmKvlV7U7V7BQ
igALLFIJrMYOTY38+Cf1jhgC8Ea2Mvw4i3t2LfQSJ6nE44+Ie1WHZMS+Mlv1KDWz
HiW0ssMJcpxNIc0wibt3qJA+Nc8QHjJsZLqw++/6YQ6JBtBNbTH1U+EFbpqwCe4C
Hp5w6zscqsQ95K+AB+u66wb8UqIr/G1340sDI6A21DU/TvTnDvXmMphq+45eJwO5
2hlHxDBf25rdQTLVOZv98CJ4VdUjw9GVxhf/XynhSeQV0urSi6rCY5fgwRS2fi4R
bFJBdEF1U4/ZRJKBc+2z/VWhxlEWVqmG9MhUZLClJG1HyK2z+vcER8X94miqjjD2
RBTfiMoRgffJ9hcZvnmLq74OrJgjT6cRvBrTQTVtmIsqcieywBn392SZXXsv1N1i
ixf3rm7wENhk3UDaFNjCSISXH3JWHzrjb1IksCW+51rHO5+dUe9ht197hXqgRAsa
qE8pt1I0sLNibiI62tCfVV41mYVbFi43VKuR/Aw7LWk41ljT6xsJ1ggjE1eaj0D2
Q93/eCVRTp9Xac1xO1a618tLgo1L+l4bFBmn4OynP2znv85u34rp3YTuObO7bP3a
MuV16/uB1tTgovFaC2HDmjdDWwiWp1xK0L9t/uIShgWBvomsOoZp4P2ki5Reg0nq
iO4JZF4yroZdenQsG94fFBBShkilFTkDej6yFHeE5/XP8GRPZz5v7mcasC5Bcxr/
ZOYRYdwD5j5a9Z8bo9WCUdID0DFaVVC62a8SzJhikn7EcEY//unHsxXwpcO7Y4Y3
5TER/YdszV++547lGsq2x5AnXK5BNgRd+DEp0SlzibeRmQIzPSbt2nitOadFwhR5
1NhNj2uPKH/7uo6N4INP6hIVjrg8z5Q4b8oUhf6rv4Ny3r4MEVy/NDduQ9t9jA7f
TslrIerhBic68sPDFf+8Jaze0dKIEJjuC0lxenXBlc+rdV5z9q8uB/QrGRgHZ03q
21aGzXe1sEVp2H4NM+KAK6c08cX+97Cme3XgnFgcU/WuoQs186lmavhHc8w3sj1X
Er5nfv/FUU60BfFGdzTVF5Y0nltxQyVtwBltZcAUDqH1pmD0zasIiZwYiBhzOTNS
itVsGFte0pwEAoyYDZWsmCFZPm0ldwUw0LPDPaIzdWavF5TpDPS01haXaufJmJGX
LI4f913FsR8kl9OS5Y6cEgqP2i8bvud3+nyxnl7gwZ3fsU33cv8d/DbUCXMKfqsx
v4odb7gzhnv3LsQpr/pQJ+/n5beERFY5YJ7eLL8em4Xs+dWwEGgJFW2vWP7MMIbC
Y0oPEnkdY09sTQRYjj1T/IR8JeWsDgsD3jQ1Pni/mNQFluSKSTy/sns0ybnqlTqd
YFH/2eQyDKToUIyHIBJnyT1JxJaUQ9R93yvQ1CsetbwPWaoniL0w3tx6c+2mc1JY
P0gJtY9QWcunwT3LxATzCGqzgAvW9ZUZRoYPvUIDwyPXsynDZJu+ZGWNK9suwLxU
hErsm6sNkN2I/DukHz8nUXxH74K5LPLV8Kv4bC3Jk7FTuKKEFTVq2B+0oe5BUk2a
wrAz9XC3i9MM0eTnQxCwz+Ovsa6tFJv+IQOSDdNYgH0SYExDp1LrzKTlOMiMJ2aT
Rwo5uLfstD+9YHJMemTFlXjBh7QvlMIMgZ00v2mx1GyT46x3vAd1y2NtqraQQ1fU
tTr09dlpua9+iBCPW+RXlsMmPIOze3yO/mhUj1el2FbhLdIvN9n98hfMoDf3d/SZ
JDaANgcq99L1tB9sM5glgm5DORoHVKXWJT4ip267nqb3vgDSFSdjdloViQPeyt4Q
KSPUFlNScGDzxEOJjR/K1P1qtPxjmwHxAGHH1EQghq7uWLz6QdlTOZ3C3nQoj4Ek
wE8ggPcbmCANY18rvEa/xQaO3b7AnDWrmml9ZTBmAFGwm8bTvcmu6gl0Xnkn8LJl
LTIglbMS+zhA5YyLd9sShyk+gA2pajXRTdEGLSbwayU3lmDdMfzhiziLYc+fvh17
6/lqWTYaw1lYlzIlxX3iq0UQ/Eqy7CQoJFoa8j7zs+oj0udJsozB4oyZPHLFelt+
CqUwqrIAmT8ozcyO28FM+F+7I6a3uY7nB3gKJ9wW6uqaEjFIo8lx/uxL+Ln1Dz7m
OwMoUoTBCCahbNzt9TJoLabxyFmJlck5r0iEHKoD+L2Uevepgeldlnqjn8xDJ0pb
DWtVzId7qZedaQS6CUXckWSzULKWZBe1NJ+dMunkvlfwJqIdaIkOuCxOg/syu0Ba
2D6v7xDakPICMIxwXC9IuD2EZigeJ79tn/SQb0Qn7aT8lBMb6QR5myqDLxdA3aEq
UE7bF5QQZ+cs1xMHN55a9LfxTMe6Fp0fMmMtGxnuy+frSVTF/g3V7aqwwWyOX0bT
9oiKqY+vYjYVPElAlXUKCBKAR3dn4xNbGwVN/uG4r85JXYdTXQf0Vl1ZIqPMUb+J
aGzEzayzdJRdzifYgt/cUW8cxF9q0MVtAccDDOSMWpa7/9UhCPQ2K0J15s61wexk
TxRKrCwQDJvwHsJ+jVK7qN0txAgXV/npf1XY+3eyX/pBYqXrk1TPZIeH1BxpG0z4
rWiNBIHyxwpEX68/u1eJ0H/c8kyTlOMjIxNDbNYItSxq9Z6ysNn7Hl7gHCeLL6S2
agHixdJERQ2NgiO2xO41JJm1uKHDpdnBG0SrRTNg/M8HTKEzXEjRdN6O3izcrew9
WJNKczB0BVoe4ULDvjXnDKrFEV8fA0w11iKelfYVMYutyYqZkZUT7O/ZkG4Q3DQr
GU6Bruwh96+SDfGfRZcCx8Hd9UpwMxYhy9SmiKQa5qAO5MZV3n85QFS5r5fXVZdR
fQAdnWda4Zhb4dnGu4QO90EBikTjR7LK71xdMyTBW9rjzjXdhfGzxhLO7uEDgO0M
CiY7+nzoJbteWYySEomEJhQLZmiCFGTQJQPV7L5CwoG0edMjt19LImucPFOqzrII
nP6Ogg7CsKfy8dVmNs5oP+iq2jvWjIlVBdzMNdLNLkXI5pVNDKCesAOo4DDtPf+J
Sn2uMplhlfDT6eOqA4QH0o/AFPeHKGSVoyD/u/huBRBEPYjOTbZ1DNjwaN6F/3cm
c2PDwzuu1A348fL/OWE3zw+Qe0xJ3gKciN18owyneN+/VVer4SyVFhEOTOUYx9zK
uUpIm6DsPTb6WOIEnHNiQ7X02I9a0qY3MW203TYr6uUL8N1ZI8IfkKfpNAz/K25T
sbAG1wrGeD26nVf7lZiJRJCWq8SElEH2luGMzljbllYWWcWoGZlrOJzIfNF56ysi
1mDa+IXDDbTtYtaDDJhhEUbvvjkVI/H3MB54d00K1A6IQD+sq2zGxUgro+oIpzwf
iGhb+EJ/1uGk4HEx94xBYxae5s13vpm5RP0XlryPA88i6eWXqBa+jAIOWylpdoJk
O262UAX73Qg9Fc9UYTi/sLLQHs1q/uC0gbfYTJueVSs8b5d7Y8h2EBf3v+mzYYtu
n7TYG60XfbZp3WzUTXj53ePC8EsMJrYVSulyOEoAj5rXzaVZE2pQv8w1HPHA1N/O
qqP13Y8/h2geyu9coD2PE6eQ+pOCY9+sIIiP+d1a46VuClb1UrH+fgp+Qu1iA9HS
Is3RlQ6PkNJuNjEF8CFhzbUNDT4fN1lspraTBGnpGvdx6wK4F8iiFf0IEGlUEFIF
SDZ8se/nFebLg8cWc/1YzZXlzyeqlmamuJB57KRzBp0QsOkvbWLqtxx5NIdhrprq
1WshTTmnnwCAtRHfHITXa9yseBaipKayT1CvV+vtSNeFPbsvFfnJqWtdAMZjIRAC
iGCgbTKWhSAuDfUgKYtaCnSNNZT78v2Hs+WQv+Xqg3cjrM9DoF9jfaB6GWT5+0SW
qwRjzPXmRZo8D3uy8FUJP9uZgfgEj9OxeNUQTu9nCd5YTmm8EtjqTBDU4yYTOhvM
OYl7p9y3fMxnzhdLS7yqEnUUCu797AzCVaWbPuZVFy0yGO0Ba90a0BBtt4Ro50D0
Gr1mnbTisT4kDzsTE2NFdb6YpRDjUuBnoI1j8Hrkq03gSTl1+cv6fbaVootqJJCX
wMw47l99wA2IJEPbA1n67avhG7qJsRTxEbkDxbtbuY53KZZT2De+o83iVzHO29U/
6/odrOeWuu2UJZWT1Q/SB6ILiRitMXBD7IU/LsOXN6NkOutZq+Z899/di6FfFWr7
tQfGpbKfZOLOwcTxpVJ263WenJxR977pfvistcd50UlSwCnojxt5Bwo+iIPgMnNf
PuPEYqNzp+Y1+i5PLawmK5Gm8nlrMbq4fhWF5LomVnkJ3xDZIvhat7uW8FU0gNIW
pVqNL1fpruZ9+REn9YL8pTJJ3/AdosEU7ozm++IsvN4LO2GwcWnLHB17UrI1+0dF
OAPs+KYHENH/ORKTlvluv/IZ+EwDzozrxDVSu3cGCsNAHW0teU4WaGwr+vR1K4XG
Z/pQVouQkE9pR/5NWOsLxYUtrfTzxkyoyahnljJ8RFYmqsLYZopzVwR9RUB+y3Eg
5Lg0ot2HkPzqjfKeyGT7PhgH2+6H3QLe8TKl2XRuJhZlYk4aW4UdyHYA5iKk5Rhr
qFg2CqcNQURrNTqWsz0A7CTsbD/GfPv/Va67m91RTPWlJVu+H+1qtv8HmKG9JzHV
7ndgWJhaVNcyGMVTJhFA/TcWteVb0m0z0/ZNr3Z8cev03r2EAwuRFgURnQHZpKhD
osxuT3dSEamAt6VPv5dkaxosJ47nClJGqJAPz/r0TFxL4EzLLQOnkDNW0CxLZ5hX
rgkkjhoqz1Onvx8nNbMbnho+qgTClYhGEALhervtkhLootocjDu5xtGayGveSIUv
/BxFoDmiaHhOh2SIkwN+HHzBRVluY+/XWqzY1v4UixXUt53v6nwJ8HoVChMN5EPD
XeDh3+tbn0cpNYYBeB3TWbex4S5RbnbkRFP6NzA+O+EhbSeWW1tcIuqfLiWf9zMS
Ki/Sm7Hc1YC4OlII62FEu0uPDTKbgJnEjdFT5SRVflrlmQm+ey/PFDcIVb4nwX1U
W28vCtac1uJU+/m3pcVLaTB3giuIE6JMvvXKu3tVA3BIBSuRwhTwzZgG0PAt/LbG
o0n+tASLM37F3sK893pDsXSB0g6881o78X/fvvbRU/WDXgvRq2QKKQpcovtEVOsJ
E4TrmMQk9SoLfpsbIu0ODitcC/U6QHLiy0JzQfFs8y7lQIH6Xb8qg/xNsI1dO9KN
LV4CeM+7T66Vqw7l+UV4vWIjvmi/3iWqyKKzKeKkWUZUaJQFJ5t9teRHDAm9MDMA
a3yCmdjANXaUJtzRxjXg3RsAU8zOPQ6TF2/YIJYriSInRX3Yso4M3b1tji5CauhX
PcqgmlboHKTbWOkV04eFR7Bu3fF9o0ISe513i9exdGgCdCrCuF8WzXCl5SZdzR2n
uREjPegK9qD5ImMeshOatL8L6WItgGVXXR41+Aq4iHq3W54MVF7h/CXVYIkKHSOB
tFIBScXlhm5J/8iTDQ6RhSidupJsRVpIGlzZJigAvjGjScqC0fIjy/KG9Iuh9H3k
5Pt1XoAkh+qE3QdrQHWF7HlzOOxkcIjZbq/YU4OvBKWdGfg3yLzUhgQ3nEcEtmoR
ltBM5N9XiuT7r48L9YUjjIswDkz9ypvr99uFtox7vC0SQwEfbrAI4l0nRTOLWyjQ
sIp7SHWQBe/o6tn+YFnHWjBtVblbUnDu7mxYLspEul0DgtbzBBHUgBwXBa0BrypR
2qe9JhOcJ71sQjSqYWSiiuriaKM/2Vna9AhqW03fzvqolRYurPheLab0zlLo7s2T
Q5a1xPD9LYjydKxAZId5xYYX3NfI5yy8dkp7/WZbt/Uby8tRhfLCYAIK4D9KggBk
DkPhr0Bsq4137Z+U/TLSpLsqc8Lr0RJE5AbY6ABtaqXunXTwmrgozHOKrA9JYEpH
3QZ3AsKgsJt3MTTHmWnxNKtL8LsRwYbRnbwMpxk+aCXYlJibEzUnX0G2FNuzKe5C
Pv01uPGTprsLyT0aR7nzCwrg4ACWyQ9UaAmuV9KSm+m97HzAOUFzBiDtTHt+ouMr
CmanUtjNDPgkHsnLdOrMtN6fMWZv12LhJ5upJDaPFBGrHmRUL9Y6Z1GcKFPQbLqA
WpF9+hzlZ3dg/mcZAlEzGrIGbBS0mQ1FzdlmAuzeycSnTVvWnrZB7ZGxA284OEhO
U0W1VjijJMCnYQq41eBBFev21Zjw79v15Wn8V4BgXltXoVaLfAoudIBMJuf16Bpd
jco9fq3lPTiyJTti4/bth9phbe1hGVaZeky/LbIKD4hmZxQhtU9BboJSLNMhVcbz
CdmPMqX4jD01Qll8pwa1ieqe0YJNG4s4pohTTXbeIZxHjcf+iI53Qs9mt4z/ghNq
C/Cs6evihBAXpOVU9hY2jPxdzMuIksLYxAmYSSlC2uYFcs7SjJ23OWY5yVwd1QG0
66veQPzcvn0rxF6vjV4bz7kBWMV00gXne5ulLJ6jscOpuu+i7tJd6xScLQ++nMeD
uW1E8UnxEWCb9oxAXQERm/Yrer4jfN8jzXSETNAAuOgIZFyMtRntUbwmMFKvlvwN
L+fWbXhPnnK83ai1Mf1gSmq/UROo0LU7gOxYazZXI4ufzX+TMB5WzPAKysgIJvlN
wq1kP2oaYNsydxBpZMx4U6V8VvcOazQ1pNTxVL5IY5BH4Z7KMW9zNP5WMWCHDhEY
3yroBonwFlyQovcnJdlrm9YbXUuEvDcwYpYXOFj2I07LS4vyGPOrar9tHAPRIBhF
lRqnT2io7a3i8Mq70rHANZ/ClIN4Lo1PT3J0nA9mFbdxSU7Vav1s+BC03CnYThiF
+RKBut/hTu/y8C+g7DdlXMUO53Ca9uNPX+jJJOtXaClqxR3zkkw3wohfTnmb6vqH
CyKiVaRSl7tl66kyywqfKhBo2mNQvdXFoQ5A9wdnMSPunddUrDBHIUiiNMmLltyp
nbpsVgHDXcvfEhzCiguyiVTWMyHqIKLbqMnZ2py10bGByb+4OLsKnaL/TXdM4T6P
TdvGcM6hLQ3w46xl65CvRoX/jIuIs8RtlfYq4KDb+53Muzxte6FKE7pGeQ7lNYp6
mC84qR8RZO14yvmZpz+GdgB8wGwCRn7bzPWS1bwK361j5DXSOX7/KmqoiJHVyx0+
t9gk4EEYmG90BJSU0prMl1Smz6yoWVV1pw5QX7FKWER5qwpW/3+J4DQcDD053psU
vEkdThwigMdgCjbtvr8zyjUK/Vz+/CjoxaLLQI7kZsBE1dDrygaxenDAvR5e0Sk6
GK+hcmE3RjBBQKAauAtFnGjOdUGPeXaZ8e1lGJL0Kl0uql6eFUhVpm6VEWjG93Cm
wzXL5k1/9+t+QGk9xAiJ2qSuSoA34x8pbNtbvgXx4WzsqoD0WYbHQVipTvXaY6tR
HZIfbz8NDsIBvnBAQ1CuatdE4jBJ/MzDLa6U8Yy/kkM6JNHrSxMRvR1PKBLWMR3v
9pxlExPNma3lDRZ0IWm557voLhPqCt3JGg10ZHgv7Ar+WJs4bpEawgRLZr65+fLP
tNdjYah+R2OaL2IqPUpI1F7ts4tTNdPTwdbzQefcmfVAQGcKaY0EWQl0qNk6oBW9
1oIl6EI8Fq4pqHI2OZNJjiTsoSlT73DfT/OcQaeDfwMFmW5PTEkgt8HEAUcNhXhK
oUy9L7mrnXl/OMaKkZe36lUvWvjo8fdKDCUAaFw/KTYh0BLe42gwjZxOLkKKjbr7
KEfXq06fOvn4qopnPov7dspgcs7Ljo6kKjoRNH5ttTJh+UZFAQ3tGlYdnXaDvFBk
CapWRGzfxElBGk/mF+zG4SsLk6dnc6TVDgWymx0Pqh8uqDVmurNKH8JwsrHy3aKJ
oM07H5pTndmwCfVQSZEikFAbP7LN69Yo40wPLgHbvprye3/ULcjbAO2cbUoKMkw6
anBNavILkY9SLKIIesuwLYjVCRLtbXPMlxbvRupiL2jz1TszMNp/2mbDVKq4E1LH
2isBm/Vm8YjzFbDO8M0bIA7FwRtmN5+eKeJvGlDkvtev2GmJz6pIplAxCGMbGNX6
so8Q8LlTJ0NuHtd0g4tNDKahTpxAKKVtaanudQXAD8Y0fKtNqXRqf96ortsIE+V2
VywbfvobqBKYQpTU3Pg0Ftd/Il/Vswceiu8aP8hBSZyAxX9QonalUnX1OHaEmXl9
kae/z1SekBmN7s4QjeWBf8rrfExHeD18NOmcJjB9rPbxt6u/19Ap5Srn+iYba8lV
n3vvIB+41BGrgpxAU0UX/4/Sx5uTakOuy61b2bb8q9+SFOdqS+T9P9IEYtbnyzKC
dNhlUb7ARYnTHoG84uEUUyETQexnivDiP9oBZibs1OgVQnBfuWkbZ5drC3whTL7o
gXOy4VTQqxkpJ14TTvp15+8dzfaAGR4M+azcjDa2UhR2PCGkNw7aw91qBB/BPvII
TKgbPZ4HDTFFXen+XgZ/hCQh785ICrPBTH1JYOZ8Mn5C7ci4p/XerzYVG85txr3b
yyAlHkIrM7jO4kmwHQQy+DZnpckYgUWwAkjIjW2OHTmSsyghVFCW1B5s16LsPkgx
xm6g+BcCsWnvrT2iwH5ycQFjSI+mbZLifAl5EIfZ9aWzqYrhx9SQlDI0rK7m9Lpt
pMj0OctKAXx5nyVYXkd/byPkUzwbSnhk/kBa8hVfM0kOcVLy2d1LmCi6XmgT4QEW
p6PCZPcU4UyDX8D+wWWK98D/G2dblTqYgUExXsBTAgGiDliAaambdUQBgPPShK52
E4Ce4jKKxnxCIBcozKlTabq97HrS0LlqUzrBzhw1wQVVtMANpd80amlA382QBign
J8krbn7jvga8K/bmilcVUJorc+7QGkdUwM2L2eRs9suS49/Atoey/+g1Kd6L3fAf
XlXWtY44XH3pVEqFu3oZXkBTB/nZ6twy/KsCHgD65wAqfAS8Uo9W7WEzQEfPuq56
csy1aG0a7qrPh0cr3vhVW99UIsstOusJ9vjMB9X/+aYGKsWfHRDMqLOGUiKOh6Oc
qKgaeLWb2Wjwexo+6ECQvZbIIUoiJWkEEV5wozYqzulEMRrlrGqrxmpNxjPcNpgo
6FR89/J7b1s9CqeV3j6OkoPtpl3Vk539V43wwFRKdR/lm9lYXZjzuGW7+aJ4s1bI
EbiTPGI9v8yuvVV+wVSgbKD8VhkeW4O8e1YEv+4h41ShXPycT8acGCc6JjzHBU2p
QKu9Cu/fCJndMa9iG9PUTzs+f98mKagnjwz7hUEnEmYgUasAYFgTwIDqEUZz8/ZN
qFVWicuvyxaXBhgsTo6tpWXmCFVsKXoJV2Nm+WWmS7j0LQIaQPinWW/64uPXxkFn
7PbTdvNuLbzWla9KjUt62UqCsP/vAHsrnSaXTfXzmpmA1lLvaw1UvQfN3kS2Rl1J
wvMq2u9XyJZN5ncE9BzLIx0LhO/NLV7qLJNUxqulmdUIhVmAyX1+XVjVjh3cGsOL
gWTefuRIXDw0ttvx9dnN+wQyJmZ0WQ2kfbU2QRJARbxdp83o1jg9Py5Z6dsKL/E+
TfHy784NvRbcUpW3CjYMiVka1FpYjD2Swwg18Mp2drl+Q9fhaHg4I4yzrJn5Kam0
oO/XF9psSvx6NKb/zgy03l7w9zXNmhw3NC97rromgNGeg5ibb8VOqxDmqv9ffTR2
VW3T35e5mPhNN9Cf2O2WLJlFZisxrqvzPuqD0jr/9Gag5iKa6bwaTCCvbpTIctC7
6byPV9WfGzZfLbu85CzBp0QDblpi6v18sTQcfgyBsmGmgFUug1lT9UME3MX/Mkol
VJFCoYeCoudiXrrvsnnDI6W2rc+0RxSopfUDQAcNdg+yjka/PX8ccBMQSUkyst6c
9MtFgquihvNGo8HqHizjrrEN+VXIAnkJzZyWZQNitwOYMsyIs57ZxEmGMSd0A8Z/
qCwdzcwSaY11mhRy6BeOGXxd0x8uYybJM/FW3NpH+3h4Ad+2E9fbpjAfCjAODJ6l
N/5cn3XgBdEi4+YYLRRJiZcLauzvOzF39J32OtbMFZl2EKTpBaElI1LX36+9s9H2
sa3sJdD3mQSzlFwIAieiKdcq5jQ/RuiULjY+6Z4bEI1i7kSoc9GzOKNwHv15xKVF
Yfur3l6F7MrdX+Oohk+5cHyEGBo2ePRKVczXaAUUqyWLKuf9dwSKmdU9W3t+2qMK
ZC4oCnqUDY/lRzO4UJEHCR4CAdhRCLQRuGi2ccYqj8izKkKQsj4A1aiAYvbyvx3R
WkO2nhwxYIijaSiXTv3+CzqrcGgEqcwj081RwLEOuUXVKLnV9Kaj5KVBNB2ibmt7
TFMM2zEg+r9+KYaiTyqgPda74RLRR6LuE4nqmIbsE5OdhusVCHAUEaWqT+PuLKS8
JUvpI6sRyi2Se7wGDorSHy2KLpwrB2kDmcc5b+FlncXVkUVbVv8JX96WVzsW5n5s
t7RRqQnwNtxO9lAucvvCCCOA2clc2ANWrSzK2QepfilFwpfLH1OWZNYl2oYOQDMM
wCQNCNuBfNmPWE1e/qYZuOXK+6GH+peEPJUID4rUNx0x6muIjzxRMMAkqXz3Wepk
EyLBKEr3SZkJ6CeWbFylMESUaTEKojmaJXsUpf3ntpyKTlCpeJ/WH3ve8DfP9UlP
pX26dk3SdVQ/dBdUeHguCfInUdgl0otLO9GHMZXJq/KuxgsfN6aQs5/QlCkN92XR
DQuOKfmrK4rBifsZZXc09kyX+7gNbu1VNEXd4z4e/XOa1V0FPfuV3xmFwc0wIhHa
s9j/TChgdcFyAUVHGD+pWszyPJvI/dCswvCEFYZnd2XIHgeAUwXbKlVrow/VF1M1
cyp2QJ3zffdwbd943lIyVy540YjzrMHYHaH+/iy6eTlWAZtTheUTHIhnE2WQQP2Y
tJCYqGhxlwChAipnE8U3BuJr6CcVInNol2EClK80W93+NTf1lGI8whnnJaqisTDh
8bWUJZgpQrWgSCWwVXggY+H4y8wrdtVXQ2gHEk4CTaSD3rcqJ20z8YDNHfxEoLT8
cbZyx3k6MaqIQ6YOWXfl7ZkYQF1iJDPqRO1RVdD8dP9ukmBRShuDBdBbeq/lySiO
CScyH+mYAsY4ViVaqiRB3r/40NArlg4elRFyQJNBpLw59P7u2gpUkti1Ft+fKsda
wPGHCyuvu77BjXqvLbunRFViNbHaffqt8BZ3tNxmq2s/Qfjm3GY1Qi+XB2Rh3yBP
R78T+VvobGnBc2TO/6E8APvGovR2kZyfP2IdlCYG4fqPYUbicLKlG5+o6qqm3Z5H
qzLwUHnP8XmpSQiQ4RJUc57+op8bqh/6Onl3nD3K6FlUMSPDQyZ9yz1sIjTPIQrz
ZkjyqF+Y7hjwjdwk4EK9D5KSAEt3NhWM7+3viY5xr3U+VHZjhKlUS/UDVZCVTRGq
HTUaefdEXLmJWuFXoHASkmuqxgBlF3O/qlKsRs7AUQ+KgvFRITaL715qUCw2ZghB
Jje/KmI0ftGdopbIgqP3Ph4W5hROhmKRo488QjavC1m5KlamhGLb/YPrZX8+Cqa7
NGw8+W8NN+UFMnXYR0raS/zUx1wDoNdyyXh4FqilR8WzvtX5cqY/H05UWmLO+EwI
ARYFftaVj+ikHTjkbDjcAQEIq2PBXhPaN/cQ34Qaa49GfckJ2G2mfW9XrEqeXmMi
hvATVNwjPyYRULlR31v5ebUwS/8WbUmJ2BkXv7VRXqqF5bUPv3GZr9Lf9X2pJgyZ
H+zH3zdxO3WAMIJ9yhKlI0OsUOITycT78jMsb2k+QhSs18tcVSlW+TuBU0kqFeJi
AC6IeFdaGvHgTCd//IQdIWb03eOqAK7z63dDutKdXr3WGRNrB6c4NfBv35nHVqbb
M0slmkmC92hSvKzy1nNGQz+IDG6M2/szHIg3eVNc0dqZHCW1wn6MRO1niALK0v0q
Z4591i7F05btljNvukdjzaQkId0/fEgVu3gmFQbCoUO+cymJ07bnq5jdsidBr2ZW
R+ms2fSZf2sfjy27lC2U6P+HT+wU+xQIS8L8qF/3NqHsIfXzGCFrt8HXAdc2QIBq
A1LWZ7b8WYII2zY0RPoLgNWf13Y0FhtjWP2AvgTB87saE6NTaErVvvI+S0n8DjdC
NsC2x4VrEeV0xEJRUBWWJAVaabCMyj6gjz1OdMb7Ecy8fFJKnJXagaY4P2hzFmCA
L7CqCt9t5wnXCVULc0v08XFZZJ1Cqx6xzWLQImnhxamMFR03diCgajc4yVuBFR9v
sS21jCt/BVm+mN9BUcq0rt+RmpA7klN5ExAQ3bPgRhouMnTJTlvxT+Yficz3i8Bg
wTGQBUgpnPY42PzTVsveNuooUCaW3gJMpRd/T5DJYRPiQ0h6oX51YLM34xs3mVcY
oU17TvSmS5zTB2PFt/V80PEtcFPJJpM0GPAyZKf3daK2RnPCd0RSH5reY7H2y6Ht
FVfs7F5gMuWLOjkfGtsYbOSb4ryK7qElHqX1AvZg1BkM25qc7qPx8kBiutY8/tZy
bdeCVx0qZiDaMT8Ht9DLYOKPSkIvzVOw8OShMSjT+if57DAeqmpeYlW952rYUFnP
41TihSnfri9ydoHYO8SwomGjc6rm9u7dbIy1o5W7jirV/yur3ZRlHpBSgetkxX3O
H+u2mXLrvc6kYQxaI4oZW5wlWp//wLrXQmVCuUSrYyMdEk8mXb6Fr0E3lfWO39VP
kY3Sb+QztluMv1MCec/z4vVBhakQebzg4iiPM57E4W2oNy+uOIGJ81jernOwVbbL
4uzW4Y4sxA+o6jAq+452oi2nN+is3Og0aLd4GhHExaE0Nd088RKupYZQXftHD9ED
AjGshGo12zW6g+mk3J7EdVGIZnw9b+ujYnZ8I4mOmn1eICDEa6e7cCeHogmlBSQ5
PBP7ikyBIshWd9PhLgK4RDe7muix5OwBNeZcemf5R2F5rWPByAnOi3qDxVfEZxaO
kV+DLzS0Vgsu00zM7/7k2fVFFORSqZGCeVaFB290m7S5p0hT66Ajgi0TpFDm50wM
j1yacblq5QyNKXPHYplyKRQMGPz2zkMkPubsCs6YL2DrQvMAsNnFSuIy2Ur6tjid
oCdeywUMzrP66kt8lt8n/2mvrwGKJOo00rJoAHUw1r0aANHsfuLxzO8A+Z73DWjT
230hWg9zFG3C9zx6SsXn4r+z9+96Yp9XvZNPCvPjC0H1ACHGLXvqcwI9z40D6eY3
9N2rl/+JYVk9yq7Jh6XmLKKgA2gTyrGt1v3mlOieSOicqO498kUIbA4LDJsFfCAS
UtC+vwUAELpgJ73/SRmPPVgsd2yOVvrVxOpYMv/hESjHsVobUGiPRMoHc36npSys
5NjjiJ0rSSZQyNZNkcyV8HtIg1HEOGq/1TqoO/eTxu3MGm/meLjj7AGQkNCGkquU
usfjnzjsAnrIEEqs1XrQPxrKyJZF4yOwQ2GPD91ezO3R19ph3us2dKKYQ7OrJo0h
MASVGUUfcF6kPWe/ZU0+vvMoEgpbLWHbMW2NJquo6aCTy02w1GEnMgp+ycaRbKGS
IUUb8zzqKpg2RjAFhzOo/TVnpMl1q+dYjy9kdJgS14VOMAMa7gPp50DyD8grou8O
aWI314zxD7tH/ZBW1h/U8EaP/2ng2n82xQy+BtogYjY72EwOLf/gy3CfHmvWzVUc
OsVEuyLizUxEQLTWipvSMnUZ+iv0hs/ofuVj/dZT6SiejRAU98nFCmEiGcv/OyKF
LuFlQrOHhWtgzYM7hjhrm4kN/t3E3E0VEQasm9roCbX9mGv/S6VhExIbbshd5NoA
BRKeLR5Uva/mHMgPbIFxZ+lvuPaiX+y7kJdDoIypbHA2nPB3ORSgl7+56N3xSUBS
D/qtOrxMKv/pwb64BYTT/7Rly+Kp0gC20hkYMmPH9P/Zoapc9OkH7xRrSmrYlig5
Kg+GxZ6EwQ63iRPx33Anmm6EtjnA5QRLACKuNZr+/Hrwl0TMWzmWbNavoebb7WF5
6V9ClRBMt6u/yzUC4Oyy61GbuGLu+Cg8SqGxkN+p5eriCX69ClOGRIWLo8dVVE2G
kWRc71u10BT2QT7NTScbyGnG7pupZ3b/gksPFhm2qPCVU+kAMVmENK4R9ktbmPRv
/TEvs8H0dHxoBmsAO4ymkHmybwNaciUx2b7SCJIFdI07UqXnW1gR+hiGELy7jYSK
7fKgZCuno16zMY8hPn1KXNU4Hdes/oQjdqnonDmupvBBtqo0IT+qEIUfdhUO67fE
t6lwF5IH94LpCuRta2/rPDtWJlzmoHhgd6ao/7fkcGKiosFVZMrzNMBi/ZZ3I00V
dyoGnk9sKCfVFpJ8g2FnQT5Dk9naG2JF8vKCpCsfYEhXYJJwPjrdZ80NksmkfIJw
2yw3sb7lihAEi6CEQEE6ukV+fRmJ+cYGOQGS3peoiKCa0VUCQl29XMu3p3+/v2rZ
3dl8rXbO429AoBikmkUThyPer1a1l62NTnlSdTmhUdDCX8hV8rG8dQ8mBU5Z51qx
BPhtNyWRgvt+463Rd8+Zke4ZVwhdo1tduV2MPVhTTbblTIKHFOTrefQKgl0W76p4
d4RrE3TPsIluAlwkv8nfxk9FwXrY8jxWKHJc4IF4O1nEZC9j7Ds4NUd2UZ59H3+S
dCcssvWHQm5l06QX7l7UxQ/2sbZd0wwbegf4hBWLGDHMLqvEk+m8vNNkKxN/GAJL
Lb0pQtZJPH5Lite1ivFPEs/zfDfFAZ8c26S30+ixjWK/Fk0udhlDTHHCk6G8On2K
XgY8UD63KYwIOtEucCxbwMQTCJfqvhMq+FebaVz56v5xjmDJks2nHEC/A8I6LKhz
I45l2cUMcCdNdffwMP7wDopmDuUAFPWYVJHMeseCoIZsKQ/9JcFJQsKQrgYJa3Tf
M8ayMV8ItyiqDiuOFuGSTuToJRE+2eQMnTEb4HdfR7egwj75VeziylE7YKQoB7xt
kB1/I8uTdpm63fAfOGv41IJbdJ6XrM9kY4nJDLhacU+2yFgwt6RepEFqO+hMJr8P
zLhVDGUNu2zrL6QsV1H7A2Psw1V5SHeVT8Dyzwlv0kiI9T+bynOr2xEkGC1h0QA7
Dr0gTtN2X1uL8sqHCBS2yvDM5Tt8II41kVRwh3GdqWrak2snPMeu5FZQU5gUtIqM
TDqxPtEZOK06chkDzm1jEYilA5epoC7k2ko26VPEp958PvXloRMXeawTrBvuUxO/
nk9LhRbc9yWi3pdvXsweWTsc28W3nSs4uSpT473woWcfN9uhZGijCCMuTWVn702o
iU763Qnm7VrZCEYI9D66vhGjpwPy9VDvH0tDKSwk1QtMvzAl6U8HaeTuSHEOddoe
W0hcSHGqw4qVHqqoR2EdJ+fkRAjfZZvvxcdPfvHgJLJrF4uWp8m84q1fJXL8E+JH
UaKx4fNkTcyJQ1BkGznYPyw/zvxi2NONEkaJqKFeC7RGWL2Re0VrknJU3c5EXuH4
gtwYSs/GlUeTL8xeGytP3tm2EHp1HmdJCWkAH+1jDqAQsrh2ePYpSnB8Hl3xGQ8q
5SnvCtnQhCxqQRo7wPsmFuMAhjDDU7v2Ml/ehTv0V2btyZ/N5tnTblvfSaWvoxq7
Hb2h6po9HDxa6JfiHHz+w0clroQz0lDJjQzJhP6snuex+6IdbDqI1t4ZOA63Z/B1
BBMlMQoLE/C48r6yAJhnb/TkaBVs+xdDSL1CkIRBJQu6YWihxtTbDNIi8TNhnogS
vrC7ucja+Zj2dtWp4e1a0iZHV2DxUInWs14DnOmwdhfIh9LEsYY/4gHJ28MZ8DIp
UmYWihSy3P28W2hq3LYAdJRq/eWvPv1kosvHj274n5EdxEkTHKYnLdiL0VPomHPl
ATQwFH8ex2wF+YiZ96mucwUpwWTJimSULP/Xnjjxwz/O53fq9A8+717YMXhaFuBV
jnCa2KtBBr2vujLBg1vH0cBPUG2ZaMk17ITtoW3CdvQzqrjg6DQPm5vOJjSQW9Nm
9hZVz720dIXvlZ0WM2ZUyfZP7UkAT8eE0KC0DWh5pvIeQAS0yIicEyMyACe/Sfl8
vXXWllkAOpIJJfvhY2alzP2nY6gqJMh35edXnpY/y6TtwBXSgEoQRw1cOu2NgK4U
97o0kyfrKrUSa6okfIhZyrNzzz1oUNTC7SfkouffgdoP/01ivoFvadgal9NHXCH+
1ZjEjFbnykEAZiXyAVZPMI29XOvIuRShi/jQ905sg2wAkWXn5eHNpGy0J6JmfSJF
UM09Nk8og5+e2DWq20rrGa07XdAlurezHV7wy6DQjQJE1m3ozXpEHEEI9Ek4eAH1
nV8VXCoKC/CpaPCUznk1WQbu268QYQo3lCQVzEMHLewA8FcwEEtUwWVoM2s+TyHt
9wZAbgzil+yh82NJDKJkWSYE+4T0wB3yTeEcfo08CmVJfRLI74YqUFq3uAPv2TNR
c0vEJwDRFP6zoXVl33RxiyQ1Y81JxomNpObXDoxAumiEmwCnARUfP+c4gSnw+WUd
gzxsahNE+bg9N5zo5UFdsBNpyS+F1lCKRbddouJ1KM77i/EXLh4ll80fR8ZxpGP6
73Ux5Mtmu1RioK7j0yBPF1q6Ual5DKzLM84sHHqGi7B4lCoGj+nbxt2HsF3Exd5X
edyu/wZVFMTD25xNb+pDuGEk2Doe/n2ahJnLwQ4aNmjd0UYIwqEnPJjqU91dox0N
i8Ww2RMi8rI6J6NLY3CnSNm4PIEMao+02nJ5sADeEZoM7wKW1OPdu2y2Nb9WCkvV
q0KacchCp5kRTmkmIy9PfeyDpS2Gc2WGyFCyfx0/WPg1+WhrTxTXQ5fQzR/vq61X
Vaaumae+EJfnL84FNKjzSyikW9AhxibwggLoNtlePrjme3EiRg3eW4k/SCklX0mT
EC9klolnO90NuF4eSdbQYOudS+H51d/bO1df3P6zY4i6hJZNmoy0mEjfRvi0lb9P
ZJtTAZTZ4JUKRqYZ9czkk3aSGaVawbtCYVQHv0P43e85j3/09X7Kfkd1jpR+9KLY
2OjFwW5S6Ia6ZRjJdsXNcoH6EquJaP51wa5ZQWAbOZ6tp/do2O921jj1zDaQONt8
DBri6IvqVI4b9cwWzCcdulsgXEuRJwxfGnTANZhDQg2o1l/bLS65kXOaMKjh00zo
2WGjAQYzn2XtZvNB0OjJXNFjbI+F55SD7+ADhJ33NOz3+qoYZifKJrb1iPBuLuHN
nYZwLWwmyWs2E+ZNZkaaNBYpfw0nzrZcaOffO2vtj9l59swr5vVSzFEACqhSTxhC
gl3hP5Bz0cGsm0UKRsGI3KFS/Kwbmue1qDXxN8PyZBxv8p4/fMqV/vEbxdHuOdcC
y7N9jGO5dqSsjf3kcbM5hUApKYwNxFh3GX4VbGMYpp1w/vEA/nojARz7qVZQ40dX
zP9O0KlshbzK1k7H6q1PWQR6FHiPSo5UHUVvqLxWdzBQtpwUvAHiCTqF8pEmT3ZY
D+itHLuTjOXFdxIa/MW1vrSw0WFxUTN4MfWhB3BYhryV6jWdwGoSv6BQ/761F2e+
pMJ45jYxSFZ7XszI6Pao5pctkx4PFw4cu2WrWoMO60ATdFHIS19yl6CC/XK6JZYO
LKzyBjlfUoPZDlSq6wFmGl3zLGhkrqQkmJnoHBzKlTKw4TOaL9/WJRWJ38lMjCjB
uZSipIQxgZ/6WStr2Vy37/eTNEc7F9BH0/OQNsUPWTj89uX3l2Px+M/fTksbVeWX
SKH4aXCDQc7SV9XqC41q8qKmg3bC1Mk1s0tMJ7vH/SEFhN1taMg2bdngd4KYWmNL
nY1STbLSp4F8SvkIurBKZf+L8ExeYxlMv1VFj5cN7jl06eYM2wr1Mwduc5qOTYdf
xEDJ6sp/jRMYsM8m5+iNgeVsfWf57DHbDi1NbmWKCOoLcWQTfwHhy4gTmW8J1ncS
IixDwPWKbD5P8W5LwXXpRaAEwh4fQkLodWPDfaSzm0JZa/SKAP1ck/xon8lAvw3p
nsxTKfWlC6poevs9fMsmc9qXhiL0DWlvQ/E7PMxJMk05iZhpE89pZ0n4WZbfsK+B
SeRbOGXKQSkjUZIiNbOkTEaim1jIP11L2sahmP3PIvPMBUFYxuOokSq7g8cXcqjA
mQHpSjir1r42BI2mSxe77Gd/ZDBa/JwctonjdAirHFZ++62Btr6VrcUks7LUphMX
b7gTbHSJFyEn8I99TA9uoyhRijJbDxsoF2+BBABfm7bfiInP6OB+6jALkavUq/IY
9V6ecuwRuCRX6SEznEDqle7G1w9e2Iz0s1pvPyefngOFHnFyLit9hXMSvn4ixEa6
jjX7NRwzABU47ClnOG68cyqz7F84syOv/WlHOUD7aOEmexW9uE3slXWKhElgTEBN
tP49ckoJP2wocQUxGQlNcGb6CbViFmNLlft+RPNHnkXf0OtE8gibqAj7YMKK8Tfz
JGisOi6I3/iFQx4yFrnwGOPFUwV1tIm9tdW2XsFI/7uvc/zT/LQduay2hVMfqvJr
S813psgVLZRj2+AKlL1R6+AwaYdzmJMBbSfEmbkfLqn1TzTvjoKdPC511b0NmT1N
geW90o68Fb31zd14JM5cuBeZa/9izUNxVEobBE4INYZiEHCqnkAndR630FFwRQQa
df0k1vR6mBxZ4DvwYr/8MNDnDjvfS5W5iObgSdA/9d6Gl3dXpt80YcEV5aYxSlqX
xUiAl+Rpv+tGbJq1tYyoHY5HzHAKd7QQVboGw5s+33VfwWHz0u/47YbtYp+odgj7
sBkEPp/e8LjUexLfwMnsifQ1xND17NqSvPFlkEAEJBRozG6xIWz+rLv3+L/eodts
2P8k62VODu1Gf+jszyTuA++nIUNpwZ5PMfPEO7Hss+No1RHqLqQnUf1IqVq67HC7
kX7RHiPmpu1Xu2kGDuMIu+pgqshZ9n1aODsA1TJWv6I31/aD/xX300BnTn/p3g0Y
51wjhEdG960i48Q/+ytJQUx6CwPFvQc4DsAV7udRPtWw3P4K21iJj+PISNz+FiBJ
xm/X/1IVGIU3xCMNiOpOqiAzCqH6ov39C0xu53Kv6Jr4lRSFrJ1VLmNV51mc7JJw
N8HA+rDD1exXYGvPhlrxTEqzPpYdKje0B6HY7trS77IcvQ+8uqQ6X2nNxRJSSDvA
N5CALnfss9bsZc5CGBfNTvs2GsPYyUAQklFPpExCfGzluC2T9RvN5LbtlKXUOD33
puVZ4skestWM9B0j1VneIxpoUQh7+l/DsvQcNUwCC9PTNX9Aq4QeMml8wlMQdVxO
mT2nQ52rn6+vUXxYLuGeiHFF52YU6kNVnANFcKmF3rTs+dZMzMWhl/azMcvDVx8Y
4BEDA4CaxsEmbC985DKCrTZIdhtNjy8qOJb5Mh4EvNPqlfK720SczA74siLld+eb
nW0P47n/xja1bbZTO+bIsGV+8fzFECgzTgaYDndh5hosIlRKNVn8svGS1rB6TBmS
rwzf+yzJ9tZi7uqLgMQ9iFd43YRiW1ejVNX4PNZtyKcxJEeILR7if6htvBBmPrTy
Dyk9WDj/J+z0yiIdgCOfZ3s9CyeH7n7cTatYplLcbsh7LZilHhCZctPfRDT84pba
7LNBUOGSZ1tiL41zayMD4D8GN3P9P4eV8QLjwWCphanNn0P/EI2ziiGCMRNzGNwR
ZPQwJ0/aZ9vgiEMzFr+9j2tqTQU/G1kUegZKCwSMH+JULl+KsOrkjXK4dyafNVKd
kOPqlOcexg4VA0uivitMCxuL7XP00CiKIw7dYSN9zQdgo44/eRxV215vIAxYAv0k
hSwr3G6RBdzvmL1MsS86sek98m0EwNAtz5CJvaxm/VqT8apLWoTPqdepnRnozphO
rPq0ROnr/O2D6VWEVNK1YUD4D2f55NGdt5azvPsyIiibkacLY1SuBIXILNqcUTHD
kmdYPaafCinAku4/YDP8PRkqffX3nwCUgQbtQiSz7Sgo3xppJsCJfDoyyD10KmVc
n/M+idzoAEXpsYq4HgD+rX5jSbJfynOn/xtr0/iDxOx/nI8zvdWbYNoyG5jBTA8j
XVSl0aXbqUs0YO/e4R+Oq+Wc1H77x9wqDxtVjzKsZhWrSlcCEOfahY+NddjipegP
XQkheGWvylT8jcOObQUJ5Hq8OmsOqmsV8S21AZc8+Iqz8uJ2Ye6Y5z1Okph6Qp5l
NbJVzsMiqJgVRE2PK4XU666rGICsneMBjXGzNY9MzhmroMcVuOXI61PhF7qZoFEZ
Sx1Pl+4GCwdOltnYM6UNEZb0CC6sITiEsyzia0JKpioTXgK8vjjnf3YyAKrUtpIT
+qNyfI5Bxscom1LEvgbSvmZv0qqxsPN0mIxzrgf3eZTGQmqj64B9uVNW+jCxOqPH
i3YohjZGXmPV+253LBxjSN5ETaD/RbCeK/YCd9pzItdtcHoqRQP8pS3+X0ZHpwhE
iFvdVoIkeFmWYCXgtjWX6TCr4Mmye3cq4fqHuE1onfDSyofA5D8wu8loXndoMuz3
srFUAfUClvgo+iU1U0svmWWL+qWiLmo7Xuhg/QGnVy0f1wDpjA4SLbJyJEtu3EkR
EP2XOzmABP045Ukpq1S/GQyJiNDQivu27QbR0ZYqojvHz/GckJZUiX0YNJsb3De2
Zl+6JK7cUEBit54R3k5hsP4XkVLStuUuvo4fxurbB+Wz4BLUDiOoN3TDkSvjqTbP
YXjxl+8iI7GTlHaHEHEptsOnpkGo5vdHQxlMoz3swYPtPjGrDplZ0OQjNn+XohvX
Fis9EkGIhz2n3//8jZFlT7vNqyb10gTFU7N/9g1Ylyvk+7knjdYq5sPidyDVVe87
S+baprKGKJz7PJuz6imrF0qiV3NNYlKsdmnPL3nycT1oeVTyCBlvk1uvgDeZQnEN
NsGxLHp3pIgd/L9t5OXoZq6m6bSQdXwqLvCUVUqfYnZW9LBJYNjET9Z+sG+bAs3i
Ji0am46j5Hsdb/GbjcyngCmGQ9XCxfa3aXHvRofz6RLoPhTfaVdzATk/5rR1ozo+
8yLw6IbIKMvFb6mdXINDcJUGrqy/mlVDqA5euDFGy7+yKiowin+nTb0gIwsPE3wo
GAhmL/QG+6S5iYSRL6NbpsUKWj0oxaDne9DBWctSSFEFhzQqZcTZ3WnVZ51ahi2O
mP61l/HifAHnOVRX9pS3a51dBj6Q2lRy9/IRZdhKYsNzKnk+OFgsleGyzVBUTBJs
Cpt7axLnn7YD4oGfKwNAnukkN5w7DwM6GOMOFDkcSXC2zzIWDKj02fPMakKq6/AY
X/ped8+RJ0gDcPSXzqfrE6o+IdtTOUN2PFH8y2yZ2g2/K1g/n0xPjSYtrq2viGXU
5y5yGo7EDnaOjRkxE9wMdPvplsrmy89kcXNwENuuAabSpR+JQbrGdo5CIx63RZpf
EyzUdp1aJZQGSgo2Os18qEba2BWxWaLthwaHe+bPZrpSor3v19CrYQOOOOGmDRzO
AotG7TzdU1a1z1KZtHyVnz5TnVuuGho2kLgq9l8juSSPE5YN3lVFj+vDC51y56ca
UU70Szi6vCvWv+v6DM3sV0P7tzXCyFSkchLJD5kkDytgYCk9hlfAShujHE/6u1TK
F6rMZSmbVL01RiyTEMG5lpRCwY+MtPJdJysgCjaE5zdz10auxh/ObadFCMPojyiO
Ao270YFLgeeNKX4RcVTibN89uS6ufl/p9lCeD1hM0yoG5oQa0irpeNlfvxUZPXWl
tMgp0M2seMTBVBN2lmvYZawux0WQXqVtJ/PwF/ebcZdKZ98Y4QIcca+20YpTjQOE
lRahtvZIMacxJLz0lrmdZxbvsmIWgN6rDgDXT7X48Dgf3JmgCb80Mm+zlGQuQBMV
bXJKRQsTXn5l8exy6u8GWsuyX++MYS2A3QkALga4Nvl5svFDGcDNrte9jMJqlU5f
82sPQS1T8Q2GXOVFL38/kxqaANZnOkcpLiyJhw/Egs25V7ZumYh2vij82O3UPLVd
HjeQ3/1mVelQK0ZKMOHGsQ7UF/6q8veGLzK5X5rvmemfwhmtIEwEHKYAFtsyYPOR
cuSixBN7E3q2+O8DrxruVQ6Z5P4n6RJpbWE3g2D1zMniawNVDdrLg+OYcyh3Um1y
lyIiJfCxBzPyMpfChXW7cChMhqS8LaSXe064wBf3/TrOTqqBxWPs6NfIp62eYJCQ
KIzF9nU8Th94m+yrhwJ7OQQrZf89uTwLMzcXaNuXWirshmoWOqPQsNPHpfHjSQjv
BUcc50VSZK9UaMd5rnw2Q4CjjD3P6drgsCv0jWZc0p1RB8kgRLjS5nbkeexBAFHn
OBN83Po1d9AQkMHNkzk2wL+op29nh5cdwVFuXzlWuPBybyNtsl6rAJAk6iUzud4/
6r8Snl3IgqwfJ+nV+67B0GK1y3Rw00V/GxsAZOpUpvWEW1gxB5o9tTRB4P1umSF1
083qyhnRmVoGqNq8e4rMBCqnrJbwKnm8kZFdk5qwyiYmw64+i9st8WvtuOg7XiEb
AA1QE/rt+G9JcONNleUyq/0kr8EkUHvvAElEU0jC3ACGppuBaxl57MScQuYKTlKr
NBSGKdykt8K7BVUZKXCwDHblgxGmpJh+WP52/pzIfGOySmSbVUzjjHKZlC5UsnOc
4ySwDImlMydI/RdCwjo/oa7OmCZDbgNyUp8JC548DBixd+paTcr4ClftR3LOeGw4
VY5an0AwpTkDr/5xd7Pi63A/vFC8NcupBigQyAsRPZ9ZjbgQtMlHsccczmxN8GiS
++kEtWujCNufJ/F+iTl91tYLoQv23NuFqVQBFAsD2weCkRYS+iBhc7kTiUEtuXCy
I5qLthznR6J/yoAYmSSbTNEN1EWp4Mda9WS56mL9Sn22IuSxTQb1qygIPIbsZovX
x2uXkSLK5UmX9hRTuIbds0QUybgDIqXzBQ38LBL7bRRucXKJSuLZwlDoAHWGUDnp
Ye29/p7NJRhimNgXiG4utUd1xOQsdy9QBBta/MoDvjJpQ93rlqrpnqJgLUpdz4X/
h83pJcY3rbw5sjxrRrPaVjTVZl+4YyS6i6NQMqgnLcLXl+6AietgCAYMrhEmgqHM
kQnhCv+f3HAAu3lxCJ14KgCflnMeCZj0yGO2wLKUiN0LD4KhO+CBNcerDEVsoXUx
9lzUuYw8dYb3yPJi7RXWXNIi1vJ0jCy6Ow8BskhnwTmGDjFRNsnHBZZzpcI6l6KP
XuZ/QClSG5rUAg+wMAtamWuqnoS2uIbqno5zqoyMbhs6InD0/7EvIVoXU7so4HQF
F1sbz1epUy0MSH0KUYOmp65KsbVfbVq8JzfgJxZqIOYB4iizAx+n7xPtUlBO2eIS
KYWKfSiMEdKyzmCDTxP4BwcQqlPT8++0/FESYIOGDWOLuv3iSVltgWY0TDsX+ySK
kvzn1Ulf363ITKYYSFhVklb4R1pXPxsXUrwUgIT9jXXX6JXphsJ7ZcyP5neIO7pd
qmvUU/vKtNhF0Zr18kMRmKUWDKj4JkWwJ02w64izt3JklbXFlTsMugonLWlSeTUb
6FVcyiMQYW8zsnExD9jGduldDI6YO7W5D3uyy/aV0MHMTuAoT4KM9hy/XR7RidJl
0EpEWD5wcRDxRJocUGhaVxbNZrzc1YMyP0JGrqpRelupMZ5xH0gNzaphuy6NF3f3
iSkoQmOi4WxfIHidnSD3SycDpGHW5Wuc951q1DPa52ehU486QbJvP3u2QMlgqIPp
W7AzdH+YZtKk5OoyvXpkPsRPzOgObaV21UtenDXz//IkaJEqEp07ehsosOO5AjK7
bhrVCzwjizteP3q8VFV721gcZYBgDM615EZVjvvbLPzormoBPnBIxQjtlWMTJgt+
/6Q+buzK9UZ7yJ3lNjQhlEuWBHSqcumYy3ojkrQMzNqPEuy1BnMgkylL574OQR5d
DNv7vQpiQEIMNLNhCMQTA0aEZAjLeg0HV9ZViF/Jl1T8ce9mvq61+Sf00nOZEluq
hGfdrkZdlO8oFer1F+ggQ/BDm9VodmLChtA+6Mq0ZLwsBt1y3MMI56hzPIHAIyBq
Dx104+fMH/rM3wIU5JRI/mn6K++9kb8RCw4MDXyUCP6EChssK3uSU5pb6aMvFfCZ
zLNN3QL1m/Pi5Mc/pE29xOOOIEwWRK/lVha1g8OgeTskOXPTNPAKPewXHV78N9Gs
O+33M33U+1XGQFjwhC7yyemB7BV3rAjb63CInoKBdR3gT58H37rWMd1U17kfnsZI
JAfvp9C4QE3ylilreFkH9+EzR6ju6PmW7Q73xDQaFxU6mLjLji6mK4dHl3YRrowv
w5oKLrf3YOxRycY+cLcnuzIbg23I2dt8DC6iRsalxo308uvvIkFbZgnU1LVzqG8b
iZpKq+hdTJQKR+owJ5lSFt4lGbaT2wQxHOW+fI0QZLjnAtmFKU+/d7cvMLmEvulA
alFKPaTnQRk3UUa5rTpAfrS3dhtUs2xYJHjLp1qSzrRKQg108bfN/9Aj27Mf+ilO
xm0OWKMs71EzeAJjOyMWavWe+lyMEtfTYkg4pTMbcOJmBrorM9kd7CLI+v0MvtwM
vXJj7YC7DP8f+QjBPKoZSaLjdy10yabp+4Gya5aicG+8RHMW04VM6HhTqhObXGfv
43y5/vHrQVnW1tMO+kuY20g5RsKH50Wy75DofIHmKXiUpMe7d3Y5Fot7vMeBX5jE
1bIAmXX5qGSHnZ1dwJC8JpE26osH8/fYj6f3Oe4e60KtXn2uoX3O5JGHNofHIRbr
PB50Y2hh+C1nBW8Q0htZ1rEeoKU1t1cg0khfySat7eyZxPNoMAGlaCnlIGOp5RFH
UGknyCN9ZhdIIR/Cl/mk4obNoInhkZbHQjcR8PUxjJBmbPeY+xmapluvfXLlMiYO
qj/JeebpAuPNOaQj949uQKf+4tLLjqaKtnheger/zAntGPUaf72pfeZhtd5D58IY
ozCmqtS7OHoNkSf9Ugja+188qm/HG0HTSENdqs6VKrYI1rRqSGNHiqPrqJPu/2jT
Z9xs7Dgn3rFvYPgAwwYJNmsN18671yjv403qU7A5SMaGLq36QLLinGWhDSabR8NJ
FgbskwgIOsQj6nQnX6Zigr7672TrKHVoFSeSYSe+oYUi43IoCKSBgE30oqYIA1FY
/kf9twzeZCTTpMLwQxk2izqvYrig8/ZWvWlJXRgKmCU0F/Gwt+lDRde9o8/4VFLt
QJB9NVUYR4p2AaU42qqNwMOjcmF9U3YLqIfEomE+Mpu+3NNKUwZr3p/puCFYGCDy
hvnTEoeB1jyjTzifpmcKqSBzCWJ+qRRl5sbv0wVAhFocFkPx93K2EmJRuR6sMlb6
wOaXTYztYCd0lNqc0k1mrsucShlSzQZnePl2qRAb54A43GPuPgPOO0RgMmiaRZc0
uQJKLXrZxJn218gQOnOu6G55xKTItlqrun6kuVx8rAF5zqczlNfwQU3dLswYTCSB
RkjmbC8P6zhVj+/NAOy+Bc7gUPOVbrN9AdDpshgu/PmJapwo8cgy/idQAweZHyzL
qb1zNVLMG9K6MK2CRYuHsRuJBnDC5/fOowNPAqgsMLqguIceRQhLztETxnvml4sI
V5goHy4Q6KQTH0qK3AEFf+HfhTNG18+ae+qxy1w/lM/FiQ9iPPTGFWisXfHEQ4mf
2Dk8DKz/lBX94F89slZshIJQtaFG7Sku8cLj870ENENSkzBCXFtaebBVHthtUjtE
7WhPuKeyiu6vRB5pNAzmPnfgqH43Fv70BPKDx3vqenTpLzC6GoFPc+Ae5Q0LVtG9
Lk7fGwDN27tWFKoQre1SrJh45PaxkY++xoL1Gcg5rQ/p6/s+USXzfiEj+S0Mplal
6vR/pV7K+IpRV6ZuoaCC7L9xYF4it89SpWzRRJcpzcbrldwj/cWVW/XvPIa39zXE
lOa6ha2AunTk6Pc4OfVXzu53rrQAbGkp0mzOs22WqUkPgm3Y8qSw1VJRjVtm7Nu6
3iG/5CCJ/JVGcqBsVoETJMGe2d7Kpr24iz4l/+gAngc2qXtUSG5oU50cW9KNLPQY
NtLAr9kgKcHepuALlalOs6TmZBp7iaxDqKlu1CmEzCpk8mM64WYPO6hCjb8s5ReB
7vfI6Kv2SylZFxxId+niTNQZydCK5CuiMhiazLCtSh3Pfi7KkL7vzCYJqE3uF1MW
4dd86+kiHjXvBTMKQQUW8NRCEWJYR89m+ItU402pW4BkVHp6GluaNRv8ucpkTrj3
yM5qskTTaWcHecY3wjflm5G/L4dZFwTBXvm3aNvceaYsmwXnwzFufhkfcHsbEh2O
8qWZMjdfYemll2nhp+6CEAyaN058fOqUmTVHSAftMU4kDktZAhdxuXNBhY3al9tw
fKSBzMkj4EGZWWzsc8b+7VVLQkHNoLzgUvO55uBSzh6nV8hH5H+xCqKp5zuOngb/
Yf7XOd6/xonsuRZv7aSbcrCOkIbBrMYfMIzkcROFXzN4IO1Ac6s/l1vDLIFpO5gY
1OGp2tp5TlkyBMmFaAJMvj4YIDAdvGryMj2hNSsu2ONOh9xhM3LRpHcGWh5Dr3eU
8wuntkH4kkq9U7ARYvxs8AzJNC3p9djA1d0U+kDuqaAQxAzZY1PQERO4OBbGR8kT
0F87jeQRKzLIM/nKIvP/B+jPPK9rN44qXRmB03Yn/BrYkCw1tIkT5GUy6SGQuWj1
bhbTjbuUU1mL6pBvlNAWwQvS/oY8qZ3DGc9Y4tbMMmxAJh57Chvhk2KcqfYlqHtO
yKdCY/WQY3Y+VvBQPDl5VncBD0B+EQNPL+L+6Ee9sDeNRLFvqLjIlUEi+YKIPNyc
SJnMjOikXoaC3yyQcfaI6PwYJFb6/gUPzkD8otV+9brKfHtiWQUYAk9CwQxNa66X
U1Cyp5F1XjpofBdqxaSV5YEqWIpoMvYKYfwfS1fkrSG8DS7qxtYlChieIRUOG+vC
EgmeXJ8+6zANyznjSj2r1xKJS+CSjH7jOZPcxRFHdHeP+QwD6zBTdnmn4SOqxe/1
IiJRtIsPx6Cf+SSizJwjpKHp0dBo9p5ijBmuxJ43HQq4jlHwaa5HyOeusOm40lZk
JomiWRIhqjsKhpAksgAq5ZHoAJMKaOIfTjnV0OaUEv6ov8rcqJL5TsFHFZceGN4i
beI32+tP2Fi6SsWKT0l64ZtkzhsV8A/NEuVmVPpyt1Uu4gBAHq4YJfr8buzx7KLm
HNK2mC2tVD1FtE1SOpl+T7fhoy1ZgHXmMbaD0iCngh7rpas85ZgS/EG4DtsRXxop
BZk0PYLpoRIpctGpVtsLs8hAW0LrLIbsiGXAIdnrk/9GqWYUjJ1c3AWHxDGbUqhQ
qbCcyUOLKwQ7uo45giudRfltR3ZtHT+q9v4gNKPs+mvNGhkmD37Hcmu0gUr6W0qV
HhBKDpRvF89USnMXaApPhP6mPP+gSAaPMI5zg7xQFl3pclnbx2j0N/cG6dUnQWsl
5uNkyipCErhilXEbjxMyb/QYaApG294V9Jbp740xA309Ca0Weowi95ZZFQ3gpwz0
8FEYpcLBhgnYIeVFTZRYcCxnG8cvW1zOyplWRq7nLVuslJRh1p0hE2Nsv833ghus
evdPZXQptDVAjT7/vqNt0Kw5Rd7LPqmlc5q3LqROhIMe0+WKPBrBOxKA4woyIMym
Q/0TyiCc4P9WQmRDJUdWvNkUEPZ5j2EelCqDKqo8Yr5wylzk/hOGeejPF4CzP319
butVV5FFaSd+QapT3DMG9ukMR09jVnOSUERuy2s+JNyIGfRgR+7uZ9u8x/nFHFb/
k2akg33DnlwlnBs6ZFTC6uXP9+mmOx3HfZ5KYkmGxZv0u3KEWwoQEBj3m1vDSvQm
J/7uxepnvU9id2W8kSafVg2rq/XO5fRkMRhsWBgeCgMnou4tIt4+PZNGzSUAXg2G
BGaNoiphmGiC2LJE60YZ9GuTW7lihlPXAnmKwg3pPfvTUt2BJoZoPe/ZockfazTz
5anTB8CwJr1X6Tq3cyOUsKNlwh/4U9byqZ+umbd4Day6zzxDLFfFl43MGlEvsbs8
Jiz/gpzjABn2F0JoBmM/lQG+utkFCRBEBjUJ99KIRnjjGliHUOOShRNAFqpaViIo
Tu2C5Oi2G/ecgyWzifIfEILLa9Hek16e38i+6R52n9BxoRjVF+DLTdGyXPVhIw7R
89DOyuGRonqiDYruckbIB72ZW7jvTGvy5ktpC7U5e4qr8q+ERYdLxCK9XdsMxZXu
3Gn1cWPUFLmurQTOCwfgA61q6h6Wem3VVjXmBbHZuH0/J4TBO3MTNnNpsC6G7irW
5TM6TLQrafIke3uFBfeFp55VodlplcK6JbPWQVYTM3TXOi17nBNOExnek0euLQoD
AITyIxala9kvhOWEzU5rRbg1+VWGyYBOUKz0hYCTYnwDuRi3EWIsLB8WEU8qTd3w
Pk3/+AwyB4oYZIpP7aB/XoW1Sh1sgC4jSiX9NwCFXkuBHjsESt4mp4Ynqirzjx3F
E0aRMTMVCKtn8QoMDTYQ1LEzjgGHdhRTNognzB28omEKmLBGdtI5asdKQaBA5rgI
u9/vvO4wtPxAF5Lv+BfFKuqDduqjS3erZQw1cnI/0ex5Y293Dztetyx7LnxLrGuU
ucqH/JuRcCiI6Gsn1TO/yJFjDt+NZ8864U3siqZZ3M5QOZGKIBhpg2/+EBPBGctO
QEF4YJmxslhRUSBjOtCvXyFmScU4yevXx6l9S95CHpxLx/LinXSjBqbktGn9RWa1
yz2s3ZsIHatZwWm6k4zOKHr8pBxyjvxts8IKeOWVDrur1BSVic2ZCzSTdDA3sNA/
1HpzhHFF14X3iF1REn8APFL25nZAyjRaJfD8sSoiBkB/N6RLHglSrn3Wq5OgFp53
Bn79wzCmvDtMSXkPW0rnQJCkTN8mDWjFmnflRkXH06kwNWUwyObLrsB3ptdq75Vw
u6K9fH0vwZZtfPPwhbfg/TXrh1VYj06NTvIeh0f9xalhDDJjheErZbh9XAnRsq/L
knqJRbREW4XbbhZnh34kyqenIOpg5ka/HrkpcwUUK1h8HlF8YuE6G9OhoH/LzsPQ
H3v09y8cDOTXSeFrTNrm2Qw6DKNcnvqaKGO6yv8OBn/EaVYRmIWDR7m/wGcqJIG3
Sr7VB+mw3vw+LR2vZAioY0AaNHQp8ho0GSxlT2hpBjxErKFtE/VpJz6yfKb5A4Gy
e6n98QQttVBOxT5VCsDMvDj49d9Zc5/4xcDFex3Op2gY3ohLkYHriQmQ/fTuLXKd
drQKHQXEHOuiohj0R80RanTlcfY9eDH4Hz7WgLZW3VsurW55tan+M6OY2RJyeycy
fEc9SATzCT6gq1NX94wBIaZqd+pqDmYD2WOg5KHlNGINNM86NE+MN57XU4yTRzyy
/mgIzpcjQPom11UvLVodz8naFe1Ce/p8kbn54B1CCL615uuDqAHzJ2SsHgu5czTe
4R5OWfRiuEAgmXAqijMbiCt3oR8mD3c4p5VlAzBUVaUhPDqO3uaf96Py7pEf5UMI
LTimaltOKHX72qDQjc0ycdTRd4/oxLtTsKb3Utf3IvTCKQWDgBM5ekgNG/Rp0ZQH
SO/67GdQmRTLUK+WcTxGBaJyQGc7j3LwxcC4vjoAGs7qrvzzsZ7DGCOqVl5YZWAn
7nIPN2X8u2Mq2ScKksQdYkh4kLGiT1YcT7ejG6nwxnr7pvnK0CoE6HLumuqv80dp
BivcdC8hg+Q4lMMv5MEZ5AjzHMj85OL6jawrfem4vYFXjVsXFE93XTO8pq0wxNf4
qxhQL9ptZhGxT05K6Sosbq2L2Mpo8pCVowBgSsmEJ8y3EyUZmJI+dJaq1fRU9xkf
vbcMIbxt2j/VmPQ3mcBoRMqgTq9gxkmc/gQSeG2QNuVs8I3I/YbgdOguOSuOsuBd
j9XDD9n5xe4E0PewLsmVCWy6pjsoNctkbv8pFD5HMoZDNaHaxxmdwmK/Z8zMddog
qeKo8mLgoScFCguQ2y9d3mvbq925dw5VwSz5CBGBgtN2eCZ1ci8o53F2gymJDFGL
udRzDIdFYFXbNm/EyTzTX9SogsWLt7xo1VwtrRYnwUoy/I3KgDgtcHnvgjeMPqjH
V7cP2roriHU9w/Tvv3lc9BFYFC80hU1nWa3gtyBspMc8+gJwSngmHcOA1SawB6Yo
FA+RKaQVvUR/gqbShRlqF3o71+Z8CWTLkLS6OI+CsFrBbac6pIbcLuQxM2gw6Xzr
YLru3OENH3XdJVZ3EDTkKBm9aI+ebqX1++CyNn/VpzWH7tgWo2E1lfmIUQumUXfl
/5TaGRsSsWYipUolHv0cdW+YXzJNGXZv30kdSfXGOZrDOmHh7xCttBLFmOtCpjYS
7ZAx2waJzoAtRlHOwAj35aO6IU7QtRDleFkRJbK2N2om16ZYLcg1DmbZ8O8Yb5HS
LMXyVaQwGbCjZUCDmXQw1zRIaW2Mi78xgOXODqBLgKRodDTVTxwgOwl2DQqWA1Bw
Q2azD5Y2MOama1O8ItpsdLP3IiFkOIQRzCoWHsB/BcVuLoot5T+iVDCpJyQG2TqP
J/aGmWnqLyBWKnxeXnaNpA051MfjBgwk/xUgQa1GxdYdgJlMFtL0u1Rfruf9/7xz
6c7R+B79ZIdwqv+5p83XxzOfobLXs2uiDlU34tCNP+e0gPzch/IJc5xPX3nNsVAs
l6mdEZ0+oDvFXfXW4wZe3gRYpb06NBbVfnK/QKF9oROnb7wDFz1hcReDf2QRCdqt
MCkunNVZ61wng6MQm35jCooGqaw8Of+Vnte4RWdCpUbQZpTv74fcTqP6V8/fVU2K
uKvsncJjfbcKII7PkB2t9V543CW3KHYWm+Hcg+mlyVQA3DKYygmWQFuRgngbXTj+
jPiesXigThb1HKbQJTCNXQpXvYRwkrLp7h7GdTC4pwCl4x+wOwsLdXfWQG6xdTS5
KMbzdg+cKB5k1WA+eZbU85TNAz+f/rg7YFw1pqMoZoNYm6JU91FQ3EnwOg3fmXHG
dxIBZRIJaZvHzvuiJaP16QbydMw08O9sIWWTj2R1LQ7pD7HfamZMUteT8Co5aQ1y
S0b+XDynGBNg2IH2Fk33l6bW2bmuT+bVrpoe0kp4RNwcxs1gEn1i/ym14559BK+w
gGrwuRGjkLwG4x89Or5mjKlCcBH0/H6ySXPlKOsn9jc26czq4y+BpGD89p5CLjA0
eFo6o8aOfMLMdKXnLFjlV38mIlKs4gxSJfQP98iPYJO1PvtQ8gHTrq3rMryeKxZi
jgeJEEVyPjkWoiFCYzygO8/hkQjQ2QhkLmv2n4vmIYFWfYPkul7oQZF3lCsGdnNj
l5GIDc2Es1ZcEyHxSTUkqAprTCQh+QYErMNhDsWBdWKFWxXa+CFRMxh9MjoHUiCk
to3Fi4drSHR+PDd69RAwiqJaw0AsRq51pPlEVvfH0CjjM5dopFYFDOEgG87S11DR
wpisGjQKRROdXST4362BU98Zvjas0w4XHm682UEOmjvSKjh3/KNy05tDRJHzFJK+
EWMobrTSjxo3TIpdfcn2bstdp+iSR+u9d2apxYL/ZC4+c5hMW55kAAdE2Sjy+srO
S+dj+guZjbxeuRB/9WC24syv/T1lZyngFRmt6g35x4xoA1+vOe3foNxOGn+WH1f6
8CCVcsncGDbfjXSgHzrbD4CrOtMvPMrqjN8GcCtKLbnLR8+wg3RXgqbOL23LcPrB
Js7JtUp94XTlkJmeCS9IiBbloEF+yMaPk8EMDL0tL4rLwzrN6V3mM5n3fNQT5v8P
XF4EwX+7x7tFgUqLzqHCAEOhe5Ob1KHcwzjya3JOU8r+2FHsCoy4kldEYmTWg0Ft
HtVkQfTBnFG6ofjgR3EXbOx3l6p9czk13YnVwdE7XLWBcaLAS0Va/TqrP8YXpu2x
rhtkrlS1bEY5iUaK05v8QePceaXuMAnp44x9+1hJevBHz4u+tdu3WPn/PlKxRfZs
IN/prAQUIXmCufzllJzQ9TETJfoobsOM9Q+WayKIBCpbh9V/nJPh66XdA9JaNDwX
rtLO5NCL02qnDwGRDYn9TMzXeixWuLuSF1jhYqiRPB7NSZWQvhcLNi15NWIRy+rI
Fb0w9BEqHv5h/4HxomZ08Etxc6yIRyd5ppGFyQDaMMo8zyKoL93VlGcE2gcVaJd2
GLhFueUYaGVwS/rr3ki7iFWmGeEaGHLuQOtG0sKV/WZxaeV/gosoWjyKwT+ZuHyq
jg8IH51o0XDGd9f2rrkmyGTiLRg9rCQH2UOG6n+ErZKKD5DP2uP2rP+RIoxwEFi1
raMMLY4X6qE84BtWB9V3VcHGCii3lN4hX236GROp1JF7HA+cN4zkfpcRiqe7jWO+
9Vn/uDf+fKkEwaZdGJfHH7PB/X2urTc6urBlxr19nLw7yXI9zm59XI8yCZrXQutI
TgqtkntHFBHNQ24vH77gwGXSP2Ss8TRPKsTUeBMorO8DbeoovJFCACiIWPUxzC4L
+U87d+vR+K4BYkL3ecA+EfVk3osXvfAVhfRaNSBrzim1/B0kK8efQdgTH8j1dA9F
yjIJ4hOZACjwZ54kakmk4BG4tYA5lPGDDTwoA+UBn884ye+KrV84jAuoMg534iDa
wrTK19W185PLiEUSouwBZaNe5VxStdXEvhfn03mitFXKq9UdRB8LEAYwbvGcZ3ve
ChBeVW6bApsXiVfvWMKnDYxDL//pL0v+AC+U6Ns79ZS4a4dnOjUt1HGLJ4iceHC4
Jo6XbVbgwru4gkIZC+4TI0NEyf3B6MEn/98k6k9AUAIJ9KeZc2a4NMlAMR9PgNMZ
MUAY/U8b9oMW1HXefC2JARb4rWIgqEksDV4bhUueZfrc6SvHoYNg0fyOCpTPHAYF
9UAw0NVI7VmOZ6R8M9Syy1hr9iZj7kKcscx+GF2Ibenzd5XCgBP1aluydwUb3oZW
qPAawa91K7tnrHTaqLAqQGyca2xZRl+DcA4NdVjkrY7PnmI230DDVwz+hCk5CloW
ooRBNct59Zt8U3K/3+1dvVIFgQUu1P2K8Xip/rv3wUCFKkd1ezGjzL3GXI2Js5CI
cmRxIr6pTmv1iRYEnY1XXVoJpLZBNfAMqwb173w6x8/1KQzugulKJog2O4TVZ4Li
qNtcrbqwgrFlJc2DFQS65A0uuIGJ+/f8QP8a7rYx6F8nBgVsEskG+3Gd3FGoba2N
csrpSPFfILPAgxHhs6klBnXtZwlfckLKXy5vZ12j0PoWa3mMAbMZcQfOitGjWtrB
6W8wkierl9xYNKfjC+4zKi6np1lCJb1KwOMO7d9rvpO6qk1AtZHpv84hhYY5Eris
CUEScXlE5JPvfi5l4FOeuM+NYib/c6Jg+I1/ue0/nYhWiXRx6pbcmAY6XbJtbj35
rTL/haPCHDyNjGUk05mY+6vhafHlUrB0Y87oHQH96Vf2m9tTCAmczbKj+x7IWUMy
PNPYoxqJXV/lSRfPfh1uMnuaH2OXYP8Of4Sa3NtFFeAhE4O0INzqYzWJ5mdGZgxD
jZfkzGjDyFmElPsbeKfa3hOw8zOtV+M+xMZkJPM9aFaUIV5WIeZAnRTXr3dgnrPW
SlBAJVoxK5smy6+CfUFFkuF6PMcEJb45Rre/ib2njCjyijCCjMu1ljRxvqbaeVv/
gwr/XPMOKPU7DtE+nj0O5ZJMqzq1pMSo25mAnf+gPG+UaF09Fb8Oqk1QilBb8e3H
1Y7BT89sGVXOZWjNjjWUyrPyhQOdTEaRAVaY1kdnV93B9CyhTQHi+5teJ04/38VE
VFOrXRmE0TEZa8ILmhxotVkYcip9usAFxKvE+JtYbwzB3ejdaiBVikkNgX/sgBhs
yCv/e2NsrlEvTmQeGe35uF6sXNEDoG9MUsR24y7m/J7KQDTK42jnTyCsHm4dxzEV
T1Vg/HkQZEMfHGMYnJlxa0tH6B6vYAhE2mrXT6lagPr58jn7vhGZTaGtIqpyMNqb
z4z4iy3Yb3W8CK00I9Zn3RUjsk7k8yQBMNEPW18AXjVVWUTdFRBd6X5Kk7jWPiMo
L80eFNbJXiITJZp3urIZtXToSy5SW0cpqQLtLUyBHSdCwpnPn34OMQCmQExsnRsX
89ZP1eKA/GUl58c8EaI23CGHW5Rd9Ac2ybGqXxVH0oPOAZAUlWKD20ZT4gl7DEar
wI5mLdGQpr5WeJx6J+pPf6vXwTu+mVOd9Yiv43vCrS0uAL1wxeGQBPxm3Xw4wGNS
qMA1ayIbs49aB4BOnajQ18NF4w+aX3r/LAOmMRwLajHZVHbuRXZ94/XoclZSVC0O
QK45ByjUxhivJPpTVtRTC4fT2Kal7qGja+kt62LC9621vPlmQ+WjPlpm0hidd0xc
h/cPfQCGsk3KaClEGmgX/j+MDyZge+8KBLjahl2Gpdx/9m0UWlw+SxqZ1US8qGmp
Gw97quo5mf91wWUW+3a6zvrZNizKCipdZ8JdqHEKuHOz0Z7fl1O+aQl4pCjoiXPU
Dcy25dN8XuDAwsRouCLRRzYdNl6YOUHrA3fxZ/B9FzM8jkL3MJ29R4poqjNV167J
n6Dj8Bx+cBFmbFhMJyLkwMCy/ZOVdOzrLOCZnmbkmpj43EB/+0JW32wUPPTDQH/2
f6HXFNwxSXwn801aLt1u3ezhC0IUBbPVAGUhLydCLUktfq3yJQdsB7KSCu4z+nP2
i7EsLPDpH712sUGrI1X8VpTVAU7Cbg5mchSceWXekixH6b00Rk2YtndtZGW2uA6m
tiiDQu0A54UB2lkYqb50NOF/xxKzK+6hwn1ejCFVwqmxRN6wu4Trge8H/ckPpD76
xXPq8iuEnOz0GP9p/2xFddxy8oJsp2d1j9WEv2wCWUZyO5z0M8ZJ7p/pX0xDyWW/
GLqqqbQVzJNg98U/cpevgQ7kIIlQYiZi2aTKW6z64nlt0w6H4ByQAFClKikergmg
MZ5oIfvy1ccNDxhQ4ZJen9FVv19MPcyxK3QjjTokOU4KN5NsA1/djqPKCFiYk81y
2t7DTBa0xD/U8dwhxLQSVaUQZs0GNLm4icStQ9eeL/kDQ+TIZ5a6A7M1nFQ9sP7a
TctPuTgm2t2pFRi10/MybuV6SbFXqi2R3TaY1JufCppvP6FB1ZXS1p6pAOKoZbd1
ar8Dkj0E3FYqX47rQM/fHZYyY5p+4S0xqFEjZS2xcJ4mQJeYfEcHhHfNK3BiJ3wt
LZr/riIYKViDPSMijW5j40zdFmZPha/1K86pg5c4EUfmNWT0K1Cxn1Fhyc0zKtoV
xyq+LaMkglpPT6rL21mv4xNJ8a9jBzUkLSmi5gEGb3yJO3hdfQPMh88Nr6jO8piy
YCQ4Ovct/hLESRyK/UBZBIk0mtUisIK87XjfoXO91T3WuaPouOgZjxeDr9FQAV3V
B07dzBhbRd4xQ6cEORJkoOQyGXz6EsDQ8oKO/uUk3Gnm6ZeqkVRA2mH08hHwaR4l
5Jd5pxlZ6obcQePGpSXQ33hw3OHABVE3xPUJVZprG973lS6ta/240gf5vnSe8It/
RRO+E1ViCdEp8JPc8TlA/vkkUhEPgxlAwaPHa45+g7/EJX67LwiCCnPmgOMOQa7I
9pguZI0fK+cqTmLdXeOKlMNGT5WCUa5unWqU2JDEmlBZnqMvFsGUFH/eVAJ8U7hn
7CnLhmEFoB2UhsYs34HtblJrtrybIcfP4jbQe3NH66TUSJP8FvHg9MqeyiJtfOBq
NwN9jT3wxuReaLF2UY9fGBH/l0b0DhGEBnDZSQ2ZugaQeYccJVzahCYfyER0Sbfk
FuNiEHFy/0KXjdGi2YKV0YDJaKpiMFlDuXVJMGyB3buhEdRBYHyYAYjdFmkFxk91
CbymmVuGKa6ND/KRKelgBJx4aNo1omDwescoLEHy0cGQmK8YgyU73tvtQ1AG8OzJ
c27TDWF7NgBJsDAyJdq/OiC2BGxIKeSsbcueKcV7NvrH+8N1qxBvegR4ZF+Ao8Or
LtqI16n6XKZ4hy7xeaNn/Q5cyPg2tnfyawy6KtfMq1m/0hG9yjlfuy6IeLLpe3tm
iwpFMxckWKl+hBACfIPzOC9Ab3N4lpnI4oV+W7ELkBuw32Z8F12AV3aK9KUrTVqQ
BKEEKmhT+NppWd+Iydbsyh8QJ6ccoi0A5OpztRDUVyUxQ7sG5OI2WJOkN+O2Sr7F
wu/MIT+FVJzMwvoRfSxGjhejT72V4qfLGjv8oO1aegnKKocZDcIf5WOUBnqSMDW8
NfeaTLYI+HlnPG2ASO6xM76FhyoROeYu+pBGesbA5Rc3riq/e6SDjT7W+LYNewDE
fVLXsNLx0wDl6WYQurX6h/wEV0PlyrauTTc7Y2epGH6yB16m48n11I/XY8oSPodX
9wPWfxcXEqny/EkGxEQAroij0n2tDjFgN1dAvLGuyL8QoZctbge27zH0AByTOOMW
bhK/KTIv5teHGytp8DSZRtmC2KxQCmnB8VzvAi1aB7rpkKdM+ILs7uXBaLasGnPF
/qtKMJPlzdociouQqBvH+uVgNB1R7rNFuGXI9ckuU6RXtwhB8wDsWAlwLkKaTbtG
DQDc8INHx4aTpz5iSthk75+AAu40i06+6Ifoxk7aDh9mufSMAjPkQGKXffJWGBd1
JsYYipXAik7dXeaCpTPM49wCpjMpw4vfpmXKy20GT1kV2JnR9nWdgoCKw+TQwwbb
DJwpl4fYqfqw1PuXbgssEAbn07q6dtlfKxgXuou8zk99upcw7wnDwri+XVLIIEdS
GbeaOqAdkkOvRT01LFyv3rMRAwRl4blpXoMVASpDvacdFTLf4FiMHH+B9QHQUps/
AUqUySMclhkmLQoaMwRq5pyLW6l02e/MqdXzQe3o3r3CclpNTow83mh9F6btxVtD
XP526xnRIH+lrgrH+SuAHynhD1MwSRZYLiKjw+w4Kogo11Ba/5uUJogbnbX1LKYU
owFNSXlfS5pAqh45/p7EsreOFqwOHZvbAZwhL7Rdf4/CEufPvLwo1Hn/3Nhe3Vzh
pD8rEWq+s1Yh88e/Tn/ay+QXaFc3l8DzN7zJtiPlDSUW6qDH2Ie3vvsIYojkdRZx
WUNaBTIsvCyl2T3YfdI3li4x2M8UR1J6yzT82QQ93WIT6ZjDmilM5n4kZdhHpeKu
5kAETIZVKD/QT+vaK2jFVQhlwbp3WyVjoxnd7DQA7aykOR6XIsKHdBkT00WCs54Q
gdU1zADvAwpEOcfJGNcFr4arHiiQuEwKwAFHVGiQv7+/fyS6rM2PppQIlqdCBqqg
yMJ10ErYyMa4Wf63jFoPgUVi2r3O6D458g9TOozGnWocvhPtbHFAWYzbTDYVTN+l
xLjMhUsAIxaLfkQeD8ykwzjhQJeOtOHu/b5Xx4Pd1+o4MV98Ydv2Pstj1FgH/jnY
J5Gtsp5+c9hX+sQSbf3I9MOEURqHiZWeoW1C0gpIETOH6pJMdJjD7SKJ3bCVZh4I
+Zr1OgP/mPu4Mr+SFkMCQ/rlKuD5ibiicsv9VytH9tIDMHsS4wquMb9ozjGtzARG
hXjPG0OQT6PPU0G+SQMQEiQgruLnueGXICSRBEOmarabq/7KCA8qVx28pGgc6XGj
JIfLg1sMqIQugRZL0NGsukEJ/NeHaeGsPAe3u8RUlWOCcxdSyDlz8+8uva51QuNT
/Spj7rxnbL0Fyb4HEzePLWteW18JJLXjJYsKwp76NjX1Bmo7RgrF7L3wkdvrbZ1v
TXIvWjl28eV0m8A6vKWFcKEML/IoVlcb1LAtfwX4uTN0n/jjpFDIi6OOa48lcdlE
NJXqPT8nsl4vb6Z/lTlFGdw/MAZbKhR0QzdeWZI20i/4XY+3LiXqFcpn/HJ347b+
QxDdbm/Pg8c2JoXfFc+3ckZ5/NqV+x8aiQZTcjWEmkg4yvS/Ujn2doHmnV19j8g4
qA2BaRrcyT4jaR6S+snEOdiq67ep7a3Ol8WLtFGWpptMfjTucFTaEynPRBEwmoy3
kaE62MeC3eoqsQwHtLeGj0QJQC8bex7W2xaxrQ9yxM3Ss2PWnMYUxKE4WLN85IDJ
++hiXhMxTN1y061cJfaAwOhFKU4Az5x5pbv7sx7YUeHgPTp2idM5IistFkdwfzWT
IPY6i+crlr4HQpk3F9+SHBBmxSvfG9S849WfbxUjIpdjfL8g/IYATOrYW9zKPtlY
KFrnQEiJS2RjuaofSsFSub/0A9qLuVmO/09bcXlweGp50G7VViwJ3Kttu9Pm6x25
FqxivDl27g2cgm+QDaMifCDgjGVNAKV+PSgdJen6VDbO/ijD0wVtAmPYkJFBGUDP
AnHiGwQU9tmv7h8I3IZFoLqBu8ZLWJvgc+7JQ0IzTwpLOtBHsiYRBxPeyLxRULYT
/uNvh6eUEod2ysj7TkZxueXmGgtxN3GH29ZqrhI647H7LorTguNSDeNGNBBdXLWJ
BTO13JZ12uGJn71zKcxNtBmy9gVRKM1j2/U7p4K1iB/0WgvyX1ZPeowrTUc/KjA+
WgZAvpDD0DuAsRadlyIruTz1r456Vri98b3OpL8G35c9Psy4AGdFGESUp8vwXyvk
y6incuLJWJlVc70KGf6ZA9fusC3CgT+NlFs24aMrJnGkyuHt/rPIpONqKR92JLHu
NfNbWgbwvE0IYSxmNLo36n0Q/toRwcSe/NTxVKnrA1SwqL+qOHcqUUbeFMPUN3jU
fB0dNt+oiLeBoWLF7uIOh14x2BqmSCt097mlSpKcMI8Lzbl3vXQzzBog9Y4H0qJE
GaFMI83/aaKgE0TFzw7pi5/Wk17EcuBGMO2+xsZbNEb5CxhLt0H7QkvwBkiugqYq
dIoxccZLdfVjSKC5yPYglE3QwTeWF1iBqBrecOfYaCIuQMG5AnpHTUttlhctHDH2
1Ly7YzWIAHbfqTtk606BzMZNsFY8EKPxVOnyI9leXI2KBrBz7L/IPn7qTJJNMsDY
u+f1nRRFQuGlAmjtdnxnt/28+mvAtp8gM6QmATqXyfk4+YxDHTkK9wyoiUmfaBRG
2HyifSMyZLUngztp7TSURVgS6tw3xo4vmPBs5VZpyNrsfvL48duGZsWmWh1wIQ6i
1gmYy9jf6N//fsSAPCCPPpFOM5vvI9ebBGzaDq0MEJA3esLSMikFxUWW2JFvjCq6
/ZLPS5XbXE2I8dSBxdUSKPxhEbPGc4vVXMVF3jA/UNTjqKe3nAUyvurb8OJu+Y0q
xj9xAHAZlBAyvozNJUx4daxSmL8SzsBDzPKUbhvS3yGFG4M0nwxklxJdG+ZurU45
jT7Xr7s2yQl4Z9TEFl7g7sCqH6zYhFKZgKWOvi6/PEdqlaW0tow5upUe0F/zz+rw
fpEUyNbTUuPQZdFwFFQ0Od686lSndU7pbqJIRDXF7KAF/Edkc+PVLgJib6tux+Pn
Da2hN1PAgm0+tmyZ7OpjsTuNSUa2zHgT2uZ2QL1BGOQk0J1XqfCaFsUA8uSdrgDA
21NmeA+Atd6qcLVIee36Ztx+7rnYa3UIyjvtcejZl+SUCATlfWYi6Q6XXhtCkzLh
JyZyPThZuTdDk6aBXnygVAv3fG1irzwcHD3UC/LMgJyyvhpgRa+qoBNaH4tNuXuo
OZehcsH4CbZOO8AgA5FDr/oCfjFNCILeTtCKGTjWutvY/0Fryc1ttZIHQDJ0DEuQ
RaAYhHPbZvZ8RAIUD3NiMwZjl0EYylkCweO4FqIaZ7cfos/hsuS00ZaMOwWkI1DH
+MPTp93hEKi26hcJhCxLaeACNs5ZXeL9Z+PK6TKqM4hyXk9muKvYDdhe0P7u5tBG
rbIWZx6xbUKJcvxKBrL+GJAwCntQEGRH9A43Es30R77UJzPfnTaDbZp+9raNw66D
e+uXVWFs/fcd1gaQ5ag+2YDDGbEDLX4b2A90MB6ZARFvo1V/dUlwBVcHrhsI3WZd
itGaI6k/uq5BCGKlKXB3z7qKyPPW70aOpFhqbhATUCA/G66M/TJv8mi2VwtE3yNY
fofEnc9gUc9ofsgr3XyBWiSLrjlF666R2XDMDVaBsBl3H5VLlYPBXu9rFKq4S2IX
Egk+xB3sZ5srAUTuLqlEUA9XBC7j0JfMMXepc6xDpWt1mdIvc1q5wWGJRhvJ55bY
e1MoZsysSCF2lXPDl9TPVkHn1JyWf7a4z8T0rBHJzKLeQPqx1Yk694Wa+JdXzaJn
27Acib03sONOkQQOLfeUat7j0d6Ezlsi4X2k14kAyYGol/OX4csAGkexIL37tRSN
gonAXGsPdzouYMdX1+/e3RL1RGloolg6S4EddZ1+ChfbV7eGinn64RZN5YnoHpmS
JeMia9ibCvNmRr9H5z/TEmIXAR1Nq1ngse6hxpoy9hUGCg5Si86EPHMVAxrPPE09
eIjAAIBsWj+usz43izLBi+BtJusPhCPrLVLU3Z9LxggADIDJhSoUtRBzT1+r/khn
UXL8o1tieeY8j0pQPJTCzo/OgCGpa9EsqKA8MoGgY7rVDIW9l3dY5/e3hdY1VF69
eGNlt+JZ2iedeJwr65hMN0eBAxFU6tegXBZrBKjcMNg8pq5qHFKxoCxvqIjaYce5
2uvS/Ze9vimEhE87hhiU2TN0+LCJEcILUOVPwve4d7JpiKHMdV64gUUpH69ySwBq
f/0bhGF3csk0+3QGpPzm7mnIVzA8MOQp1PbCzlSvZOLB3aoqSP3qbGmI0E4++8yP
lT85qIcDw4JxryfYcxfxpAcU4G74x6fMx5C2mbVMXdqu1xlMSYBgDoDLtGEmIZzI
Qd8UZk4lEals/Sn6bSUsE62JxfPxSfKrbn8B2WUXmVQKur3PiAybaL7sFmRsT9cG
NUM2Mj9fdfe6ok8vpXCHuULQtXof1u7vJLrdDWGAPT5IC7SPgZ0X7GoH1DPtRSSG
y4m7scM5Vv7cb+814s94WEJN+jHYRVAeP7poJl7MFLV6cFWDqcgWTic1uBJ2N4Ji
FEFF/fijWhyeqqlRr8BIOxMOqG8ju2RLTnDjd6clqZ5mL05RPKrqZ7BHaqHFPI91
87K+xXjNuXW4okjjvrd5UtrIAgj70IIc4tTqQr23WYvqiQQGZr+vYZj2Jvk4bDbp
GLVvIKZHE7VSDeeoUbICyDTuZAhgJqne/DLx6Yvd5fw0PcwFzMo/z0dEu3sjqGVq
mbLVqw/lLq8d/HJx84jFdrLgUSwBRUx3okNQLWhKf8JYQL6rsFWpQQowJKHc5/a/
HaPsTc2zFkyEINbDe98Wv+h5VxVwjst8hspfF8dSxGY1K3KeD1hwjP99b3sRfY7E
SbIQwZHM9hYBxhfAcKHob/NAisKIYQqm+nBWEEQnYGb42b1FpYHWK4V+FxtUHdRU
fWxnl0E2XwdMZcRlAZWXUvWwsd4Yw+e+ihKf0hKBx+vbJajun+sf8/vyoU3RU0+o
PRlJHVytkR6ZlqSBY194GSzPW0uElKCe132QAwE6QZjutYfxZIqoLP5NcLcYc8VH
fsuXhtuijhinxu2TgvOvxp8sHvm26bFe2bzPdYuyfM/hzKSeTvk2HfzQkfKFjAd1
QqPN4vessNTazD9gbG4Ni/6k1DciArcvX14MfGDWmZI0NlTYxOwhjrjupJCFbqRE
LYOc7RViUCuwVc4uSqfxI80M/HFdw7WeQ4Idsu+uyxIB75C2bBLdl1weTG5wYJyl
Mysf//wlV+BHMmeA6G7DqaSPdadSjVDN5bHSP+JzrSq5jqkRZv5sil3cK28zhhH0
iPewRBIfDxgXVuNjWa0/ds3QbaYzSmiNPYX3zTxOymFYljLEZdmYPw0ggdWLxuYD
/nN861QvJd0se+tQkmXqbl8QHNQT6tz7LMfke00lb/luqXeftSiSMi+oBo2N0WRU
sTHragRMkU3kPs7VUw82SloN821AxS/AuoMRx/Q+ZZQ8pJEueHedbrUBDZxzWXdG
SawMqTmw+rgjol5UEC4qdxZIDysI9XBsv4CWKBpKSF+URzyvIv4SanIfSfUqzagq
sygBdoAxNdXtOqkgzEwhMYg+DYPbTzl3j6eBJdaFRemYHStJh2lNoLNrJtyb3gby
iLpS7FjjvgWa9v2bpqVWzsF1BXsCvVw9ak7TcKDfWOAoTyerBnWcP8lJkbC1IXJ/
ZPuvRa86sR6u1Gd2+yjaRO5KRDS39RgPFyOS/1AbMZDP4d5tTdweZQk6+jBORuvY
ZdmfeomJnqaGgFTAGOIOPds6n/PzUUTNNmkNS7xoD0bj8ENnOC9uwqoBY4FGh5eO
CEeeasLL0jXBiv9OrBDWlFTvKxrcNS02jt3XZTOiPYbdb8HhtR5xhcGAv6djBxZR
R1Sxvo0AuSR6kvnYkbE/krn0mDYhfcBGsh6GZF5mKFAgSLXW5JxijF306Hn2mEzS
89+g6Ls4lbzg5fxyUyeZPHefZgbwdPtKKbEa1vOQ5l54PkDcgmTioL5CfBkQWttN
acD2k6ZGiufYpUp4v5UiK6xfdqO39hT0R80Q0JMvAk83tyRlJKlZGT/WLyhM2vNR
Gz8DlwOfn/hpJwbY6/TWrfMINH2cWDgnG6k43Yu0lErDRTno0uh7CEI41ftzmAYB
aPBkiFazXlJCs0uPXWRMtg3vCdGWn4ptiKwVojvuSi8p4y3FSrIc7IoxoBS0sK4E
Etaufas/HsxKhKmHZGNtBb5TPmFiIhGILe/iWumMkFk4tPZ+DOZ/liWoZjH3hzNF
2XxEwkY4T3lE92M5kBDFpkEuV24x9SEtW4A8QT1FiD0rIVeFbRzOjTXnf/Zpw8La
oYW/nOXTqKMWaYyyGvl/Lo6w554PneJ330t+dtiBXRz7uFMC4uCKFiwJvfv5R5E4
JyxQGBWRECkSKCGgYbJBmDCM761jGkxq2hZwp9UR98tM28OZ0z+mGsM1HkRakefm
6d7YpGsQAuUU9f24SmvXl5STuajS/aH4ouJDQBOTAiww/oIWat0Pq6RSKDnJDQ7J
iwtn59e3iXdem2GKKsW+87AlScoovtKlAXNvq1ivDXWn8m5jYYGu5N2oeCFCsXSh
Zw3SHpyppBaacQs7nbu1Bw47zrWCnRs0aGJnrHo3fvhPbMTgJr91mR0JotNKl31k
KiMHEXzJMMgsuWT/JVqusvM4Hmab/f+MtEJ3NAuFx0YwWFvlJKhpNyk8af2f6ZlM
aE8YC9JvXaVkwlT2WBLul3uP8p3cEwkEwzjoITY1OC/klMNtiSlt5ojeglQ8tTr3
ROWfB3HRPyPM3IvPUy8lBeMPLfgIzNv4FpNdd8yiLGdIEi4JfyzBXVcx/OrXY7Gn
oI5l3yBArx7wi4Ph1LVuAB9PbGIxZ6FVLDW4s16P9pd5tJMPiKeBszzc65SS6r/0
0YpMUvirN+hbZHJExlH+Sidjt7kRf+dJrWBH9bjTr4nv3Btkz+vtR0w4ktiOeehZ
Y22kSbfv/PaG2+JU2Jvd4XgJRQutSzlOJ94zEkAm4VJ+jZhwGR5/XWG9EbUjFkh+
y7howxDoVeDC8IEuUqrq9UBYgTWvYlOkctkqV/mwGoQUrMbw/wmh6h4tca1eSQ8S
bzHeWuIQ5BO04ImjvU6+fXAINjswm03a2kVZxM2rFi0g6KBcQEcq9tamf794GFqn
AsmOd/VLHrMzgcIRVPghcpPqonaoCeq7SYytcWRG4OgqRqUfuZcyABNjMJesbE7k
aLSYNtAxtKO0uTKs33lysxN++zGV9ehJTGaazLsb5cOgHg3RNp4Tcq5qtyEACVR2
8sR9aurtwmhx2orrqZByd6ottRyJ05o2WHS5zA8IMkEA+mrC63cSsnlaKow/6/jN
5n/++RaS4ofB55OBTGKUs/FBJebeuS/QbrHnwOWtMPNCJB5Y7O42VSeigsa7NNCo
NitF+RsACLwsdpgzBUFj3DaD+Dk43CCUrkRXZJzu4ZyfoDTrlaltm6tP8H2ZBDDh
rd9xqMH/oIYK5j1EFVFr36RCQbZN8ULw4NBJxC6oi3vNp02IbTU5a4VQRHvM04uX
BGcKKSz52lifKTraapp7CUIDbpKxOCAFB+1LanJecKr3LWOEc6sjaEAZEuqBaGbs
RxGfyzrsObsIKT4YvEmdql2byQsGdIECz1RgeRMIkceGdaLKQe5d0uVgkKxVvf2M
WfyboFUWjDmgO+omh4Mrf/b3UFuFdK1c7Jxx5qI96DQi1K3no/e6LmYbN0YzICAW
CKIxHv2uzcYdfvyboVO2s9kxvjaPt9uCgP+fAjXfDy2G2pHWa3h5uimWUBz/VJdn
26nQwSR76xDteOIfa1dv77/WDvW7t4fRum5p9iAtYVAKpa5dY4QXmQkWTBW1A1oA
i/OmDvOwVJOvC/sApupZ7OLuvxHYHigyyGBkaX0XcrtaYcEjFD0guLbKpqtmSk5k
EKD2VNk3GCrXGhkPS7k030C1hLUuHgX8TmpH5jQd/AAHLXdvJPAjtqzDiRqQ6IeR
P+RfYe+vsbhAjsmMAdSCJXYFUapWNJO+pHw5NLx6CtWNFrD89eUaeNP5/9O92cXN
ApwymVIVSFAdgJdzEKnC9+XEBwRwiAgYA2Y2jITd6VsZ4VEUrJCe3wsR+yuHDiiN
+gJKeOE856e/3IZpGsa+VyzNdOJh6je80lFqNL8asMCbISuICDA2NbYdmTWyheCt
Ncbj4T4vOEVCzfM/CbxDzG4LjH4aFMa2Ombq8DCgeuVtuWIDGdgu5rbbK0EW6x9h
aFinpmqlwfU+NEY5GdyVRg+7H+xWFjL249StDT6mkv/r7WS0mcNLSIGWxHdJHjUV
awOZljBDjZrzK3y0zYpLYtNfW9pvoZ5svE8yFCFdI2BGXkx5Lgp44M2CbTFwJlNS
lQK0naxpg2LZIM6MpKT1megIf3EZafcTrDIN9RrWTH92BURG5Z/NmRbMdn96otaK
6ZuKeSPwBL8jt5U07UWjlYil5NgcL4LpNPuN6eR5NVrFelljIiPra4vGDGySIO4U
ZW1zMtcM2ZGXh6CPGsj+j+CgkZ3cF+j+xkwoGiRGwsJi4pBYK6Y+eOdniTqdaCTl
w0FC/h76NwEB/4ztXrGYwZbfkvUWXBXh3RlKAtvevFCKvcbfhAIriC/QUdGiwR7M
h7U9GA7Oj0m5AyUt/JTjcwji2EZchfgTapxqZsLtxo4DTO95AOg+ECGulRnfsjAF
9qKAiE6OSoBqRmSpJXYn5z2udMBuBXT3ksIDihZ/GnH00BVI+oLvwiuOvUGlCqEY
iqJ63giykWcv9ZjE9AH1Z9iR7XESMKPe5NdP4LF/tHcSvBTHr/6vvPTXGaGxygdi
Xp9VhkCl1OfeHXT9VDLPTZSIq1IhUetjzSE/mHzfAuzHRXIv5iF/NTPOglU4IVZ4
oW8XRJ0sloTb3fNsdVofKd9BSXXLAImhd0rFDriJqjxwAy+z+FPf2vUbeUtzfs5h
L2eKHOnNYBOIyl7qWXTRZqfMkN38SAwZzHtu4V44Gq8sub6HPtYXvDc2OAIHJ2ME
WmG5HmbO6nDzHQw9CIQn3W68tLam/JhmCGSEeBAajOoZtbleFZgFAT41XdYn0ta1
itb1HHRLwIU14j4c2abGnCg/g3cgZk2QniKrbRU9EPjVKIkyCmYilLpM2EhVF7dE
Cgj8VJ7M4iIjFRpDD4Cthcz/jCSHFAh+EsYwrYYhec0VnHRTAirXjSDskqCdhAY6
OXiijp735tmTOQuJQP8SG2G/L723nlTQHYhSPAFTyeG6kKg1VOmEKwGcz/O81Vq4
PYQlg+S2EH3e5fLdExFe1f8GzJA4eH88a+i7mn5cXQyzXKhLsPYPnrMg+6bKCz/k
40Jt+Hxic7Ei2M79G2LW4bihbsMBeknW0roe3K8smpEaQu6ueW6/zE81taUb7bP9
cedlLjkJSAXOInWhhhV/6l3EZ+gHLz4osJiLWXhiOcK/fVLlo4fA2nD5OP6Eo5yZ
OHn9P2pipS6jsoyd2gPJBIM7SggzoP48AdDSA6luzrzxRII324US5le1w5XKyXZU
1ZllYauIAfFUufahLX8Zj3thPlChLoW4cN0pRYLDEpWf1362Qc1P0w7Rrjp4cheK
sGXpSXiWYBdQ5ic+ljLy8RMOBw/lX+rcM1uyKHtJizqSli77z7uJVvZnC8EzPcHn
RptQn/0Np8OvYRJys62WLeAKXs/uwac700EOydn8mI6W3UjpXv80Vx5Mr3nT86MO
8WqAPS4wkoix5LJtf7ssaOTmBEXXDJyvZh1lL+XSzWHJ7wR7HBKucePcYgDWF4iI
KGgbLRzaxsi68oHWcCbqrGqDZaTdo8ALAlmaYwCs7JIXhkpO8lHvYbkdex/OiGAv
N+osw8JUytmk6BXr4qXW7a72kUR3g9KOHwjV2EkhcyxvgH2nmHiUfYze33wldNNn
vhCmORH77j0UXWPwsu6X/T2wm8/WhVHPTdIskDQ2PzVW77MRNVcm+IKJhgiUqMsz
ZYjoyvuJkkWhyyvE13ocyfln3SihUIpFHfTrXOAswrlQKds0uBxdTvTixYJKrN/E
Md/+gk/hI6hT9oPs81CckbOkNRRFUJByF31CnWqpPaq4r6Jq8/Ifwn6UXKoUjHWO
YJd3luCT8YJ1buUT/XoqGs1s4MR7A+ORosE2CC5OjSjvbR+HM5mELaAIlVEns/mI
LP+QXW2TxfyajwUoO5jUL65XeRjPf1qhpsuhEZRvI49i7WUwA8quJrwkbj8Tr575
UAaaTeTQe9FvItAGFZ71Qz3VVJCFVRMK+TM+YU7jrdoS4/V/qfwq9aPn6VjC//ic
QiiVtpLgOlw8UsXD13276jGNMyQXqEc5vhDlFbfv5MkVuJqPPcs2pyxJLasCiueh
94jGB7iXpXdxbaPJLZpctRmmUnx0TelWXzlldcmqiiBz82a+TOCxJ+8FM/VtaAS4
XDgy1pct0JkovwpBGsX1I24PLmelsGEawCO3qNyN6UpjnsmqndMOivR33718FHFx
CA2GkQFFyMLnHnWztUe16Lcqbxw6dNgji0CmD7l7tOKRbI5jdJaBq/+DnWvESV++
Y0LIWA2aigcjom948RUAmfwpj9juSqb/60XJaQUSDbbjNRL2A0j7Jj6tIjfBHtg6
S8REPRZpWU6jhmI/zZ0baSTkrg6tG9HRGqlsBpwNgBYFy8rJQXXlMYz9bEZJT6oI
mCt9yEEXLRiQoGK9Avg8MAkOQPTnvq14vnRR2e4P/2nSFXV9wXfx045c5ReTWLle
eXgvD5NBMxERDe+yIJJYu2so63TxzThzdzaM6NVXhXtNJ5v9J+GW48I+7kR7arim
ZGoBj88fK8rTWYkitrrGmg1H5v9xr1jHeTfaIXXxyQOmVccU03Zb7hnS3TpGAkkY
WLcTAjWbwNg0zpRAM6hCpaz5GdOfCESaLC9Br0I8l8rxGkf2JxFCYTaS6eIu35kB
l9zxUr7f6JMUfuXFg3jE18SsDE2spcdiFEaYM6DYPK15quhq+aAS6VzmKnLWIGqW
bo11F1+ZZ8+BeywqnVQff11kWFOKmiwoN57VjxX4jOyO5XSTpM7mjGah4dHQraSx
GHN3sh3KS3uG8fwDhu+x4bEbLZAbxViWLoXCVrJVwqMhHzQg8PRuHoXdUMa3Ar+3
bCAw/W2GHIpfTHMsmQlfEDnmBXTg/XXWn55p+NccsG5gq09CkLe8tOQqGXBb5j6v
mrXbqLWpsEjunPncVNurM/aetBejFHdzldFhMQRAclzSPa7dIatMa0TSuHdUpe6N
4+QFeByenLkfae/bh3VdjcV3g1hsgZk24rznFRhaihROlYgXE8pnH11MRWEgXSo/
Bp1kmupT/31z3fVd0XYyRzc5D6p+b/zdgZonHfw6/pCbcw3OcauSOSCjrVkOljC+
Owax1FeRpTviomJeo0Lu0DP/dFdn0bkPduE2U+qBIwaY6Kh86tDiU/VEZseygYC9
3O2tFlhgpl2g2mB1ncETbrYXSyk+kogSExR6JNrpaEfbTl3IEnoDmwwuhau0ekkx
cABWEZ0xaAvTjxzlZE0jlQWZG0WdLZ3+02fU2REd8AIbo4ahs3Nh40C1VoChMIjq
lZwJ87EQDJw6Y0LoohF1YMdbOcGxROZwnqFpDB50it4F7ezON7WQXqYaCp59IPow
aYIhXhzGL+FzyHcCTo9yArGnXYluTjuPAAbQcNv1X564xk8R56GxblDlrjcbat4S
qowOQOwmqE9t2g72wVM1JRwt0kBK5BiAP/B9zmXNgy+O10ypytyyr4U9so2k+0Tn
BseTWECSVFRmbzbSs3xMTRCM12mkXJlOYVuTEWBKYCcrqQYmkcTVW490UmzXP3PG
jzBK3RNp/NpbsXc+SFJY/v74FQcauemrJt3vTE/D6gr6F3RHiGYSJN24P3h4rNIK
KNnqkwgwa3Tcg+L6AybHZfkYNNLKI9BrNTHNk/2XuVQKLNCe/y00YkalnXZ8LANb
PsqM+/0PVoQIhigSpPRo34wGFldZu5e4/Hy6GgxrCgK8AIroCFsEad3FEf6/0FNE
ufOe48KxQ/Q/4b0nKUzGiwmJj4Q3va00cfdIrPCrB023jWkaNrME7teNdAIyjmmx
JOoXSPcmHV4qcgWe4ibi+BT4h1YfDFCKIay0WUjEPByKbWPm1qjjt8nyQVKqYvzm
DudH3omtl/nO7GdsbHl47i+mXLPGlON98L4n8mEcExMh9EL4/85gyZ/Y/7Ey+WcJ
HSeg66G6gwfgqNw8ZoG5kZAtH40CDaIT/YxfRCrEt860kAZn86ydIto6R1ouL/Ee
2W8ENqlCqKEgmq//UzgnL2HWp0KBfmSWYygWgbpLWICjQHn+F/SB8tBpIvU1Kr0k
NvQfTVJgWBt4/4X5fIzf8UoR6JhDpulnyDdcn8agCIWNO+Fm8nN5tNqPkTG1Nk/R
4xU7hE50J9W7RF3+bOc9UEiB1M0WvK70TKtJAUDIp2vpspiu2NNrQDMe/E4ekgFw
y+ybNEyJAcGvw5P+xR1xIgEUuR/wVIUHU6H8oC6j3WCDo5JdBEL7OqAHIc27Qkem
7TDNrP+cVpReYH4yadIRESa2LLOPlglBzZgkYRDZ3b76LdIhJIB4MgsKXu6OqZmP
XNtsugYNabzJhtVNk1IG5SWph4v8PMDHTGasuJ+4S4T3v4YG4/RMxC5On4ZrjZfE
hLGFHEMuLC0dLu4ahL5iq7idMXsLAthB8E/4wo2LjTyC8VEYIgCuZx/Zyi9ot76M
Pt8WGfDY73ALL+ssiuNlnTPAzv8UboQvPqK2lcIftms6wGInT0y+LMa91dgx4ymR
TVqB40s1qjD0mh3n0rva7EPbBDwXRbl4/oYrinaPVu7HcPVLUXjflYgrP1mYxfMQ
qI4EMys6MTnogdez5KrsI8Dp6Y8VBCQmU9Y7FKUDyY573dHwZiA1QepGCO58VjR8
LqfAOFcK4plvzPGRfWut3KX7K/9GlShLjcd49fFvmmHSuyBNlc6P92vWj6WrdPVp
RdBjp1A6SP6+KPHuzMP0W49zYMIJF3sqhQtVbGWQq3Sq8AES0G6YwGADYNQ6tT6/
QbCi2ZTKF+B2QxIzI618BZje8bR9B1VugaHLFbJIw1evYABRr5ZIMkhjRR+CopP2
MTQf/hUX/s/4r8u1+897tMRdMABxdxaEKTyRPsTGJ25TLY5Fh//n59ZJ6x7hD2Yd
bBKS06IJM611t4i0b4p/x3Sd6r5reWSz0QUz7x3BuCRqGex68O3OFrDSNjsASKJo
OKYwovlkMjDArgi3NbJ6jkLvH4M/RjNqVX8OQ4JVPBvvfYQq0FUGa6Nt6MewYVgs
2lASo60TEzYphPohhbpDi6jhFuSDm5jV566TYreSO1x05ne+8pb13gApDQhz2hVQ
BXFVv7Ms+Kz5TLgy5KrVgs12CQ7l+KYy2Oqf08d2Doi1EKogfet7lQCYKLg4w66z
lZ5qq411kRUWBRJOgLNzZCxx6JZzLREpTqN4D88sa+oUPghvRK8swnay+xUCshDa
IuO40n2s9DQ1KCA+BJYbP+hnvAKVQ2aRWqopcv/oUpR/9+0yFQ9/p9tsnk/Q0w71
89pwrto5QqSZrU61KOTdJSHzVw/Yusolp6uCs0xpG1zFjXQ5ZTgbU0nM6/Y0cu93
6vTdlwR1D1+/NhrTztX+fTJB2p7MLq7vGHqHHbeNoh2L0lOCU5YmBz4DejRIb8Xi
RAIKtXu553vo9hHm+I94DIoD/aKFGGUsUXH0POAuNneOq09B61BPWok95hGZeP6i
quOnUp2F4Gw/M6kj/vc7SKhvv/yojLPq4HkFRcwleQahGh4ZTHCbB4/onWY1EguN
cDb23to/79QUs84NmxYhqSFxkPLokagN0QFm/RzYbHg4Ah4kPbJ61JlDDulSh75R
CyykuToo4zPAAyD/h0txosVutlbNn26cpk3Mfc9OTHVtEJGD5D8PXAQ/TKAAHZWi
wDuRvD/QQcBx4QdI6v9V+0A1NILo4CDPDuNMZQH4DOOKsNKAKoMTys6kQF1jv78K
o43wQNB+hgF10NVQME3zobtqWCnwZYFXYT8TMac8ZEJvIAPty53f0yW3NZXPY0+o
F9Kdc98akwxs9CqrxI677CU+n412TgnV7zTDuDHY/uPNCMcxtlTuBhgiebNZuRZt
f7KbuHyzFu9WVWKJBUwgL8inFF6we6TWoN++EjurZIaRGlp7Du9hoRbJE1VRaJLO
DmIo2REuF3ULtVCvzcchL2XmcUkoqEISZJi+dkFd6kzX877s3pw7Qle8Ln6PRXfr
vizH8sfjGmtYSSuO3HPbtZvQNngN/5ed746dZ0fptylIvV7U25XTVWWVKM8I45RY
3YeyKz8D7HM66ZGrLn+IGjl0D9wsDBwnBt2+fCrUUwj26BX3zgQMqteNFaXTNjJT
RtLRkk/C2+tjbYNQuBlpOukMJYyA5BhrL20aYpXE5DjCNnmhA31AHEy2GuGnv/hr
98AyGWpMXOvRyfAKSU/xlMXVHP8G9D0jMBoXprdk1SUvlp1OIc8dDbTvcfgL+I2u
wT+2eD9OFqpvbs1oc+OQr71ul6CIZg0c9d/IlsWG89wbrIk9e56K49xjv0iyZUEj
kE05hgD8DQwtCKrmkmmDb48pMyTdNnO5HX26GEBzRKoGgN5WVSnh0/wVw1RvHXL9
DKh5yJ4/o/9D0hjETY9lGHEYX7VWu38DQHnlxdEuYf6UtmLfbxeSl1tXQuW9AFNW
UhdVHGMSqM0okEU9Dznm0+rpjFRYu3obFllds2dwb98btFr5+PHf9A4d01Dtwy9i
HVHM0TDh92ixQmMLzY1VaaSFJ8bnMl7IiXNhveKTmDu/pmWuuyT4OXRW8YFldy85
pl9lWrfyKSxw6DEQIY9dBAm21KMMrU5ArnTH+pav3pHcFJFwo/se08AbaALlYT2Z
Q6+rU67yzGLOfqkEooppRY+Fqdu4rehtvIFwTNcFO2m2gD85vgX/3NjxZhzdD/NC
CNRlO7g/YYVjisIbhgD5ZPTOQ2tCOZmGIo/3+9ZDh14TzJ2L8xBAvPVmmrk8sgGG
JHQBS5I4pK4HWa54CoEKQGRARDjIVoMeZrag94yfhHef2+PTzxP7aVxsN3Vi7tBY
HJ+Fv/hjggy4bG+ZhJisfAK5MbSTMToai6Ax6ohGQKrbCw/JhUC0cVOOD0PKOWqG
8bdq0uUE6WVDG8f2xDq3u0P/JXouPm86ILvyUmjIAceNq+NM8DT7/N7pBIW3qfvG
RhT1tcIYX2B14sD7hXJTMnDRgDj6pJEvDQRZenD+w4Y18F/pI6MVsxJuUllWFsxc
yXJxNQHOP/vwbYp75UnUsZlFF3aN2NVdhtw8tQPvQ/Vs0d0ijN7emuBbixATDj7w
XF7rGJMok54RLg7EMmSZ0B2u1JgzPisJ8yDEXRXyNXhT24BCI3YVd+DeeACkeRD+
5Q9R/V9tlh0H93hUNED8zot26D4kVblaSMdbUlTdSfgvJUek1MFEj4xOUwmLmrk7
p8HyCTBIFcP5ZydMnG6rBoxEHzfKLMHFculT6IFeooefe7+mNrO6Pm5sUv9vIk3m
KysjOQ2BMIhfXM4atT650xmVifTVRWaPWA3vaHE2DzT9c4JQyxikOgYU47oeINkm
nOVkZXqpivm3qNgDI2stFSJUTW05Dmyy7sq2EpgmhWzfpnWmvtqejUII5y/arCUP
DF/9RxOUVPQ4HQGBpSDMS/8u3JpK4mtZR8hxAaXCe6iCDToxEW1jn66VUsppuIMU
iUmbKCzZH0XjEtao8iu8/o/FOM1OGWlbKusvCa/OehZe4AjGqN9SxkX+MLOxwZz9
7J7lgDfbZ/NPV+OnfnfnfMRAs8jqZfkkzkgf2viDOf0U7pJZ6BrCBxJzV5fwoWX6
Hn2/2a4Hr/5f5V746QboiCSvwSY/gmuhhw4ypj4wPvuox40x+4iBfIquC0dTd4tH
iGSkTNkM4sU6xrsiY7Kh7FTHmBjrxWgx1VVVQgMWUv+KukIOkIWutA5ZtGJZSSXC
JcSI2dtouoTtvXYmds6iGx/aXo8GqgGN3W5YiuinvCP1DdLKLhaghr8n1DTA5s+h
2qUxs0PKLhWzr55ShsNXG+fL0g1IuAnF276+VFlxKkdg5rh41PLNdM53QeOKp56C
1RF3zAdV+zuJ/lkAeCx1rS8E3n0QgTu/kLLYfKSCi86yolOsuHq38/1XqA0FE+vi
1/D756/eHCPC1BzBfsQD8Dqaz+budWRRPcfRCXrIIdr+64xdUvTxfcBjoJQcSTZc
pMH+DO9LHrXyRlAGH08kGpbdsDTvJTd7G9GvAlIw58KL9p+Gy90oc5lDVcjHj9ty
Uk/Y5YaGjv5pLEsKoDT2+afwxYXhpws1BA+dvUDq29PWDtwUQ5Rb+8KK2h4sAEgv
8UwJ32eZCLSIu9mTjh6M5IfvKh2AA2YY2z0m/myw7qRAzquwful4opTQdrnksiag
EB7XR4T5bxkh+aXcOIDKdPX8wcf868eg9fIZaM1uq5naqbHqjjFbIpQ9jsdT4YXh
mm3kLexbKexZnG73aFG4CPdTPqTWPLSoTitz7+Id0aNcyXS871SWF/bdHjkcY1d2
7LTkgUgu/a9dFr90w9ImG96TMNW05EdFp1IIU6XPUdEvZNrWr3qQctANyOaELVZo
Ieyj1d+/OBE/CMgLLUOL/8Ru8ebZ6BZisMjX/roh6kKq0AbGobe63Pbb2rrdVCfY
3V74Atm/2/PEwht4fE5v+V/ffCQD+2+wAlTWNGUetLxSHY9YsRFThvXW7kvaiWWc
TVnF5KzwarfhCom7KF28AzBEWQsgO52FHG3Uw8NTXCs/3/5EUw2bepu1cZ88NhoH
7VfYJ6MJ3172mu4hFVJ2jiBezqaiMvKPrftxdDzhchkWZj12FJxsJsscOXS0QkpN
wpnABS06R9nAx1yBoEXKuQH8S5cmIS3Se5urn4w1Fe23WRmVAaCI33pdIJ00NxwG
s5wLNzyoFpFUDnic1fuMRcEKjRVZSVViIDtgxWGdfEhd5bN5QENzW/n0UimSlUiJ
idV9sAAFn1ZVBG9Lo7hwKcByWDAZk+BNHCO1cv9K6LjPFlrxAr33jt9LTzmx9oBv
ssms9UOU44otb12TPCHDSDRiL7o2X4sHyPrcaAS82/wNWwKt9MwgMfaYWsYlJk2c
cm9ctY1Ii3q1beAWy960HBR7rpAWmSTDUZUT7A7s7NYy2mDYBvwCAEAdqKANYq9o
t71qAsXJcaqLkX7kBsYlVQStw1v7CZ2WOym8ffln9QleJOzSFAU9rH2GwdcE5YbR
U+YJXYaYIGAauawjVpZc12YovTcrcdzTj0w11/c/3YSUPSDRfQEHvYXlWioBPAct
Kk0y8X9qV8CjqxZ23UqK44ACho1X/Of1AEgv8eNAyu6HzXWSDIEZs5D5bc2lYC1y
WfQGq0Br8CJsaLGk9BatsGjTJ94Vcky9W7xURKxAdmIUogg612nrgeWVm9cMPNZv
O27e6Zwff3eh5cXyfd1LvGBxaUXnZWRKSi3tmis1utUYegUXizinLppwwu8w7Ti8
3mM3wZNO0GFdaV9o8JEzffUydbBPO5vmwmnMx7Fr4JBoFsslX5SU9u4+NPSOnkD0
sykmhJ2uPhljtBmSSuCqxPjU4TpY6ZZLLdE02U696MKLl9BTXu5TYNGri8uRrVJ1
9EcvrB1toOLHbVI1RchPtrG8iqNuMavl9Jahw2tunCjkwtOElPoLw90FxzY8QNxW
Ln9hJnRWw/bmwtCQJZABnD0mODez9dRrIosapusS/74Jj0+f8uKDUNvpGIu6Id4X
smCF8wA6hNWB8qqWnF5xksFjyrEAV5vdRcrff0INWGhFnRhWK62GzVne/zl7TnXp
o/Om5OlNdITUnnft9k506bu/pgRWVoGB604DibK6+mctVjxmodEukdqjDmkefHVb
8uU0wwv39MTqLOazQbS66sNucjTlfnbfABlMbUc4yjzqcUSwfKAkKB/RJTbHQjoR
w5rcHXtune+yGIxEMYvSZhPoftRPRZ3xnJgsG7TxaFMD6+yCA85PPIWR2Wu7nwBF
YRE8oAcri/9ijnTz23v9KEKmSo+EXmH8PE7oUAdLGEu8TB0s46H0wGWl786Kx+Tk
Q1/s3el24cDEGmMOVOulbfjWbGgI04jGXar0K20jgm0KsaB7Wwk8az5C+9FRvdiy
RwDBEfj2BFMYoAhAH8SW1mFeVApOA8yQxj4rnJEVaczB8Jlr6C4f/X+Ky81mp7B3
bgIHXIQX9qsxfy82cOzaboM1brmWhe8uY6BFfHE35iclKHBCjbF3ag3D+QQ7shQJ
ZQFRtna0E0nvyJSXZ9neRgkzyBiR0uLmgRzIQGrEX+0Tg7QMbP5SUXG9PSwGtayX
wrMCZ9hszohDr2iSxX/v0JsabUo0VEGRFKXGIQt7Z81IeMjireUZn6ouhEHDC3ok
R1Got8j2caR3ZiAQcpxBkFHI6MtYUku0yCWhBJ55YL1gNyDVUYur67YYkxyjIvR3
AOYPMx19E442JuwJ6h9UYkgQT1qkBJ+LdDLu7j60cKhAqc9cncMwfjaZmu47W6O3
EevmUo7jsxX2S9IX3VSkM+nq7kc6j9oX/OpRHeJvReQP9eow4v8OJiPuhNOFZyHY
Ho5MZ2yMx0B/3sVUirvqn5YTMziGTDKWapxXyZdwADnr7DmqJmwnPV0khsfbjyb4
ga1s9+350pbObkiMqe+feZp9SVke4i0tHDABY7un7Mp7PxDejuqXCrrhuLk8hcq3
mUE7mB2HTgMZbHwAALxQ37WnrM8Qsi4rvLGSzcmCwbwQuu3ILq6nJNQscp96sEl3
+csw+ukxNMwgDwgLLAan0b96DYb3+fo/CsQ6/wxsvF3uGNSk6HkxuWbXsY4Kb9vD
QbB7VjX0QPGNJZ/oZG/0m8W2qVw9F4UNcFeC5P6Hm5CPJj+dULQakILVb7kDKY9p
Gmo5D/9EvmCHEqTT9f2M3CKCl3b1iPMDgUsywyfpGg6kjAYdI8CmuTCu16vNUzOp
LGNsBq1RTiFk1Fh/z/H/LeWh8sY/KXLWWtA9fa+RTM3l8vh0CQL0RVZDmXfY6ZRy
v9i1wz1k5/6cXeYWCcUNlVraoDiVk+o9mT729FJ7qgMoc8N1f9pZfImNRiSW6NMH
p1ciDeDFnpDLjRoOBkKmH5xccsNgzmF2mQ4uexyJO5RZ5GVezvTwDT/qX7qMdJrP
BHltUuKBCmIP2mb+04oZMMxzSTkYXpnBJOA6g6LdsFchNIS7L4xFmxhhOijBhu16
IhIultTVGjMzNuhcuor/jTesAt3mP8VNkr4N9s064488fbM09g9iAPdlXjX7j7tF
wf543PTQd/AoPozr/sxRhesQ8xGbYzF5Kc9GMNyVVIzFA96P+tfFkgVziWSOkxOv
08qqQMWVui7bbRw7uRKcGEHz1jZwZaN9q84cRhe8f89Zwgo8LNSqe8uOurmB1gQa
ULEAotSyaKAZ4Z8FDZmBryfcab6lPCG+kPksWH9ulk5EmsRc/HnLzy1Kzka+ggKx
D5h/Yrjiz8La5Rl1Yh5Vs0YNKYXJ5o05nJeESevik8hGRW6Sax5AWhaOCs2N0IqZ
L2whRavaudghVzsFxF/RxII+yru9K3Doy+e7iV/8vSKAKimFvev5VzlMIb/mfCvm
JphIzGzfxOePH4UsE+dhbBVitUMloeHNXr+evHB4KsQ9sURzHvJF5j9rDbn5aQGv
5juvm5m+CEdSLB/yggM6HgqfuXr6U+ON33A/GJusqgN0qZ/x3KW0zuTKnvEP053F
mhi9BL8q5YImv8RdIDgSF5AsGoUyx7FvoZbxEe0YPcjbW/wqWH/rBlGJfaHkHBCF
3VCYKjKl21Qw2vFPzgU2lkS2DFDA3W8DlsdCOSFM2LVKH5ST3wks1yfwV4w1fyYe
J2tl59SkpVjdYxJWPta/2vhkVK2BEcKJuwiY/2CfS/GxrysULckVANyWoltvxXx2
h5GMW4z48nE+a9moaJcCUln0Agjr273mwLkLKAaSi/R6P8VAI/va0YLhD5/IolJF
uFLbE5bUNJfmhs1rehJpqKvAh+0i66Vczdy+6wt1eZZTTRcfzWY+ZpsapAOgYx4f
ywt4bzFNdNFveiRELuk+cnnPIlldLaM9rZLam5gXktBeQV+DXBPdnAkKwTRTw7bH
SctDYTuaEjOHqARhK+d/Nj0zc5CWAIjUPN747/C9Zb9MCPIm2rG03rMDlKKPhGy4
nnQBeLDDBwT1qmf8KuSGQpRsL20a8m9pC2Me1TBIj0H07LmwJYj7YOcxW6zYFxyu
e5BYH8KUPUlzWcIu1j3cbJz50zSZYQBxgkUVB4D446ir/7HLoYd6wDmX1qNwDG+S
YR113bZnEH0BU2s7o5+jih1DNHa7Jl2EE98g4u9HiV2s4pRI/BSW0N3ujy5KSvwH
IDC/UqsdmT4fdAsGzCXWMi1z2nhnrInBtVqZKQh8DYyOS/qNGYxxsivmyq8lh/lj
4GcqmcJJJ3GLh5vNFagg0PI5xQBTWD1p4VB2eSXa0NtG+7YN09Sp4fJjqnhqrQJZ
7P5OXqPLxlHxeDJv9sj0aotnA//8ZxV79+jvsViHJi0hEl/Ams9Zr9nNlC2smMC1
8qXoYM2mQwPdRCqaoJhrOfyEGxClvX7WiXeIGXObqeUBtf5V+sOZVxoyPUQH1yxd
EWGxkYr9GC89JEKw/0T0pg6uSeZgtlNBvEqDs7WbajtRdpiu7Nql+hfwBArgceHH
BA5ylM4V6p7pouJZ5zUVpfPxTSl/P1/7P+lUaCWs3sNVzD2G90WoydM2wDlackD7
EInXMdO9k+FgTtac2RAQ3hKhl1DwJFtFvTPwW59usDHURP38LAEYeKco+ADvzSj7
e3/RYswv8C+22VQoU0VBRWAGNzIudsl7yZ1LvHn/w+3slQQ9oU7dfxD4IZ4G/A8h
j8ZogZcPf8irT7NWfmII4vxcWRPIKzzz+mk4sUyhYdW/2dItIUdn3ldqdSBfjs3+
i2M5JUFqzGYsIYj5OWsiKBZiz2yRkEIJILnMTuddkuoNs1za05jEr/z65s7ramce
3nCsCazLNHCvU9Fz3i9GkDY9J96m2r1BnDQ7qLsaFvWgfK8tThZJXBmhCAwoExiE
r0U/u81alGe/j5TLhak1mZaPufsFTCc60WuLQbvcUmf6Xy1DyoVOxRRud0a+cvvw
eoXyNCql2fDb6Cs9GiWh70IoXN5w0Px/3lF82sQU08nZ6r8f+rlrr3AtIQg3ktnH
lxgYuFdQCtmoYnszRwo3bX98fKJlQnKB9s0IFzrVqqSLBPA2n5vTJOoInEV1l0Gz
HcZsg1+0UCO+PaTVrVMjePRUKZxcSprcFGkOYcbZleduKZxR4429/NvpsNtB811H
A7dES3HbziuN9MOwsL1XNDPTNmlfihtWolfDkU4dDknMMnFWDwWWZl16a1Gy4neT
vmK6I1PQyy2JWoa+9FfVPV+nKLVhjAKHH9lO27mmFcmnjUl/AFEc29If7EVsX1zl
uzTbJAP7hl6q5RK3lvQ0CesS1Vk4eQF9nEkCSftee7+4+/CsQnEhTw7MeYNe9fEe
cua5EjoV48OblBCgaQ2Y/zPrOMY4iakBL3iFXKr08e+EhMTRr/dhpn7I9A+s0Kd2
vEKrP+NYyzssry0lW3HEVdScVtSbPGsortYtS8m+9gy6EWiWIcfgjmr5Pa2hdyRY
5lK9znoQ19NpLB1tzPH7YoNkdEPuAocjvGo9suCSsfPosy8KsUxKiY4kQg6aKML8
7AX+Xj2S5CSTAJxAUTv++e/TgqA8F/yxanGlfzsH7R/qxjzezI8QCgyRBaNqdUas
D1Z1O9yVo/VFKlI0GHpdi+vII7PHB0r+M3UNyh+GFNoHX5/AecGfX2TVLAFWWcNs
d0mllRtOIOOFAAFlavmMHfwvNomMR+G1WP+x3Zdv/33HftU15qqlbGyN8TkE61nT
ZuDcX9BslXiTNARiK2zUK5KtWivy07NZ90KccZdGLhB1b/W9Z3ns2xNer8C7uCzu
XUEsfVX/lT9gCLvhaSQJfnberVVQNc+3POUTScrqSDnrmjC8exRCNfSM8mPLfsZ8
9om28cammSNFxbYlwhmMNxE0RQSvdf4ATCU9P8IPDVfe9G4Gs4O1ZjM9sPIa/sMo
5UUOFCs2pL1wKcaO/78lkB5hL3tB43RNsk+aHr/6CtBzBVBZYzlcX6WqAFQZqQpH
98lFeciXEeu2l0czmt1ea58UleMQnTpr6OlrbXwo4ci+kziZpaI5SOVVxdZHKQtj
g5rT3SNUFEcEe9pKdy8WBpSI+oy1zCShvytmXHtxPiwoypVeyOBUvAFNKYrqDoC/
6a5MXTiwM4WChe3++X5eiRoKc2foEAwJ3STzEkPlX9YvG52dB3Uzb5gsgRh28GyL
n83lRip83lcxW3RtT4kQPRqC8kZqCUFI5xFdX94IssunzLCOxYj+jxUCnbOADEj8
TX3MNBSfSMPaMN5MuYA9JI3MaPF8ygiShMM1IHpie5gQ1Kn5b32EyoP9U81tDspF
HZRM99mGxuHW7wJ62QlWyc+FiGIPjg3EPc8t4mR4Q1YXNSgiR9fRnnfEAFho9qrf
H6ObfA6MRLHEhMXlKA/5Ni2pkaXYk2Jo1RpUFntTYe7IOFVFR1jr+DhzgqCZ9djW
6l22/YaMyyzVdTXrivFohmfVr+xBBwQ4b6sPLCTQxktPREEg+d7CVv4PSxEuWKM4
2wr9FgB6m8Duw9dCsxO9vD5UjyQb8H546vGPyB09ccybJwdkf/vT95e1XpRm2YEz
I3P5ilNv/cqB7ipSAJISRAclmXWfByvaLnsRMwttNfeM3oHxT6sbwlij8z0a/yW0
qW/rgWOYoQUPvaggAxrkRDzjIBrMvBJHYsnCK91elI2F7ekpmmfk2t2ZslZX/rY1
lQruIzjJdIYoxF2zk/2TSqDxATUQScUlK15dHk4zGM+7Z5P28e9O5yU9swGtLmBd
JvMKEBLpdzCTcA51deG1zg6z5A82oqcN5xXYYFXasVtkJ3OqxGhnVWp+Xuf5L9oA
2jP6BxE0eQdQOJ9TeUkFB2NAf4esVtkKpjbO8BrAqicMFZdFtnZfeNzmzAtnAhRZ
5rhywli80gTwbQALMNKf00eC4alnGoVhtx0YMxsCUwQe27FJU0KCb6cAUscRiT2E
EMxMDXf0KzCYa4HBEhqP7Gt1Ttp5uZGc7vlVbeG+KpqaWUikXqgE9dA79iNO4p+2
V39AKyBZDWHyUKq55phYEV68hpdIvlngkZ4WcsKxO79Awl3D0stZJZd31Ll5shxj
YEgdL23iGVIVSE0pXHJ8uxxcbYQ0n7rmR2LNtVOUnhR/IphImypXo+metc1k9Os7
A6dkH0+3ewZ5jkwSwOY5pHE3CqFtEZdwMoUlB6cS+Tr8q8D7KmRrT61xcGlmynZk
J/bzlVKaSrRFerLkR6Ayxl4n4v9Vm53b2RynG/5RpXqlrbaeZLYb/WQrXidJKdjC
O1Fs/UXcS18NUmCLkIJgRqMpxDrMcUuBZJdWI8CIB2KhbnOsJt6Sc7sMrrrRm7eU
BFopgwoW8jEQSIiNBDZCsPgNd2MHwJFN9p9cMzDS+qOdfhwaWB1unllthRYUEXpP
EROG3+xNS7VrqbedjGFD4knrvFZgZ/gbWkocdsJ3+PQ9Bn5+kLQILD9jwZUvqAL2
8aYqzqnTY8qaPBqGKBRtKWVL7s4bn4VLYTBiT5aC+q7PBzgy3I8pL+ANpCAo3b/4
z4OtdTAKZ3j3pFjsv9QdyjGka9bd4krim0lj9+AGLI7sNAExWUC28JKam8iqaVnK
IrkFFm6sNkIzbQvMLnaGiPhT3O5fLpdwsyw0ZQnH8ZcLAZZrOZQvL1ECPqDcAecJ
i5+ZZ454+QemOhUYKU06bpsvDMmI9aN9ixEk/+FPjukBvoLzz3o3p0VN59BPytVn
Xr3dc5JidA7/RKjUCVrsxM3oSY2ZIpFfYhOTqQ0jPckRQu+4PlQWW8HKtB42hmKJ
6dzBi8iaxSaNQVOjH8/6NqnXIBBhUP63vnlKSigrbaZa84ixxXuX2SJEXENLEhDN
ut9qD8icCgWFQbACu3+uTOZtHnXxdoCMdxySxkdYSfXqKshc9UPtK5sr4UMTh5x+
1X/G97nR5o1muYFuoyD2fSSg3MbIluBsfSEmKXBsYaiU6j+uWCA6CGwxukIhEdty
6fEjjb/6rkMQf92J87vH+0AtB7CWpcNLXrrbmdWciq8JRaGgn6xS/gx2WHqn0PAQ
Bzx8g53bNlHny327PkO7kuo+E/Ia001Yp+6xpPqEKMiyllfysh+IZJof0IliApZJ
iXTD46gPwCIBoUml1/snd5K5D11S9pTXxcbWgf5LiYni7Hnwmks9dR6p8ODJYkbq
X4RXznxK0X/LkrifWZtGYLNjupj3Pvq5Mi5T8PmHS7s1EgcbtWtMckOgSgHneoGK
7/9Kq/ba3tfsgMTMZXsXatR49R79NfW9C9k8MOmaE3oH+u0Yjmz0ZZU0QBEi2Glt
1g7gbPaH7CxA/8huPbo6euaUrb/XoFC0TqSmLnomo6UpImxbp4pKdXiIHxib1Ao9
FHuqNEOOqUFvBm43rANaPREEp0gPAxBQUP+31KPATxzUuodL2kVgwjglSlHKWNgF
bSU5vInqdMXuEx789Kjps3bt8t3hWXhMwnQa7+oPzoam0URd6SfMzuEhuWDKaHr3
9JyHHDHH/ZcAXNqem3sL5QARVGSEbVNEJPYTUZsjigk+ABW/f1Iul3WVERaTtxA7
kg3bjEertNuwUWJHfofFbJ/N7hnvmc+wRNXV+w3Y5Eq8Akbo9Xgbex4n06HlaC6g
0sw2SXuwWSx7IIZCpBN3khgDq551WS5Tv8U7ktsX/lxEsTUN+aD77FYmvI2eVE17
25+MPx6ANwr0/ZW+2y3794hwfnxoCyzW4uuC81vXBTnyxXQZ9KBiRLW/rue3ssN7
8lF6mLT1ZMHX86bxqTuRidKG/4TtvwJrxJJ5RikJBC5gEznnQ9C51TJyLTbr/+tS
dfrWDLTlxHBFxcd3cpYT++Yv/TMoRUHTv3FZfG74NkD1rLqbp/ysGlIuSMLHI4V5
bkhPgqhzOqg3egkf/n25LxF8gKZEKlKnvpO4rfjbptqIV12zO5yPvJmeDiQbZvJb
IYYYRNEKqklcC+mm8np9eR+nQ/FXfufVDW2BsDC6IdSnOXU/M99K1dJtke2slJaJ
YxwbD6txb+hIqKh8M2mnPV/FbUnKoiIQxveYydNSqhsUcq+bZfshtMRz/3zd2fXz
ybVTUsSEFwd+wDeWc1Bf7Z3Vk0BFRHXrJ9eqdiEOL9VlXkGnnoQFlxJny++jkXXg
regS/Yk904ydrKEa2YWI66N1geG71u+DsrKHck27iSgn/JFgYSlr3c47XHM6c3D4
NG71Jm112pJMNCR1Xg1Y41p4TsMADwf5jwIgMLm8dXu9NFsjpXpqag2AAidY9HJD
t+QsDTRQnTvmgolH/V6RBKDVSD75xWjBTIxEDAt/+DpNRgWE1y7XQwae53lMQSmU
PBwLf0XZrIlgTrh3Uf7vW/3WbU/qu0K2oAGXRvCAcIXLbILyPXQfT+JlIR/wikfC
eBf+bni+f1kbkQWuDMlgVwgD22DmyEQdEKGiKvpJXrOZV9l/avea1S17ec5m2FaF
AWjRIaljfgVM8sfjVciPm78VBdP35Uf9Q5DzJNYa7SRZ1m0OkMz/sfVSlmOEfriA
adAEf9Olfq2rRGceaXh8fgXz3/2MxxwJfXdTdAGRL6cO/0TJe/KUIcQPwulJ3mWg
iLep5H4kl2yoogtYjdRAlG88FmyiypRnO5qyn7gKDyRZ74B28FEmJFmdAzGxaWJ3
E93Fgaj3ZBes1za3E8QNlhBOeKAaopphyHWt7xK1xyrnRm57BzVVSQp0EhyX1Kc3
Tyv+4zdcgmOtMb5umZqctBrcqf/coCsDLz3/U1mVRVonxEcGU+Hx4hZHwAjtqs1J
/cYeRaapP0y0FS5M0hy2bZiCHRWGJq9FNcZqM6/8D6l+vRGhGsq8xytAawMPba6f
9kXyIBJ5R1HtGb0ZV19YWUCb9JBc9ys7I3/0lfq7jvAB/HUYWZZ0iGkK11Pfd0kM
GeaOUW8gDV1nsp/wfGW/+Rw87gtFn+BQavpYP1vzDdEs2L13yKKcZ9vYM1fnNRgP
OIG/qns8iNH8zjNP+gXwEyr3AXl7UNI3m0Jwtpm42FLCcV2nmypnUE3jHnTL9j7i
Il43j9AtufyI4tSNozTECmCLBy68U49YGqGYoTP0zkStC/NmZA+moUMssZl51R2E
8goX5ehLJeIKMpEQaWyiBOqevDvZshrrrf7QbudipEq72WgtKm+dzqGR1CBVc1a8
1SCzPxvDA41ti12NzxMU/+wpglSGZDxpWjWhdSndrNa5HPPPu6dXwxPkSXWIXPDK
rCy11NmVzFd1kPQ/Pn3ldzMy35iuqcKIoVW0k7V57VcmISCxAo2PgWlpsE0WuKdS
ID9zsyD4hYO33MKpHQFSdbFkxQVShMPWzs/959e8VYctyzI4ER9B/RorJ3Zi9uyW
tOawLgL662VJvfEiTDRWPlJ9xmQ4M0Tr44nz/449Bz04mQdHzaDn6QO4N8RhDZNV
zMfV4vhQhq6NsYaD83t7Ww6SDfvu10I3QPaqlSA6Lg0/lbh4ppp1vC2VWaEzgpj4
+xx7G/aMSB69OQkC5i/pKG5Ufk+gADf/H++8KV+MhWVO1ghA8Gs1vPCy/aGb655k
NjC9LuHIsS9XEqwhzaxPbG6mszYc2mI45ITrFagPv099bWrbI9vxuSzlAEkTdhtB
hnGKShHJ/4RJSpGcE4S6vp6t/MtJwEQQ5t+bUJNmuNRdpw88++BwhK0vDJrQXfN0
zmHKFTMT34nGsBzvym09k+0CVA6YKQ1MRpbNI/5kJe3XVEv0JjcrUOCg6sJwiUx1
l6lA0M0vIvhuUu80egSvH+q1vXFWi5XW9I+h55cSqSoQwqePOE1ptz96XKGkDBHS
8j7OgIa+eP5Yao40wDvHmA0N4uIdfMnrksiqGeMnrGkZ46MLXUB53I1vwcERICfl
fI3bHMKd5VmmFfdpJ6dSxjJ1KDnWnholfGcIk1JLNA19dEzkoAmaLMFpDwFdkADr
aKwJTPZKUWINhp7hM9c4ooqvDDi4AUK2rdclony/rQpCwR2Sr1DKxENf9QvrZZ7e
pXvCxQcBfHZv5mGd1DVmqcsPLkJr0QUV+vpVjgbVP76e2T5+M0I4Si5MGeD80nUp
In8r9YQEq9bDIbPiJoJHwWAKW0EQwSaLElGOBnWUhIXC1Qne+bI2kQW3mKpSaROV
QpHkTjeA3bcaWcA1IuhH6aBfEdZqwJfPbrTinmerqTmjGt/IajLlH+zIXliC8cLb
vbhuBTSgkFkqxZ+Cp6M76SBktlKJBXiFeS4LB8jNiEbwMfA4sI2x0jEwIeEBZ03m
Q5vkxc8UwZZtlU7NoKPDV1vdxjRvsVKiq9wclE4CGpEgB9oB8844VGHzjgB3ywNX
0sw0R5OvwwYxSR7kRXkmEP+SUtXoGtlGk0ULS53pJ5d08PCpNmFq5HoNy8IUgJEm
DBh03q5K3FkPqMkJomTU+BsRmAyarfCl8FUmAI/6xccr5TOIYqJ3vWX6oGZ46ib3
Q7NAxfF2B3zKCgH6LocNQNhcCqTAH9+d04JMPxKSIeKmmSLSC18MPWXUHJfEqHf+
pRtxb01WynIfv52V3AHbkAM5/aG/nB7mbznCWWE+qmdlIihnosGeRU5EJZ9Zf4YS
gw3ERQodnd5pSsPAZUL79AZdSEYeZ0UtBMxsa2TqjVpZ4e4X5PhozpVD/1wc+qYC
5UM94WMnAcOltl79rIBUevnGVGvkVjm3FJwggCoXUADZ8LdavNb0BGuWzoLLYeOo
Q99a00nRQGUcWR5v9o/hw99+4hUO2jKuWg9c5SbskRqGx6Va0Rhf2lYS1VhGnm9i
KX90kMzDc0+iMQOUa5FYzC5RVUd8D23MX1ux6tiq/7DW4R6vGG0afjcIHC108p7+
NhWnGh6mNyJYKSQE49VZ8yPQ4RKnvtm/n5V4olDiMyDKK7x5UeBnaJOPA5gqQE5c
jK3HqtanSGvMdeBrgK85VlDGX2MUsXxq822CzALmhNd1r0bmhiOBsiT5g6tP1N6d
uK2kWz5Fi9obc1/ok8c7muGOAhIUGuu6ISxGDUOcrjXBz6pydBHDz0PDpGl5DhyF
8/6NmN5Jv+lmxLvKXIpKka4Izgh4ZsF5N0e2FcxFDR54Iw+xjPoj2Wjx213DffvS
uLvGVxWwH1M0wMm9y4d1af1LrAXImcsYCailUede/+SJoVYJLYz1axV7gzWxqPOu
AYdclQMajNSF8UCf28lvfmbW6qhnA1EmYZIh1x1DtWngYZSd/eenE4StWu7GtZeO
YBGsnarPxsHHhqXHvfEHB4OnDunxFOOUmrGnBnXwffHS7WyetJZ9pV11Qm/TZLak
5+i1+XTcpg0qQPVEh/3jokab+yFW+mpFvUs+REP7Trk9sgWJoqeNjvTHHVIPGRaU
A830EAuUNbKH4/1x+RztMmNLnGmffWNNWxMxxQGyKAz1nNQ1fBxSq0sRqejlUvfr
rY/9AHg7yVYzX4r8lw1aMKbDZzT1WITrUYmdI6K+CbWm9GaUp4/vrEGU6M57Supt
d6Zdjdox0mQj4+UaF8B2RDNR/+FhWepYVkw9PutTEXG/3A10UCXjFQmmULEic5xG
ClmJaJdrlf5gRUSua1SJ/kUtKpKjYGnlpT27b27HWYRaoUAM+OuiO5Uszm6R1MjC
4sQZwri5RDMUQWja07qe9XPDqQl4AD8RJIt681OTyIDOmf3LDqwFIq5P37T+aLoC
sIj2j/OOxaCci4bc34CMgo6O8w1RRqf81BRtUU94ha1V1ncaNkXHRYQqoDz4GW5W
RDCcOUXuAMS+c+J14xClT6R3ueeOtQEAciko8Q3QYZBQxFyAhDAfbkKRv2o7SC+6
o40D3pANKJR/TpjLGuxNlIW67qYgdv0kn/0/ViEYJ9OBD3UsvsuXTuJOeTvd5+b2
myZKcfy2j354w75O/Dy9DND8jk7G1oa9Z+m2oFgZ58rGpBB++jEhULjDFy9ymCxI
wzGf/Y4EJ+m6coC9XQL3dTb8ppt1Zi3Y30G3VUPYgU5GPThEiCKjmsKeLNvw0VIi
m37+zpt/i2PJie92t3+IfyObNP95o5iM1i0HK+mJ14cSbRsH1oOyh0QAW2J2FpTD
FzPlA++22BJYERWKkRDy/b4VYyeK+FlDsj9g0ooBgYXsgVBjjqDiETkKPpb79xYa
gYHxtp55z7VTMC/ffYtrnojF6xGWhjPxu2eAX8rTPDkK9ncnInJGk0EbQmweNAmY
Q/4Hbr9BGtEX9nI72NrVZhx4g50tVc2v9WFQv5KWUjoczDpYTN4INz7PE/wRpT7E
fOLjTsU/P0WWoPHg/mYbygewkp59Kp16gfXyRN/dT8EhcEV42g98ECMOyX6//RjD
Fwgo0ALDJc7c8SwnqHhbJCim5/eDe93EtyE26FIwX9MFA60+nrDCCiFX/lEOEB5W
CUcMjvRWHiRz6nO4R7XQgZWdgCF0St18uVKNvPB0h12+5zg3lZ0M+zaSun6uPdaS
xQNORQmQkzR1+kNnvIIl+EZkR0NKeTNawP7rEIUndf/YsDIjYhK2yjYIRwQtm6ul
fwfT7UlV7vJQC0Y+WeAh1sStzVDW2ylXwr2dlvBYmM/XuVLE424cTHUYqtuJp9p6
MUbi3iKLwAAID1g8PA13bwoUPrYX/RwgJIhdo9JdSEru0mQsL/vQnLlnoB+DOIxh
9bNFgvjBWxw85OksZnTYcz90RA3S5/3TUj6GC2XmM7SnLNDq+LK4pxOQuWgdO+DH
+4MczgrPRsREHb08qebX9FVBovg8Vnx+iShHquGvD23mqL3pPu0Egbl1xpFTcJ3O
Y8EpFKNg6Lw3NoYCsELDuJrUgT3HBegkxRYDcocKm4PA71bZN9L+Jhqdkiilc43l
Rl8vnbeU6H88pQjO3IU0hnYcNhBdhdnawynsJ3FgZD2rABPA0TiV5SXoUL27OpPv
rIBQyR6WetK/Z15Qvyj0TtY4+Lz2gecIrBAC2v+0/pjD5hovBsvB8MiS8SGZSGjX
LIQsXc9XILsOs1/iT/SL5Invf9VZcb2jRcaqKOt5JUU7gkRyC6leTu59grcTPdWI
5MxRZFG0KikLuLSjtHuHulquRpUOFq7EIB2oaeip2JZbrcea7Moeuyrf8gIJ8js2
Dux3x2NTGwhzeOP4DMyznC8meY8R2zGyA3YdUve4+fygeEVQaqfBpOeSglFN7TCR
N4cKWFBqzSlTsH4amjQM8Nn8ivfM16RVJlpHgvyhJCft37/uNmJy+Nu6eCW/L94t
qrJMX2c36/ClxIXW4C+3CpAzN+CKcMo3L81cSgXeel3fSRENMZGkeTCCloU6/5dE
ltJfxFIjn+nnUtIk6ZMfoYpPANhjX+JvyhiVXJyuIr5omV78n5yCfIBS9BxFxY9U
HxB96UIvxWMmaAzOYIxflnvtzrX7Z0xYOn/W8eTByPCQLrxG0TU70BkXE19earI/
vVJXDzROI/XfqlX8HS7a48kpPel/iX72oyVJYztWmjC+ZXZBfkbiXrrNqini3NKY
WqENOCxX5jsL2nTpZxvZTwD59W1btLzoOi1Yg0mHXNGrKFYA6l5i90wZBc6J+1mW
43kAfuvA6VeaP2wgHeL9uRp36df6Gn/nsAnV+aRORyy9D8zPT5JM8ZKcRPygU0MH
7Oogx7qHGrxIosON7/JlogN4FhZsFMvLaYXDnOKxTpjsu0ZKYs/TMXoBS0IQeK2m
1F07J6fCs2wrL/sqC4l3xKJWUpiIk8s9W2BQGGHIwex4lZTbxDOFPiql93fhsr58
SwkrPOWOt6RMlIrK5P5BP/lY8Lr91viTn+vr4HVs/9KDJrUn00yuqLcDXVGUAO5y
o34JXguRQ3H3FMIWQELmeQbx3umXUAiQ8d6tHxO4vd4aXFmGtwGh9Qxzw56+/0iu
F9pKPBBA/+JL/d8SNUU06XVT973ZKKSLiGkFNnuph6BBG2lCZ/ckgh5K5Xzhg5MT
XeODKGu46fBWxLAQJvLBBqmdgCWqU6P0bA2Xpd+V+kyF1kKaNNlKVi88kkumVHdR
WNiCHxMXh78Gh3ZgCBn0pT4tTc5YiHxbka9rbLvBIFPoxfb4JRJfMucDBl4utUEu
4eSYf4HnBiAFCuF53J/bt9ga0YckBPRpnvBb6rvhdgcy68RyA+bqMZFYh7FcTBGg
7qoD9vLigUfNj6JwVltZxzudFQbzZF4l3cIeIOROyx8Qqm0CppZxMVuTTQeUlMQd
0Dc4KXdZwXLn0HPDCeQJm+lmtiRGR+mSowZoS0jD4OJkjUwKEZZZ7H+5TU3CmkuZ
/2qEhjUjExZrNx8Iaq8kWNt5cI7JFy7Mm36p2h5aV/h0XtQEc9FIvgMBWf2mZwFU
G7sIda00g8fYuIW9LGNZ/p/qUd8AJ82iuA3hIFRpipnyKJ42O2aoinEke04ASilg
pYoGSzUIdFjwJozGOaMWyIMHo3KSQnpZLf8q7QkCJBgYvxnUZPH0W+m5mKBj/fIa
6EuIs2T0vv/lZ/0urB/mfkUtHkzLLAU0CUzTz9tzxGcxBNTDaGz/OictXp60W0mD
Vr7LBAwbxttUzDBCGc/dua7wGpvJYx8djHfzky/s2e/WyIvAARfh815crqIcYv8C
ZfbFynaSIGyClbSA02anAc0Erg4lKs8WROFCrzaKHXm/EVWHssUOijIoe5v0WRnE
57o5JQoxvDhfbmB4N5RGHcPRpQX7bb9mj8oQ7gUcgNBH14oJkv4gDkZeSIJGdsBP
IHoTzBBytUFmXs6oM6K80hTXkM4oRUJfUK7ucHbtabzPSeLOi/OlBhSKFIrWBode
retRWt6uGuddlerO6A2YnCA22yrmTS7bk8nm21BRJhv85bJ9RHnwj/dVegcls0vk
jXezo2x321hKQUuZxD1z8trVnhUeF5yJR+XGhkESCATBv5vHr9bVnzZGa6OzJzLl
G43+JU3F/DQ7OHa2CQWqJarj3RxCPS7eAM1CN/xbQJ2/buAwwjJv5Z+zwyPtpjFg
xrw/isUtE4lp6FhZe+n+dOul9ZyIdiyfSh9kKelQCaVRlibjKr/Rwqr5WA7f1ndA
dKt2b8LQoS6fqDJFEWKjErs/mxBNQSraayy24Xh26saAZjTyHZukHkS2GOR6VqW1
LJYMtALvzwTosELtjnnbq7AU7RHs0Pa4GHsZ1TTxpk+vVcSFysBb4HJfTHMUz3SW
vRH555rgKBMzttgF+z+sVas+7WhRKEV9UqFl+cv/NAjAfv52Q9PCH8n4INjNs3k1
IW7LzL/l8F0+Emh83ApaUqW0rmQ7mtHMm6uw4LNC+74wyCcGYKcVInbVgr5oS7Rr
d7lHB0rOqJg+NBaz2Gy7K4BC9oQErqmCAEZBwxcGHC7K/hM4q4KiT8SwBITWdGto
QTaVUN1e/lBg6+jzvD2w1Nq2xS7cRpmPOFASzJ2pC/JiiMyv+EEWUrhdmjumzwkB
2xype01Q4IkjnWWy83oBZmBjvyNAaD/HAK39UsMBg/SfVNNXZacMg7d5Kbaa6tmz
DlGpGW+PKYY7HSQXvWVnZOaJlN7LIg4uqr+gYTsva5l76giiiFEuo9FmzRJgqfjR
72/j/yRVo+kOfjdNePVWWxWwZeh8EsIRpNOLsfP1P0yh6gi6u+KLbLtExpp18raP
+4WgdFv/lxRErTEYXq5JsUW+PSDubV6soBLNIUutkMEurzoroke4tE2yJFwKkGwc
hkAUT3eVNsfTM7NnZJn1mGV4h9O/nX9tqbcaG3/DZhl0/FsEP6vgwQPWB18vOPIf
mj2P3xSP5JdX5kjDyHy1sJlvUNEf4V7BOf4UqgVsk1HmxkbESh5+o0B3MsjRQrOd
Dy9GvPLoyJxr4o2Y7jRctZVROSjfIK+mjxf/+QXH0niXwBj7eMNl+Pu5vtmurHzV
BF4XPp6K4O+nCgot/AK001DMWTjb50vpxWids+CT63Qb9JL2BY9scq8OOzrxwJa+
J2CkqFzVWS8yFHegqsZWnM0Tcir6q6lmOvLol5rLHuZ5uajxuFwV+v+zQVTlzvdc
Nz5ddsjCIRTJqeDMDX8tv/XgXAy09EJ/O0S+imbF4a9FNJmfw4bNmGvCcwsnViuY
cZRnXUDhpebb7OqeeHVxrv3Qb5xbk6cShQcHi1SLxpSs/W6X81us4ELy8VUOVT5T
jIWJTIZqNLt9JLM00IjzezNllHCedeESV8x2iiW0yDyiZnAp/RBVDVS6H2xKJTrS
rBHn0LwEx5cuj3XlfwIPUGVfL8+E6s4NO723YznYRsljZuYp1W9ZJy8i1tueZKTa
COrU5PdAEnOJaEMIpAhjwxIJk3WIcjVUpGA43KNy3JoIx7BP36ox3u8C+I0qx5Nb
hVI3QSoG9PKfqLDPFKho5Hj7L3PVQ765608+cBFqagz9wt9AaPymwBUW7rs7MuT3
nYutkmDCzwGWtsH8E86oBdmpluat6CxKQ7bSmXyfXmyVQsZMV/Adzhl8LHyB+apg
ZEAXnlDLL2/MBwvCQGH6j6MDODIXY7GO3ZV54C7gc/LFqZHjEe31tNiczcsrItOr
LThOB7Xx2y7ZrAwQ8D8ociWYwcbMuZEhYepqwHDDrvB3XKgHB6bnhLAN7mm7vltz
di69fm32ErTXawt5ATOxOoukhdVy0t8Eip9d3kgy2XwhNeaNrTEndZdVPsvAM7N+
WQRolZ3Btig8Yz6jNKS3PXLZ4tAc2P4t1ZEw1UmPINXKyNTP9pVhMEK84KbUEKq+
cE3WX6htv121oCv+LogPan6cTdQKmdhFcSDD8hxj6+rQx30nH8e8MoI8G1Mpegwi
0farTx2OMj43D/7eiLydNP3YOV81krlhSSUV0eTVGOtevz8xtnAcfSIOVtKHPIM/
V1tUKHJ5voK7dce2K0TEHitnRrICzjfiTlMyJCbgR82IsPYJvLY5e11R/09wkgwO
2hMrg8uoH6JgAKDIaeE0ZzbJZAxJF55XngeNuG3q0+bPYDwcCiCjv3c/Se1u7fp0
9vN6zyWENo+ceVOiYF+jgFEDk0dKBKLnY47y0K3ABylsMQtEfyyt5GHM+xncqALA
8KKEJOez2K5I4W0WfKQmwavZs5QwpBg/kUFQpOXoiMzYHyXoLKy38/4SoySRYb7p
krNQYVgDjLHaypdy+rNeQUYgBGQbZbS9bYXTZS21N1JiPGMMWmPyUgnz8UqbziJY
sT7jjkBCAo+tjvBj5HJs1br/Gy7++ntRnoJrJ6vStRWrA/BFpmItmsgNinhJCM4s
1XKGZZ74Ep2qCDz+4Re9P59VOVGvOENYJcs9KolJ68s5uA0x1h/0YK0vbM2LSgei
lWdiMhv3KgYVNkpxrGjS1syKWuCTwtPTPsA71ZSho5c6jz90VkmFzh+gOZSnXFkK
0YYKO8cOy7QNs5Nqgzc6/cOXtOoJJuSAykpXjT9K3KaKqLiu69Jh0l3TKU4+1A8s
ywCS409pNU7cDX5tDQzOwKb91UxNEsvuJijHIrXBAOcFU4B1zkfhX64M0eJr185O
kv4OArd+Lmedk+EVTQpKHR4wzgbFp30jI7zPdOCnrAymPs4P99gGjbyf8KvLLHZL
D5rrlh43lY9jKYbkq8ouqozBraGe03Z30sS2xKP7g6pagioYppRijcEDKQjJaa3o
gc7Fn2eb8tDOKCdbbuXr4QiDGYBQoGIEscf/yU8nmvtEhEp8hv2HD3/xGC1IblmH
L26X/YUXfIYE8xlujwFGp6bjOzdqyrmRYYyT33gbcxMu3bdkZc3R8BvhYK00ltT9
kewXlkC4ZgTzciQgyLiAumk7akoUUEebKIANfJSBz1Hbg6gGquolOJy6NbHaZYDW
a0gSZ0QqkPPbkLz0HLif9msGKKaERh0sTMj1Kry3SXRwU/aV+3zpytdeW+kgueFY
mrmX0/K8Lgukhy6uIhV3OKrojUEBX+gNox/PMzSc3BCUfdJIpNTCAJcv0D2N9Edj
Gndz8G76l3+c4q82e6dBsL4Cph8XDrFrwjfWHRep4vJPv+ij7Y47+VL+CI2ZAdY4
XJC0XZwGNFmdcWj3Y/VYNN8E4PQPpPgk+Lu07jkBiT8GD6UE1St7LnS8/bztUc86
4AbNDAiEnaawX/mJ/W5SeReUAQuv5zYsFQ1CzKa6I5wIoeptNPNihGVwIUpYwgE0
j6Ftpz0FCcJlF6G4ZS5btwWGFtOtCOIYSHeUYEzGczgqcQ5B+Dvo13EVS9YAOP8/
Oq0hTzxlzP2s+9xOG8eB+9xC+/MG8pFWwVK1tTA9GN4a4aozcZDFr88gDrQQ+0Va
aVHbTU7xzynISwuoK6vGJXyZ+KRznt6EoV6tXWm/6QGVV5cNeOXe2ulFunj9/NPx
9fE9/TYI2r+d5tImW1a+4f9h579/fE/erZUZY0SuStS7kuVpZOGUv9VbVNaQkEhD
Dx5a2Unr63Pe/VHnP2JbHbd52t15BhFL2F5T4Bnx0ysht/DyJCljQVAykoKvnw5W
6pDXYVJ4cAci3ujbvPDsUoKl3p0SaShk4OB2GNdOizGjtOW7XiLmlkWnUwa/mvl/
bC3UEOzLNWwIBC+D6hmimveEOp1nnNnxO/FsMvLGRDVd+mKfZ7sNzgWKBbpmifbJ
jFLJX37bPoHpWM3o/AAX8bxBU+jXh4Fff2CoAIyvsSqUoNT22/0HpLK/wLeH0TMD
l5Smpo598mgaWYcYRSkTtlYMGQYQO7tnMV5gLrFmkyzdVQi2ilh950dlx4LG9Y8q
ncGQBY1UUXK13VECgP2HHgmIA/FE8xQ7NoWmpXCTBPenC+SVuaVjA7O7oJ2WwqGR
A4yf9D+EvodSOhalVnmfB6oYHltHFhrXum7radrGVhG71KMUAIBdS1P9Unj2j42n
T4Nn3DLa0DprEA2udTow6lLMQCejqYB020OcodZYsTfPG8qI537vFn8IbVxjKe3a
f5pdoBE0ARpwXPpGUDfs6w06ieXDfvdyjgzGet9BsEb+mtg4UsCD/FL181HokuG7
ZU32ld5abbvzYKOV6/yN0qFjPYR5qtKI9cxNZcqkjBdA8MSK58v4z0aJNfyNidkN
kPAQhzv0rCuqNQoenmWjKWFAyJISffEcH3MIsKZcFosyKkC9YYz9tNRTQh8GHqKH
I1EPpzQCGL7NtC7M8B9udbZpZLUxW2Y0UdnIbhGM61X25skHHCr94eKd3PmSEHH5
6sZtYgXa7pXW/g5wTgMbcttmoM8LSwnpDblzQkLKqVb/sg3QHi4c6AklwElnpBhD
2uYmcLvb8+x0XNyzOPBRpBNhklRkEg23c+J1nY72ZwpCkFgLshsWkRHwEK2tUeZH
u8jbYP3GlUgBM7wp4ONPtGl81sG9COI9a0hCDxMqTi7HK5kKS1Qv2fCVlDgOSkKE
ElCysTeb97j1xfnjPgMIumULtCh8HYlBqCEouGCkzGUekjphECE/8DZThIyna/3S
k1u3NvrU4KIKfLtYYbHwqkug9OJcLKdI4rQFoJPO5565n//XpEzekhBO47NyCCkV
bDQp/3YvcCilZsb68UxxejTU5DwwWLcYnempZreQ66g4bsCoqwRwrhYuBBdnxOFx
BALt3NJ9BlsA1gitjyWNQNOtYeBm/BIel/uFN7wJex4GLh2bL8oScMynbDj//wrR
rHFRS/cLm8I5my7cc31Fl5UDFPkvYMwX5zbFqEWdkZY8BPM6Mn8hb5qSCVWufsXJ
nA31asGxyfBSdGrUJZEMZsBTdOEyI74Km+GUBYa6IHx61leKyi0TIFE9S925Ri2e
MZxAC0jy85GB9F6yP0P/PVn2Ecei27PZ+N73rL9/xrPE6Mk/3Rf4fp6qRSRpek+7
RlWAK1jpG8h2v9kotYwZL5mzaLJgE/gYKVNnxK1xhgtiZL4wYjOHPRyRhlQ1AQUA
c3lhm5ETki/E+WZhRQeipPsa47dkUeLUxwvX88097kdnfiIJSTlk4A0QXcRYjVvf
3U+gAzMtiThijeiuJ+/lv23bvkW8h6V+G8fbvfYDrmHt4fwNblaz0ocWzd7H+rkt
twuvLVuYD+XVHQyQwjUUt0LedTsN+go780TXH6jIT2XENVaLMBZnrgD73p36MB97
DczDpxgDQCDHs0R6xO6V/5ofDHnUhgJOaSfKgIRKQFqfywF2sR5Orv1Fbp2DqEWT
UGoeprZqQqngm5FGuQSCmVRljDqVkO/4TEnXVXRQqAJQiVdFhRc2wTfjLDOmbJHP
6EUUL6vblK1Ez1kMQtuRsCXF9u5ia5Uh6b6GODLcKMCnp7usxxeYrRnYnbtdSkQD
QPBr9juOBZrAibEp4mDKHHqD8+pMrnX3wEsz1RVAdl2iQgFwU10el0Bq6BC9aDe0
5VRZrkcLhISaphIO9SCYA2+GaO3LYpuUzfjcp0nhLNsygPF5y9ba4IxxlG41n5dd
PTcPZKu0nU77uj632JxnZXLvcvNgBEwrUhWsj9rrh1Q9Gc0u22bxKHYfUIxVeuf/
IGtmJLHXZDjg1YelRHqATCeukVo/3u73l5Zzpy37yoPp3Bg8Imft8zerR2mf10WS
3wfEe2+6KnIZp6Y9izhyGw+TigF7w/fojVBCFVxJV55nGw7i40i13vWvinuuqE48
YIK5pVdu7GJFdbZ+wR0EEyKHlZYTxXkj/xbV2NjaQRsuo82k0TLLkYP5aW7JSAy9
a2L0e/SEx7xPciZSD5J0tNktvu+5uXjFS3UgP0e/XEpAAdDVSul7O6DP09IPX4iC
uaRIOH+6woLdaBUhDqxKSKfXrrgffJ6NYyS4qUpBKKYztMJJhSC+Qtmd7b8ln1UD
YAFCkfnFNEI/N/CvkOM2KW1OtZW60YrrpJekdpsBFcZDehdXE/ccvbIzsRGCLh/V
0i0l6ebw1ox9kUIy2z8PhReHPIAaUeuvhfQA7Lc0+sGZ/HIKETnbmlWRRTuOhink
7PXSgrJ8bzF1uBCw9R8XjVNIdjQ/5X8dRaXOAiDdcd9LWxuEdPnfdac4X/3xjkCn
KR9FPYaudO3A8+jzVYq3Hbed0C70c76cX900+nPAUR4a2CO2YeUD21XLKNeihcrR
cUx53meZwIUOeG3RiB2X6FWZPWDTcsj4jLTGPR8hORSvGFKTApvZOoSgq95FhiUn
RoIntJarV0ROJoe7WW31Z5vCmxozfP/J1oLF4bFQld7qpAWCCwlXlpZPm7Fwh3i1
/WPX08UQY0JcdE5D06H8VGcnn+m6n2567NL5UGggz/tjXfnudL2p1Frjs6F5W30A
heXP0AJrioM0tm8znnqU9bZmsg24NKmsS6z2R4mNNF4WoxYGaTXmu1tw2edpqHyq
7QLyL06O4omXV1ROSGibsmN7oCC7AZdataWvFPuwCXNon5Payl59OzLDuDIxRlBq
QrSYdpn+UGKwLRd7YSNvxXJ5EgyOrN8U1dByTuTbTLYF0TCwJycqEKfVqCqQMpZT
NGe9JvUJ/9XOEUYwNObujz0Ez0B1d+cldjPVpM8/GI1xcOyJp6gM7lhr/Fe8JsBJ
PkVN7/bqCPMlr2Q9xnNoYIXZ2BRC0o2pHMs49tWzmptSfW23hg6+cMYM1/qhZEcW
YcTukvgLM2DkzjOgh6P7iAGITMzVFqm8Zj5dcjztLWjDi1HVZbpCsuZy9oL3/3/9
IqGvKCBDWNQl2ZeCchzwRBWlxd2U36fbwiBF8YTXbCElUp0/Ao36+AXp3+jBjDPo
BETYS41gUwhqF7/vjJn5wFWzE0vuflghp1RaNGrnyxuaXbc19BdYcquFTg6/4ky3
kJnYeV0esPCrY4Z2kaWBLxEi8nZ5xHS6f67SzeYHfNX59yBpoYGJpQdla2a8x07n
ltfNmLtryFxByNwKgGUWDq48p21vlK1PbGPUzGZDFhTFnvG2P21C/9E00ggf3k8Y
YX3yRSPXpTajOBfnnnTgBp4l9jBz1vlZotkaLbLG4l657CFbmNNZ3Rh+jA8AoIq5
U9MCfzW/5/GHKNab93vkmgvaS08PlvDclbPZN/GYZTpGc4xPF0zXYWmxo5OuGW3t
k173+hrKiGRAvr9cRTFP6wNhLVRCDHZlve+5QEL4B3an6fNsPi3HdkgB0RBVwruX
jmuozdewzMX36JmAKoC6yvc0RwoGvfEjVbwAngXAxYrzIPZy6qqkYu9fkiXwQxWS
pklvjSFIkEI390Kq0pp9Jgk4CjlM/HHLaDDJjg4TAN+maj78iFTPx3+TsrVyN669
MXftRfchP4rxSkuy6Xj1TGb0gkrEF48+JWCKIXhn9jg/dmxGatlpysWAHqu+Km/V
AgRPBAsbi76EBQJbzTumRc1dGOsWJeX2EYiUjmWDSsPklqpBsWAMelAKCkCpuSe/
nGEyVfgScAgCM8EtBfJmIn7XAQxA5zqiVFv8GOJwxkymQ6/U4ZQ+u48SM3ySxFil
x8Id4JBgFn74HqcgbEt13Pe9s39fOsDQdQPtK9CjHfNSR3Hfx0PrepjOa7npzdpf
1cIhCllQbxGqZqpH2GkzqX9m+pscxt4Vqy7TXEOYmQUaMEEYkhBGVCbWrrFMs1mi
ErXBkG6K4iJOoR1eG2s/COZvbfGb9KaT2lhmwNKf/eWbzR4C32Y307/+aBc4d1d8
RA+/Fnz/1bBO4qJmBwAKC802HVulgDwUhzc7dBtFDDfTaltw5Y9WDJmQWb76MuFG
kg4/MNEMufefQmEx4Px/+aCWqPPraeW5z4FXGE5f4ZVCeS7kKZMu4rrhYYDoEGFa
UzFJXjZolQtAmAMX0TQU/B0Dn6Us6GPVov6c7rurrjiddPZP0TNNDgNn2dg309In
ve0aCiNDHDcbEUGIJER+NOcLYdJv3cMoLL0AfOHTZ2RsEh5rVPQnlpugpMshT3It
ehh2/gYdSV7Tp2HJVv98HSdbniOjAmT0QVYbrJJH3G765vH+lSeE6nn7diPetkqM
j5Z+MCG3nQIjpaz+0p49XB1OCuKwHHeKrDqlvZVFhO0+9UuGzY0nzT1A3UCOSb/M
oEQS5T7QOnoi7i83QxyhGhhNRxoH/H6h+bqYzLgoLUxwcbZduUPGl/cKhfJTC6Iv
kBTRMmoI2lLd2R9NmpVGzj1UcCT0GA9/Hu7NdJ6yxjLN+vSaUnJHo1zKau0bCXOA
RPfAjFDWSR9WW43D9Sv/sSaMV3V5zRhPukUwOYJA5+xWPUQwOP0xnbs9orN4/1n2
TTtPevtZX051wlxiyDtPa9Q6TuZ8pQBfruwltbS/9uAwBpTzpG9IqXOZXLVf+79C
viBa2Or3gp4j0l42CuQHMjkX7pe+UfqMNp4gBbJRDRzhucpOxGWhptTSJdjith68
dFiewNUtutcakE8hQiLkfl7IbwNbyx7iWzEr3fSa1t/Y2cOkuKrDQWx3tZZZVO+Y
ADQFrZy+dpNeM1bKY24bPQ8MZgQLCWxnEME7iZ0fOMSqfa99ipzyVrSl8j8Hrt5D
KoLRt6szkQ6h7JmHDGkJO2Y2dgVRVJMgM5F1J22Tl7LPNJnNI8m22dQUbwS78s2y
WDhKSqxP2tMtUOSPK5BnARBpQA+a9s04sTpDPRYzdvlNhtKb/Bbq/daL4tNStWW5
C923hItrUlUvFd65fTd0QYmT89sBRujTEPydPbPENOFHAqDlzyM7lxSQC/nPMD3Q
drX8XKqxUg/CWkuYwCAvsYaa4Q8b5QeIImBZ3YixlrlXTfp+WWr8PNnyIsyovAxO
L29M+NjokmyzgpoauarIsdfXXfuxMCgRbPrdU7D9JzOxnUCo0xDR3+bs6Ulue7XG
kT/ZyddexQJeF4YutYcrz6rUtaBT1N6D4WPnQE5IJ6eoBQ4e4Cy8ZmgBPQHLYKUo
Fl0PFSXYZGcrZrApb/S3sx54sx63sCHAbKArQYjEmiVbvVPPo+ctpyzKe5ndT2y7
Qtzbqf+XnzofFTTTj3hE+dbz8kaTuDnioZW9El779Qf1xiQIbRq6Q8ISzDuW1xaU
Rt2KhVqm2WqlqR1vmmPxbFJrALYBwyndPbT9KC5bhSY+6HtrU9e+2KxECQCUkfIt
9c+YvXOEysrLfreoy4bQ26vqhG4zKqJk7Bpv6k009E2gIeBXe9t7IJcsygyh8paD
AgadwxgC/zX2pZSWnw2/UH777qk6kK3WYYWJ9O1sFPOo0XzDRBTMjwsFzfi8JJPx
KcdBt4Y8+1tlpKDTZG6934Zw4pDFAO+6gQoODg5M4I22U815wKj039gS28Q4DjkR
1DIRolF4SX+bdYfOsUcykyxA+iqxM4zXawxepJiZh3FgieS8stisffgpJQfibDvH
8kPVGNl/xyIBQCvHSTeogxhdLFABGFbXDHbCZ09HJ6din+gQbakCP2OPho0UOjgz
jBPw38BMKgzjWn4MpD4dDl9RosrOiBnb8mwaU7bJrmdMnVEr8STuInbfrZ2azK7l
Zogq9TY0WZUQro//Qsxjgb3okuw77YPzRVDgJWGTu/pAIO5VT86jBh6RCJck+Qys
nJ++0EBBIu47cUZyM2Ifh3Yikx04HhdpBkqciuITJzbQSom2sZfG+tzQQOv7sHeB
MlXqD8iemMM9LhPuaWrs6m8/udP+/cefnxo0tCuFblIUqgEto6Rbl+qz/faIJlJ4
9D0ewYV/mtVThRV3nJTKYxxwz29BYbhdVR+5uFEzrJ2RK2CQrcWLKt4xSrgs7cgX
eprQan44CiNqUlVtKFbyjH2/PyokJmX3raus/WHP4sUKJOhrPic0zIryKQb0VWQh
a/QMUczIb5i6LSQd7ftiATka5n90JKt2cN4h/BGjejqnFTkDp3ZaD7MClxU8/hVm
3lwSxI6xzvp0pnhmV550fNNE391QoUlC9vF5ToGI+9qYIXLAo/4W3Bz6cfPn+EoX
fU86aBum+2ONdNXb8xNrvJroY10t1qVwCw1PshG+xGEYhtGe7BGaqItPinWpyK0w
rfN1n1Wl5AHiTZ+ZVsrrt6v8mCWWQ+6EVHog8umBCEkUJp7LA7Grxz8InJnUIwa3
HUyBApVEnaFylqC8a1oTj6FroV89tMo1WbRr2WuNVU5HU9dFofDpTJf5k0RNglxW
+Xcg43qw+ppcl/zpw6TWmBvwPJMMGmNvJSD+RASe7j1j9w2MdnaSzSN35ii71fDi
SquLXtN83jkWXJUzVawkDZoB0/z1nKti5H8UbyEPkQ5zTjI9X7oQ3MSfFgVIsPh5
aRjKl1v0C8lKOmZEHTK9L6NXNsKw1ZoLjDWlpg4hLOwcRN8b/LBP5qFLQwD8yPG2
YQwVCQqxshTxkPtaXLC5RQnJyY/zU+wh/dPeG7DaZUFVx1vudMMnL1o34jB0Kmnl
59mN/el2oCjz3nmUjmyXLQNRSsiT8DTavMVyLpWiyHbZOzK1YhEnJ32cIZg8rsFF
x6PLJLqMqhqJM3rD36oWHgwTB8nynake+G5balUR5M9QjRqRGGRDeFfRcyRt9Epn
evWCWYmVql4bprlPh8aNZ05pbnIhmYJVrFKRQzkcHLTySlko0fjctN4OPtepKN4C
RsNt1a4kdlfVKD1CBC8kfXUnQ3Qjr7GtS546njuWzC/xeZFoZkc3qwBXb8QmIx8K
+KvNIZQspSGJcWBVYiw34FsmhSSmd1hMN+rjdy2CZ3JcmS1Ckwl5TGftWICvr+Ws
LjRlFJoHFoc9HtPB16cqIA6C5ZBFwUY63tGCDo65rJQx6EDlcPX9Qv2tPM8cLcDs
mhf72DKJ+MqgVHmeri6rd3GJQz5q/rBZWLfCmQy3Al/YF/GvcUlgHRUpkLYBELM7
i7xOze74ZAqvfb7IrRmBmAbcJwa02AH7Fq9wqNs1oHdwLOzSF9cfetMXpaiNDfvd
S3Mkkq8eCQluSNGYNQc0FZdFBhtQW8Kds/ZndNUOSiKFABfm561kI1KEqETJqSjC
aPL3T30P0wbSl2r5VZICEHk9+R1G5983gcp3LwE70R8tUch8BZdD9A69xQgcJIpk
mpuiPviZOTEYvy+hbV3JRNVq5fPwAaf+a6707pgtWKqjGuahPaw8xyBrIaki5Ukc
62CfT6cO63ICj6xDxAp7QmG7/8Vhvz43hmro43cKFPOptoL+UpkjDQLS7lmyFBlK
gRARaFhyrTiGeIh1izERkoEclnsrRLHYTCavmts65MNpwoIyypd+qV6dzE86Fd8z
B+hkIbpof/40xSz0PeNwwROAUslZXiq+ZjROhZ0u0D5gm8EekAMhm09xFX7eguB3
MqX71ZH4JKOY1dVmXTG1kJoGazdVcYo0SNuXo9Y3aiG5IuF/THGq/v6548vbrw+1
FbdIxnrUJdTbOITF6PJP2RcDoKRkcWObH89xNOr9blVZwm/hXscxuzsXFgBcrcRs
bsj4G5YitlbtBYxQGeDXyeJxylucrhUpxEsadCSlYhe9ygrzC1YEbn+rGp/d+EB4
ezcvs7uqHSvYrGsNuR23L4v9MtZU7RIQR0Na7ocBNYcHUi3QYwjb8jO8Z5V+i2zc
y8ImIDm+edyyp5z7JMd3nw9XLuxQT7lrAZYkiLvzkPext/TVQdUhxWmRSJvx4foU
jz9JVfqziAQKPiGIlvOb0mazhx+VkF5R1Kfy5Yc/rhsJ8JvvVwDPNtuWQrFjSLup
0uMwqmFx96dzi8lml88GvvOOYL7BvpSvM7RpxuS6vs5PnCWZ6oZyMrIvw/kh7Wag
yzhAmxtx9JFwi5v1IIbQmOu9avLc6IKHGL8Re2gBwkrVpioXLR+t5v9D2VQ60PNn
9i/tjj3eAEVdMAxDrX3j+OZ2Ln6J4NGEASvPu/2vmRuGu0zxKTszTW2mWpdpekcv
bWTjult6aRrT8FJCN4YLvz9kawGbeV40vYMjmLk61qlIaHJ/YjEmRjfL+f/Mrre2
9ZdtN4PVkBJsGGSJqAHs2as4Pn+WmR+9ZA0JEDIvlBJTc5oMwPq4pN34HXXM6TRn
r4ZnyhKSolTFMKttXUpwLKYjaL0H/YXCgdhP+BREe+GwpHLvUT56UIfOAjownTVR
F8H8zGOnztMrnVSfFOhT54w0gvQkJFpNfu1MD3C8/qR75oWIQ66FKMXVz0vTqdbX
x4Iz33tUw0tb1kymKpSkLUVIFhvagx1A4KXhL6Iv7T6hjfb16IZtuJWH4xdqV90X
+lZ0J12Juf+OxwoXazdjTKA819sz2trxmSsaLIASe998+pmc6angztRwIpB/2LpM
guognd8v1If0Uy77Z1QmDWXECO1QKfVEv9jz3nkJPFUOYlw0BizJP7n1QiB/h0lJ
tLYHOUpfNU66y+gtFD+7I2CeJjpAhVAJgUwUHRzlr5hUguKni5UVFWCL9e5oE3qS
7tUGJszoWo28HaV24gjkwi8qbHV0I6gKyiDSXAzL59qElmFIGoiP3VgDKuKjo+p8
PTvFS5/6Dh2/k+SF6aEI2YDRfDUZ6/f8C+RDTWz5aBSq64wripjBvOx2epOF/6zU
K15VtOoZ0lAq/4nvyJ2k5A+BRbIl5lG8IhXLPmOgWEKBKHPokfJRpOqX2n6HpeGX
cwMJQMFUnCeYruYWp9dB7BqG0ajf4e8ATngPcV9ROknip3JonyFeE8b0oo/mah2i
awrxA63joltSvyEd9pRUqy4k7iJQWv5Bss0IgAv2VPohWiC+oEgQ0uqBNvDOAkYH
lUdyNBlPR4UJlST2C1Vjvpcw7hYTwxC0UAPyrM/eyILaplVQiuOLF14PoRreuI82
PJ7Vw/MxVAbJItA34OWih39NHPWEzVdhV+27tA7Ym3Q5DEcIv+viYlRildtK9AqM
QBCR8E9TE4Mgk1yI1cC8tHS/JKic41u3u0E17rKKDr/IfJ9A8/+o+S61hA4Pa2Yo
YE1z7U6yBieQOJCuX2LMJRJfMsaFl+jrwE+5EHWpQyo16LgYF0atTcdogpaij8cR
OPW80s9gW3cUJBYPyvEH5AWWCddDSSY4ciSWTiU05GeYpw2YbjagbbyBuyZ06NvT
syBsAVNlphEeYYabs5O/2sJmteZ5uOv2MFlZwiceKkORzVv2GOZ1t2bj+iQtgRFz
qvxreu2nTK7tjvRly2mlSB41xOnVxw4cb05AgVwL1+HTbPSL4kPr41F0l3C3QhqF
DNQEylJYvnhbWaYHazh1gX2qvOt4cxgAQ+UFH33oBs6TbQGTcjzZ8v//CfozGZyN
WXSJMp2rIvPA0T2PEiUIcm7eouPcx4tREZyv9ITOIfxpSmqZQDg2FYPvOn5khiuy
KzlXlN4BmVGID6esFMJg+QLtAnIad4mZJOg/2QaKINDAiywNCR+CQHj3201ukWyV
0CZVTJmkic/ZcpU5WEZXZQYpXHs86858l9z5vnWYu3eGSR8dS20i7goaSbNfWJec
FiXeaqqE83d0ezvLfqZ3yLXq56ydOxaHfjtbjRJOabILyVI4GubDr3pNX0DbQFug
DCq/O96MksJzqcUbkEk2m+imaspqbnFjpXL+UdV1jV/qwQ0tBOq2jTuBoaQtDKJy
EkPl/1+s3xyW/SAqya44fpU4zhfJ5Khy5ITtB4AtD4YERncGh1N0wS5D8xjKCrXl
vbpk97qcMmBT4cp+ueaX5jG5ghfBZtUbHEnpN8Vlwi3D9eG9fdb0RHbEBARfNC+E
KaYM4OYTQoTqTBR/6mRVGY2tJBFrL3EfD18ZWXb36Zlqg7ShKmRDGh2jAuFxEw+y
pyWR9+uCyz917zohxxIaG8Z2IC7Sg8wEJ6nwT16O5w9sM+Y9ilxXZdvfW9gztixx
fjvcA/L/NgbSoz6Yo8lXvPWJ7gWjQIfFyNyjrbKw9gC/FPiCz8ddj7Wje0QAU6Gd
lzOpOHLDZOG5584sGyll7LB9vwBLj3XScdw3BVNSv/YXY7CwdsxnMOmzy+YnOAop
JjaexDgjPMV3xPaEJxV1e7ublAq9zMzofQxJzDvVt1mTDPCNpZcEKJfNJA1v10LY
ebpOrt86oMOC/q8ZPtfD9Wb55zhc3fZKgWGIUGoBdE9EsP96MoQkjM3jn7aSpUqV
SJZ3MGbudts4397qFdGmPu3xMufsLUucVKqcGrpDmcdfCvP/cdrG2sY7lq50paqp
Qj0KVnpseTlbw5n90rdhFslj7MeCl7VJLj+cTp3QXJNR5BFQyF+EtMOEH/4rEyFH
HhdhsLl0ryDwWk2NTgbZDM6Vlb7k2bPghoCuADEEK2YbKmtUl9DWyUUodtUYYDT2
D0l0oj+jnSNKjZ04q5fhcbd2W1nyiCqPnAb0DArwakEcoeBUpfYaPYGu71fJ08IQ
ppjSoUK4zozcs4xxX/ShOGhJFRfDWDQI/K9Vi2VaANMguA/8C9Jkmono0N+nv4iF
udoT0N918VZjR5xv+B6Yip6xY3V3SktIec6W7QYzKp8kbRTdzkmvDzZKjjeLmvox
6Ql39BWQJcItmC2LWsgPTDc8zueNoyZyvqIbFOQBIXvsTtaijcEgE6Fz9+3rwSiZ
//B8UYXHlOIjnzl1P/g9gUHnZHpQg7FAjgnGOOwEer1Q4iitImWRFTJGjsqmLo/G
ipa16swuA7Ax3uluv5KJNyYM47aTI5e2RI2kRPjLdwxjqd/ByEpQ8UzrjrIuSYuA
F0LvE5d3ImpQ5xUKaPbfKFUnDFW3RBCSMebCOVcXNezqLY7a1pp+gVmGXTY/gAT1
2B5s81WgvdfEG1MmVcATf9DfBttWY//HMH4Iy+WsXJJ4QYMe+DuenbirSOxOEANY
F8dXOak+2KgfTZG7orBMdoNGTcyfwB/d84/2oFPV+QWLcAcncQCm2GNnGtHy3eHb
GadcR2oSkt9NDkMEc4A6LymRJ6ACpMiCXNJtj4MpupevFTd/Ni6OMrkoCbisgdg9
EFGn2qyzu8Ci88o+ANoTeKm/KaGX5kZP7MqXu+eO27vIlVwqMrwObrXCvXhm/8TX
mZCTENeHGz0dL6TQiOqgzFuIpLXA5DrWIIKwROLsvQfffCnY8yzhqmKGpnGf4iLm
ZF2C1eifs6C/PWZH7uEMTp1fRtSVpCebBNgjEC+9AP4tKTFqCQw6VkZFGuMJn8nA
wFIxz1CFDk3NUgnWPs2ydWFaltKC2FyTc6N4deW3v6wT+dVCbBlzzf+TW/1v3tt4
TWI7k9SiHbSwYptl8gvXryuGB8bR6tdukASoQhS2S5A01MCDxKCn0SRB5TitMf7s
XBUisIhNTzkLesSIQGe+CXOBJ73mIXk81RqiazJmD+p1NWKcq21lwNpV1B4cQDwr
mUHDiOdQipCMjNIqJ2ZPGlQJ0OHjj6Zku12ib24Wi2/5fC05+hqDTImJuCUKQghe
+RfH8ruiAdXCOO2XzC26QolCCpYJtkuR9/jCT3cJoKcm9acsaBpPEOlXKBsm1h6D
6hgakoTTd2O3WY+7YmBuHKJ0U4w5ovqB8xvQNv+EReoD9DsFAnEfMGY5hEOTQ4Rz
W9UnJe5dOnmGgbu4F+7r5JbsZnDhPnVixwosTpd5x08j2SeWiph5mI8/X3ozDk9k
TtSm4+Q1Y4eJN/2VUI6vc+f9fcRsMGSKegpuTNCkFdSZTRtCT92CZenuvrp90XSD
OfmFfiGsbOpbK+RD04TTjye7Y8LOGglQBd8uoyOvd7JGtLcrBVsBFfx4GjnMfvki
lnF+DqOOtYfmj9nKjVzx3RwUh/iXj6/2z9q8ZNVxp52yimfEzTC0pMEdV7pw9kiW
YIf7NvJaY6BbKOg5BCHTywuSR8L40t7W9dRtraYF+1bEYBf4DqlcSNBavZXAe11b
iWlLDRyAJRWAkvlqewChbCHTNUdrRrADdZzwBCOlxaDBjpr1DxuCVOcjVkEgQr0M
NEmHUVlpao2R6dKbANjotAbmrGhIUkkK1aqZ3DljpOyV44sGfwgTaVs4l4GOHt3u
fVUoqfBxdXIXmOxw5mibpQuxN2ojNuss2CoDUF1ccfSvAuCKAJlkf7IHdk/e/XEj
Ly9H+GwZY9fsUIbts4TdenI4h86UL9bGjaFQagMMoYoGD5VTipG2e1Lg7Vtp4ePn
VwvSiHVFKi6iEuzE0sejCyXnTxJSYyHCwvVD5yR/9k/brZAsgYioqZ9MC6ZtLNyY
IcciJvH0wO9TxvQVAVC17UwFGKUWhnrnUuGhoHqCLIiCBKKrGI7VfFo8+ptifKon
mpmICzhN4jdLoPs5BYvGVuqYMySHRioFDGvFnoPkX1p6FLysFd9iP3AnMGEJnTRn
jFVjGf73EsReqaRnERDA1uAzXI4teOx1yJ95oZRlVNKSnlz8iF1EfvdeMCFwc0bE
iX0TiFruvF4J9fFWCwRi03zVO/BECWKx1nm6Y3xoQV3dhXU9XmQvJL2LUeZeuO4x
gqQStJfhZ97EngGKWzulK6xwYNR815yBFauUpxdE0SkyFM72fVrfMou+fAiR/DrV
nnAxbkW1btNqKq7VsQzeNZzmGgDtKPk7F+TtB8LgKXoKA4U5ze4THsurt34/fNQz
0TM7Uho8i4YQ/IRSq2MU4KXwTh/AtqWVgZRHdYxxN2ISu8l/y5TwWpuJ63+RxH3a
+aYLxG/lS3zqLlkykuzVSafQzfE2ndUnIjHWxGJ++kAihnDdSBZE545AJ9RkxHPU
QExciVmkvS0VLNHj0EvE3uHDX9twKKUe1+xnIW5VnWYmkjZ3NpVbTPE+EokW7hiY
+hiwgwCDNVRvFQj9iN0Ive/k1tF4XIPoxVxzG6bgYP9sorU0DBTf/8ehh69E+Kp7
A8BFNlWc2zFNbYGhibiCZIv+NzksdzitnvE69D3o00ZqotuJN8dGiCawqanFRipg
mF9qBc8zYjxzdXTVLtGC+NTt6O50K6QTYf/D0jmGgKPmK2Qq2kRUGCOsSyxmmgzj
4LWMc6RAX69aO3V13nOErQkDHYWYf8cXLX9d5w77tWkDG6W11HuGFWO0Y08peAij
AkfSLBrIirP4FVPeMufn5T72wnypfm63uH0yi+iKz8/uEKKwgyF2daopDrZ2SR0s
nOXh4aX65tHF6aI36qFG0bKNhfCOsqRxMOSfKOlLHD5PIiVzuw74B/hTcNBW6aHM
IEaJwF9c9GsjmAXdwEdlbUxMhm0GxFcX0Mmtutwrazlo9KKkSFvJY4/X0hpa2lcH
Qnw6atqsobxx61db1/tvdaikr1FyBP1KV0JldJJKfX/XqeLrXHlX/hG2EU18EF9r
U8Y4/JIsQUaSzw0K30H90eoj9b5n/tbzZqyREbSqsuC1vV3ccOn1FAWzylo/C3GS
gMjmTJcvbYZJsassu/IHGzHiVW3GI+/B33ePC84ZIU0p4n+EiDUPFk+HOk5fwH1f
vlWuJITgJUDCCFE/iEfiS90YJXgYdaIrIKnPKqXltWgC/oEpfQNgyeiRwhOtFOab
OqNRxgNMURlxcYhzd4bimpfu2WS8J4RSXPMhh0TtjAAzBIl/e0kQP2w4lDt3gGNh
t11WKHyGqwkBagHeDNVYvxuE+SY77v8BiRwzRfAwY46gAIothkTcTXFrYr9zA0Fe
0oappuSH/rkNjv6sdDAWZsFMZpeoakYtsbOYW5mfsi/S9AQySgBjPBd5DNxIOSnP
fU3LmERkflsGwVbCMf8rg+H44QctEg8uGttaxwn2COlnGjWvNozSaUusQN3MW0wB
wl93UMWifwWvaNIfHRYwUe45CZuH20jhD34unVH1IzvTaDWWqM6QlRPk3xqLdzuK
kMVp5HfL6dMKEIhebijvtfXwi8J02kKWUmTqxXkLzu5deqGc4TOVsoJbd0lqWmWG
XgnsRb7G5Q6Ug7EXTU5xFYkKreBMogZTn4L2/riIRUlsQ3uoSaMdwoHJa8A8O5qa
Ue0ZdXypsxxzcjTmkoswxI2tQI9VfNE/GW70xTnHf9I30yu3VooNL6DI4r0Rc01J
EHRI71eEUz/qJkSkgE6bBeHK6y1anqop4CkoGXGdZqrmgc7mL82aoQHWbY0xcT8a
6KKWO1CrA41pH/zvs0SPdTsbY63isHeQST8mXz8ls495wkixTCgmDcbxesE22qo5
ZreR3OpeNKppGM6UAIrsGO8e9RWDfCmm1sVlGyuv/7XT2hxYoBWiqfh/30UNUMK6
K3dgk8vPS7jfV2hcnOxTOhZweME/6wOSennhqqLSGYvB6G2fIdLg0PR+fyVj9XSz
Q2bmnH3RHw42VjAHaT4Ht8VTFaO2QcaNIsMvXCYjBmU8mfpkouS/qD57XQkWfG3A
9eqq8/G3usd5z8f8QfLAiKkyU3RlMg16HxoFMAw7djz1EEsKLZLMwrga+kNX3Bpi
KjwIiX2CTOF9wSnYbWVKb0/yyMDx1O0X8zkRQSWqrtpBxxRwEEytUkqEx7W/xmM4
k6yIX4x2/+muh77uye/3qPe0TejgHWligZbZHOXR56y3QSDLom63ZDRCbQzAhCcT
BcNjU3oTKakMTUJQdyjQadlfKsTlZHdDzSmUOMMTb+JhPP6dhstzA1VDuQ65BcfT
uAkiv8A70hMS5CfP5HhpTg4sZQ3noR+K5Fnpcv+dpLSyJneHDvDIy8F7URTU4UB/
nzL9Pm5aCZFNUguE9k6ScX8d8ynmOl83kwiEH4UvD0BUE1AqVpUxcoU1mvHOFCQG
bu9azzJ0uxvcdfkAyPOzmRmNqF4kSwcjSGq93TRePs5kLKfGK7eXdIVnR8PXqnvY
pS6+FfxgcwtIdjWfIxwPKjQxVqhONrYBTrEgkIuo3LpsuCNQz+6QwLvQkHBwH8Dy
eT20OYFbHUHAacA7JNhVzwaga80UZt7/Wi0flPgvTMoo/FtLeLMjBlP5w885dsWY
d7u1XCXv9JM3Gi5UTcG0DwnuBwFjnEXQ+Ph5M2Fl1pJN4jMFC3nR4A3UqnCdING5
iZY+eSJsLj2j5ZOPezdk4PCTpkbFzqwckqEDjSurNfU1upzlLi2lBIa0iXoNy306
wGqZ0lGRnc7owTpHBfg51K9BZeEVPjl/A8/hH1KOEXI728iYe4nHFbn+uOXh9qd+
q7v7KzGK6NH3HKwRoUFYH9UHkbxJKlz0Y0txlBXxXmLr/ePXW23nXooZr+pEO4Kw
DLnuecZzlkL2KNf7zCJLTucSfLK2zyqE6b26w0YY5OKgXK15laOxN2UuM1/+y4uu
zS9SSERFiPy9qXvA2LaffrkhXx8gSJxtuJDPjM4Ywp/ohGyKkpAH/hXqVgYj+yLO
3Yj/3u9QQUJqrIIla+qC6dsZK7pI77YQW2XOtHznyne9Zo6lzCsQX/b/xJCUBxQs
IqpoHF/RNPBCmGAzxMRHKKCxt9ZLkC2T1Pl7XaAhyt+ep8dp0Xihm2GLLPukS2Ws
flkZX8oaadrVvcZmBbtSX8yQ6IjJo34Or/za7Cih99NqkMgu/MbtXYIBVTIufQ9f
cZwZjgViRWYdMC1ZNM8tk96LW4/khmGeIlCB6e9qHbM+1yYTUig7WY2tBzRVj/Rb
vQAk3OvEIO5OBX706czqYSj+dP5WzYKy4pAZOewF3wfCqJF8bsAUTprteKISH2XZ
jGRj534evzqizBRu52QxHPreyDlwy0rma0oUNA0SmjmRU+QuECzhNc/w3JJbsKyM
i/X8oW7tfBmVpaDT8nIZXWR5lXwOaXjI3vSmWbuTeLZ09D8LTza+wONNnYceOg5X
cKjrLZQwxAYKX/L7YYZZmQKTzN911TJO9C0HIv5hU1+iE9ita7Y9r5REXjQgjnWa
h9mnImZYLJtfTpx9UKATfWCe/ceXtKWAJft3/ZlHgLOBntgInEiEBMN+jMIIMeCu
BNl8q3i8o+H6cnxfmqKzRQbrn4xgSBLs96cUnTJZ8obJSrfzSLIsWFnP9YRFQjfv
soYQeF7bndLlt2/RLdHVys/mN6CQQqjS8qwpXUA4QxFQbMvmP8dlcenHfBL7vLB1
Vdwb0q3VG5Irwa3L7JX9c54o14DgZhn/kUeZbMQiupAASKTiBDO5sLPh/1l77xTU
9KjQBM9lgsF64HNmpPZrslOpu6kkio6XhiqOoqQl40lOsF2kHpCLhFo+raUk8U6t
Zs5S4N8+dEXo6SrMleCr9jncvA8djJVLZRqsiPBbUinloGFiGGpCxeiRhhfoSsMT
OMM1LbCNch+ZHfrN93RmkyB6F1EbZpubZOU60r0k09LyIrcrGAcy8sBIQrFKkn34
0OIP9Pu9xnDLZ3ZqdJmAgCey1ZeulNs84UK6A4owASMxGWa/J6RHbAPErPGRyX7i
dS2r0vO8lvN3RFOYOaSZgsakjwC5devwU4Udg0uddK/yXdvQ5MQh9bms7ngga37/
tXouQ5ZnR0r0wjoj9EjMUs3DtpP1+AJhjsbn5hD18olaD6Plvv0dcrr4KCrEmlRO
XjTlZ4vzPrDgjQ0Ri7kwXK+I4DdoTOMt70dEFsrJ6JTtWiKrfNLYe/MmmzzLoJoQ
Ioku9tT+TOTiMSA4fQbLyvNCheOKWAn46cDeSfzzaUMyZfSIgrg/i3lMN/JfaL/1
NHbiksS9t2F7pkylSw85RF72ZyodQTwAtxeqRPkAJCLad3fQucJ/H+4BxaWE+Nfi
+Ee7fUiT75Lj7uFkvoxrctOX2SoqZgcWqQXtj0ophYisTTTfnyvcdWRpTtrrR7eR
jTRHWZpf5+4GUsSOq16S76AgL7GJd6O/BJWsF3EIha4PuB19eM2Mk7DRSY4dFNUB
Z1ToO54h2pC3OPYvtx0Up9ER4LidlMit3fCA1WXNBnQm6QwITuNfPCeWw/sFvwZ2
Xk5MurZJTFS8b1fXtSmtzrZ1bFUwm7VuO+00ORdo1MFdvtaa4QRhgHtTthOr/oui
A0HJKIXAN17VOOXrWivUqfDLViwWKz7Z3cQdAVm3L2Pbt+QIkELDul2GzVGJpfyv
YHyeDk837nPBQH6VPuhiY6BvOcHA8+Ji6IyAfCtu/R2RAgBXEZtFHNUNIvOU337T
mjrxOT1BEq2G4fPR1cNCyHiO5f0zbjXEX9v/LQojwuYfGSUQ1nDXB3JPxCgawD4E
JV0m4U7QTnt+npjSUo6OcmSepuoroblK7xaKSgjg5j5zfXpk+OHAq27i5Le1Vo7C
Ud2WzzaQ6ip20E2gDo2hmFRoYiHOBEWTjca8s/daNpqq6NIrPkbYkBQht1OfKtgT
TMMMX+hdGLJA4zNBxhaBLus7nm6gumK0lYPpXYLdI5HEBh0FC8NctNCwRn9Xwlb5
CaOZpyE7Px18yCkTeXsFBiNLPJ8XbZgzGGsoCs6zbU27L6qlnLX16OUcxT4DtSSh
z23rtZyxNLAorUEKdd/eHqaZe45IgdqdgiVvm4dgXZ+wzqtbu41scul63/GyCDam
QvjmSPUABVMXPDmeOVq++r45JLlgt7eufPVUzwy4G7rBH8E8/EGicKEx2RT8RHxy
8leWdgiVMawHJ26giv/fskKz5IQbywmTcRtaES2dUB3p8C/LcVn/dSVslrUxUARv
iFaBPBxMfvaeZ4kWrGLze4uXoivqUJo5GHkeaW9wUNryau+lD5wcCZG9DUp+FZkO
ZDKvf+VUqC61n7lw4ezfcPzrmfJd92rFqp3G9AGGO7VAoD48ltmsGIow+KPvW6di
RSgG6j+cm+wfvfU1472QCRroSwcrF+UB1jXqnBvGC/NbSsf4MOjFWj+9lXTFgLgm
ra7ITvGRWJ9SXtICNMG7SOterUD6SKtqT4dS1FnTkAUwgmvFtYU8X5d8y+JBomRX
GReVoXAvVV/3Sg3KcH3YEReJLnYE+anRx3/7WsVB494C9DTJTXUXoMt0kprJ0SEa
qNNv1ztORpUDbTAsMrq6juSvPegIjsjmF0NIe0/UPMGsWuTQ5fGIERNBUg8CKLde
70UB7bLnNdF7LEXKXnBSCOxLKLTGPTcGsjjbiIBHODghBRNctvHQ4a9zQsJPaRMD
+Do+IdxrUzoPSXcc4ts5Phsndk8sQb3bphCMc6S67pgMkscCnOzJVrYYBzbYGmvU
fLMrwWKk/BMjC5eeAAutrd8ojp+07SulP5/rnnDzOP5iue8ENN/Ri503bVpocV0B
bpmQhR0znEFzzOVhHCSjsj9Gyk9WoMGtQzI4UkJ26/2uhd9yj/vwIGjwMytHQgdW
xMhHxv70wv7EpdWlXijh/BU6SegV9YlzZmQdyx14qgDz8lb32tS141OxOyXH0BMC
X6zTBLVLwn9f7ERVIMSYy5V70VA6i5y6FhsrvsqxM9sYHwm6havxtCKcK9g7Kuof
XNe9FnWvP5vkCqymxd2nwwtnc0EZ8wUYUNHYhpDUMdPTxA36nlyobGqhr8PVeDm7
1Dv4D6Y770x2d+Jm/1Z1SyVIZzCjOGIxOF6XEUAWoqUMmzdOD0Ea44FA2kjl+zhK
an9i9tEmBP2N/k7zoPWLTPE6r5Pm6hC8YweFvvsjwNAC4YQvOQeIVWWio8JZPv1e
GZr0wQ8bnVnPloxk+bsdxvaKwoIpTRqGdXse95+GzalbVU31O+vc7HmdL1EI5OdX
zT7JE/rtOJ7/UlR3CswIu8UBCB8txWGt8ZNYTAvTLOvlzxW7ItdBuuH4xHEZ/XWd
9vbsNFt72RYCWX4Ev4e6Cm0xHMGyJQV81Bv/eo5c0IfIt1c9FKIbOMvev25JBLCj
fSdUiMNGx6AC1gC5pvY2TbcqT1GeRQAptAMXxymXKtxH6JD8TXFumICi1ylBJLuS
D2xU71szNHeyLk8D17xuVI3Jf5rcVb7Byk70dcGAIjQ1rLOJ6ElYjhEiuvZjgf8o
uTwyTosgZIubj4FlGoy6byYt7k54W8un3fhAF7iuP7LaTfgrrvm+irDKXIv4h++J
C7w3O9XFF8IIFVeGtwXynMWpCBn1Rjsw4Xu2m7MoJ8JNa4LRyNq0pjDnuJvBzEKE
WfS5PGO3aF1hTdUwX419dQKyl2cseLiomZK98THGj6SHqvNBJlLaQ0HiIg+ezzz2
Qb2bQqSDr60+QblJqN2r4FuJVZHSONsuVTLhKZnoDrljNNgVINx30yZTZTLLvyCW
tCU+yVvwpHofF3bp/sB/MjnqL9cz6JP1KBX/Mq/ltKBZVZdFdA8j3lIL7T+wG+VN
LEMl0LyiEEkk37vxUujoKkxzqkYL7MS17ay0mRjMqM9jISQbY1RN5y9nF+RguFab
2lgcVuWj76scPRrOzTMv2LBv3YlttlZJ/ZRTDOY2iVjwk5cd0syB7mBBqNmeycjB
9rt5NK9Rj3ixu9D1JuhaAY6t1o5RXlsSq6UStC14Ci069Q41hSlL+21Waa3xKpf8
7+qBKIHVLozCswCmyORrjBCosYyCh2I101GbgIhVvEPfKqPj2bXrtLsD8zCCeI2J
/7W4YFYcZt69lp0vWqkXtZQWIuvU625y+/OtMrLVRoKyl7q6/JcuuBvD2tob0+fD
qQ1095s7kJzjRV/UBOmcBSKyrssTSE7vDGDbwixrzCICnCi3/WJh9s2wKgwHszKx
DLs9hG0Lbifzz3zMC9mYPswhYXN5ClL0vj2mXOD4t9kenL+Kz0CH06eklX44An7T
h6eUC/aCKDfjOSeKuJ1+xfFLIlNvrmXGrui486Zy85n7GoBG31qtJ+SSiI9SOOpl
bp81uAB45x5Dj7rD2Uhll2NmHhpzhl/0EmZfOFrAi5z9r2mWEfupX0jD2q+O+tsz
bjecre99zvNlRj9r8u/nXanozVXY8xTN+8lHbLpAUh62nIZLbF5gx3jp24P68onw
R9uV5Nyj8BpQcYyPVi9FkEWpipWzlKgAP/QuAz5uqd3Ly/c/JD+fBnQbXnhEiz8G
xL2jt8XYhAEiOrkSY54ugo+7wJprEKbzcP4nXkCsZgEn39PeT+/16K4r0Jl2NRL8
xrbCuyj0r7GmdVcfpAVRJBcMOHWItTnsg4Ibql5dD5o7/y+Vob1bG0HwIHC04upH
6uNfaSt+3XWFaVwRkhfZxkDLni4AU+0MBR7d7cDcGSMMEQ8UuMBnOHBgQR9aYCbX
CWa/w+WKrGC30Xamfy1HSzmo0AfgNHxHMFNJVLvXHyHjE8VP79+xb4nMjXVBYIpM
IEEd7J/CX388r9FwVzbB66lXTLqO6LvjtLZ8BHR33PEsTbWSEOqGLvA7V3Sw2YJ2
7P7pgqrNvBySMB9j68Gu46TdsS9JJY/kUJfEfHVN43kI5hBhOHJZP4kq+FWQl/9X
pJoS1C9owoD9spZq06APkV+jARD1xAyVPni5+OwPgIE3RtwQh5p82NSaTFUA+3Xc
ABrV+8eyfuLuMuYUX+dyDGka3X4Q0rjqC5byCZizO2UPxff0Q13z+i7YJh6Eh4Do
n19v552VBZbR5fpkB0V4/1FrTPIs9jBBEdpqxPaq1UAgd/4PhXBVeJhvd4gelVa2
H53rziejcWyTU9Phf4IkKixQgFoI9juUD01x2bAYdpDekorqwpjDHNGX3IGG23Ij
vgMdl69avnnrSsq82Cr2xS8Bk3RdPFfwmBnsTPGzxj7MXXpwRTI5A77QsDtpkxv9
oFGGe5ISqlnMOpUurKy4CpHzKgAMW9U9y1jplD+oMInEvRXMx7vat7o8D41keFu/
0qoUdBpgw6hOtBK8ffv7lSO92316Dr3/a/05ZDt4dSCnmTlyhXLZT3HJsG1AD0qb
IIbkBzu75PT0Bwf44Pd2GrvfspSvRTfNXNxqs4Yd4lfkxIVpy7GUKIwInmpVpiEV
P2/xpuAeqYBvpOAXujUko/SK7+0pnyRQ1+QOt5s5tDQvRCr0Abg8XnoH3b64AqgC
iWzbjAS0XJ+ZW42wyUJpZFka2sGJ1Vw8aw8E5nWtfHD5lZCJHxbZBfkFbAcTDymT
50KsUptrzvlhF2rA6/hZ20Sdz6kcRMkdRvD6nrBsWuSLun6D8eY4icNq7AIShxtP
JQn/TxxceQALodbHg37IYfT2vUPWKqp/QseYYe9vzg0yppSZdiGuKN5HJImaddm+
1RnwKKxFzcpLPpvcMFH925N+HEmIpRPizVt86w0K1BAvgKeJ9I75G9VEATKyK0I1
UR7tiOmGX+q0Iz5DP8BTsV9aPaOtVvYkXFK3URo1n7+1xjQ6tORjwgUJjBxjV607
BGJ/weHXsdBHdORHdxtP1B29mGoYNzbf/sJ3oJZsfkZSEow2AlcaJ3NDUw9Uyz5h
IjKhe0PX9oF2/47W3CwgccV5jpqvBu0X6ISXKZWC2bN4N729ZiaJQT436HlMdZRb
LV8hZ3BCtdRPYdzJT8bPBlg5R8aFgv4Vw41AiUu+XnWpilBAG7I1ws17dCNQBEtS
uuS98kmg/1gAu9m1w5wo9eovwuNZ2l++wbVzJSRJKKMnSQl9+14799LwVttlG7mb
SdDcSWcfMJHyezUWiQiIh4VuqOCk92O7nx3MVYdset+m7yGk8odLCQ7gMq33NFeE
6tpI5krI+/l1O6QZcHH5PSxllmkXsv7XSWJkTV3iRAh8teUJx13IyMFzv3VpX5DM
9SdYQodwD2jF6MieZmHOJjRU1jHXmKxOhawrFCjwzOqUNZ1QeHEh7b/7bqTslyEm
rDNlBsyt2H+nyzyfxktuGvAlW3D0JSuaVjGQ2af6z4QKWK5bYLF8pIGrJsdhRQjs
ZZkKlj4YSuqJfIfWzFMW/8WvQj4eTx1oqCpwVeGA7i+IRi70KFT26hCYQVca3kwH
jm3Id+kQk2YTEASwfreEdLcnu3A8atN+S+5UqpRacrTnx8Kl35tCco+7ZAe4yC9H
WP6knelbk5CZy5ICFK5+tvqWXI6AYEpmBgEn0bcRq9rjSRc1/HiIb8S+KLmZyBKN
KLcW02D8vPqcuu20GRSQ+VOs+RKTEIKgidGl0/CjPSurHJ1bc5bAf2ounrAkpuVz
eFHjdk+YLLCx5hdfXqtIuBjtvvNyu0ybruUlg5MbsuEW6eA+Jr0y4GTnW0roYtFv
0LDkGZI0baJbohBGqLN0FuhN4XbqZ+fUMQnixyKdeu8uahZa/ThL3ranzHx7ZM4y
Fu7N7JP+8djMGzboqQgkoO6Z4gZUn/JIo4sxsWiRNe6VuOMtwCRHaCVFAwNDCSjg
a2e77c1qsZWVTvj6cjaYttMIASmpakrA2qn0mUVuxYh6QDMH+45XBrT4CWCwxyYS
efhYztG39SSrd7a/gpzGx1PdssjieHQdm170jGJP5/8zz7RIrUvsX2k1oCif0ugn
Mz+XG8Y2zvesAgbb+N6m64nlyyuyoJeKO4Ha6+Lh9Hf4jsoSNWxGKwMQSevWC4fg
iIQYvcznRHrNoy7H7fFCPgQOrEGKLTqec4aLIwrgf/MzDtyP2wqia8SJ19ZjZ57B
yhTexezhSdDdpU5pL/29If5pC3azWgGvGKxFk5NYAU/8/M4N6/XiR5ghItbpxmJ7
Cncf69xnCHVUbPsbXu78DZxSVadIjRbgb1Hda6ldwyDvzU1oAi/v2L98SRhMggk5
KTIO3lFBF/sY75BbW52oGVukcdaACKrKYjBOzfiLirkAUXF0W6+fu/zvgq8WpxMI
xqrX4gzUh4/jcpvWy8aCOSaDMB58yuLx0JTcSpC+YkhvtPuEK+X6XMTRAqB6uxrW
ARNOQPhzkMAlF1Hg+ADVXfQs8RnNDow5lM/l9lgaCkXOiusPtat386xUI1OLRbwF
3Ngvdy5rDYbmq8Wb0i7KIjFhFw1471oVKfvKdxKuLWHKz1FbpmA+LGj4m/nyf50Y
k6+9F9rC/bQIlmWbCZ3i8hh0v6/utNa4264EzyRRm34IOoAM6AKqR3KDF0shfUVy
lWJUgXJSmyImeNLDTqjYYYbNerz3nDhMXPi9ciOuG572k6G02STiJwWD43UIvRrn
Vwf64UOtHcMRhv1zm1v5w0pI07lzXZqZmet8dkkInZLMpJ/ISil9goIc4J+8lxdt
H0wJA1DJZZZWpSh3xVqNO9FhIOsLzJZQuXTPknZCaw2ydEsMmD4GjIRyIbBEJJZW
C/df878orqYRBPhcahtWDCMi9+ByWW2Fb81C7A7xRfDDYda5Lt+JAMfd5bG81XXX
wr9SGpAwmu5wuaaSERysvAeu9ZnQfG06rT/R/eH4+waxZCNOd8ye6Q4XxrK5r7Qa
4cjfewrw++lsBqMt9mSDuH6TAai9PvTjOzUAke+lKd1ni5o1Ibd3UqA6lBmOLmoh
OyBSncN7rZYqXj7v85DU7lQKbLaaKMXthaA48y4u6mEA4tSsGhZDU5x1cNLzowAX
v0lfblJ/0i97b4tBKfsQzMS6DRGRtfuVhB/hsNDkdxmgn8IRsxwy5n8J1VwKjTxH
cFDFl/0sI10spylNpJz5xawd5EWhbgGgO/JRMMCMp8i5AEr33v7RNQ4LrokDzKy9
0+hj1pbBIUY0/5TpC2OI5Tnsn3bZURrqpdYuFqjKk8LV9st7oQ1SmEIysgpB2K2A
Resp+e5uV5FhSpbZaXGf21dcWySXRII83Kupt2s/7rswON0Eq5ctcUcw831q7D2V
qJa02TGryfkvhIYBF4gJNfhlL8as8rjAt2O5fjfPfbo9Asi8eIFa4Z7nafdqE6xC
AGHzal216RlG0UryayIegHg3B0pamqUaPEoUhDwl9mnH9dqYFI29mJ0zA8tosr4s
+uivh0RFV5TDbvUwWOhxPgmJvSICN9JFUKW0HqUzw/XX+Pan3jcKy1nd/mduboO5
GfKuBlK5E90+N39GIuWEmPZRMSq9W2u3yEmL+91Bx+6apcLHs/iqgl9/Tj9gqa9X
ccnTRdlLwS79novU3PauKDHg41fap2hFaGB1eVBfB6gs/Ee295oRwEVXFDB83lLA
FG0/yRwoClKuAKUsNOfOoeISAKhPJnlG3EXgSRCcoslyy670mAL6qOO7kG907+vl
WdLFbyMW9NDHi6tEOiIPDAFCHHTmxMnboj+Yg7HMKOBOOtdHzOKL+LPWH5cNs4er
HdYYCmjwEx3c6FqbORkPDd3dQ6n9giDpstMfUdvZfmZyYJpulrF1v2gzvxflxv1n
CC2+kJAwIGNEqSW+HpxYMqFmLm5z/pbcXG+Ya4IljWMy4NrID4KfsEmFyc45xh4e
XT6JeM7ZSFXQhbZ8SvPs4v/SbI9kBzF+KqN42rG1bqRdzEHB1Vm6h+g+7oxokPLx
nzo+T9m9leI8I16WCSC0PH530XXQVUPH6f9kiDg2TnFldHL59UAEb1XrzjPSyOUj
oVwFnT8rQ0f0oTnNzrBmiMj8EyTfGHEker6RCADgx2LBfLxIPTcuBkdoZLfMqIzL
ohZTFPmQ1Z8fCz1OzHTG4r/hL5ZWHDFxIst3mBJOZK1SJVf7lRLw4OWqSm42Kkl1
uPHoEKXg4FM8HlVbpegj04RbLB8LAtNArCEjL4DYFcj3lZut2/Lxabfln9hUyLUt
cPtkT2G3XASZ1IO9ghyyIvwgULbAv2YHfaFZCcBdopRORjqchbodm+7xUkR50JtE
vHg0oKYOW8KM4QWmQr+sX03yPWfMsJEMsaHE538scpw9pmhjcp66iIcglX4+I4Tk
euJ4q70cmAfagPMYQiQFoXgUIht21/KV0P9E2NrEr8CTQizFOE2oyra/bfTOZj64
c37T3jd0flGc7DWhgu0Y4A2AOKK23NuiU+eIoNTfgpLWw6jC1zQ+jlN/9CS5w1iE
rXrDUsBdau6kiLfmwUGWdnKthjtWonkk+zkz7EzS2RPWSsbMosmHnPHo2fT7SYAh
3JgeL/tevn2VpRAlbnNLGNfU/tdTr7JtgrGVEF0EGQmHncMxkigDkY9+ojTifkY/
TqcMzKo5P9vv02pa0AdxEnjvPCo1UFYN/bnBuzSzS8iQ7Jd6PL9kTAzrxlxqNZjo
uNrWvOw3qlPHH3B/8T09q+mnkIy9/aAW2s9a9982ks4OzXyvcuL6FRxkRqE5jCWl
gTMxpz/MqJdaM2bR6TYk4qMaAKLutU5FzcFXRYVA3Bqe5DBf1lPVVQFH/fkB7EdH
b3avFCh5UtJZ2rIi54Y712DpljM8QbbvN3cSJTfevpRBmkg6zG06N9Wu3kazKSeW
8M/WjS014vJhKXyTiuhJzksr6kCF2wEZNxfG8cgSFI/fV61x12BGIZPapby91/AK
61muJBkmyvJ1nfX1iYGU5ed/9k+qL+uE/jU6ZgAbgAlPH0IgWaC7zxxe2/pHQEZa
AoqvVBKmS5nb4zJ/9YigMwOi0G0kT8jKR0Gf+GpVYx22/MfgDE+ENtuW2j31hI9l
TW/eoSuDQq33ERnD5rGwlzBvvtvH/zors6cslXKcVovgsKt2jvPiIThEL4toaCBq
rlt6lXsz4t3Ypi/lEckbKogX6j0pZujzGAFyItwvt1zU3Ui01YcPJk60fREIp0LF
P+6mxp6GIRP//YzvLqB4Jy+S88k/yPaOQ949DDcPqVPQBuEOpHImGNhewBNEpyc/
B7bwDPbx6fPT5XuGxeZz/zkqdRvXddUtmQYT6bqlA3xn5eHGEXtclE/lvt7yTQw3
6+rBSvQ0lxXwoukpZA23gXGF09W/r9+6HCm3YSJV/RGZZfz6MvcvMHSaf7BCaF+6
DM/uI+xDSzKyrMYQSFR2WO/Sfm9NOjcJ2h03VLYe1UX04pw3CB9+IaBKz0vHMs9z
qOVN6gPGYxJ9Uh4VKyrWHIo5g1oiYVuRe5x9Xo7xPNzv/M3HYh/n8Tci8LuXvarK
kdybTXxZ5S7UfHNdFsx5dvxp9rOMVi4sYT+uoOVRot69/+1JHEZzzv+2q9gUahON
db+7OigL/zIG4MBJ/9ridT+9O4ZC1HThPm10vAvigWzXYcTtNPUb9MGnU1ziz7+9
AMhiWzeTxNm9jR8xVnvyw6+DM9G0Y+CyER6fa3xB/h93JPqXIerdGyiN2VuvzG7U
a6B9m98VcUajCIybUfL3qMgYTjeJWukzYV7wBoKy4uCvJ/RvHAf9ZN6nlc2SJbDn
uFE7EZGrWAuxGPp2pHVrRBdoy97Bwhmt2E7MTPhEAeFcIxj85p//kJtQQoTrkJiq
IV0U68+JjuvuVyjnAD5uXG2qZezathcP/TeK0tzjTlSVWBydWfSl959YjjWAVoPH
xGtmsXooX6qpipvvfGOnNw+qwWazGCCbrfN+kDVrOhTW8MeK1xMAOhYB8EHqNC43
WG4RuEB4spTyXeGe+CMYaPsnmwZo/BE0ObRjMR8B9TmztT8ihFEx8qkFWMSrOFlc
vW1sqsJU7kWpP318TSitE0nF7E6RNL3ob3KOIIELwtabxEDQu5z99tKImCm7ZCng
F4ZRnyw9zmNKTmnOIaLS8EDvvvzbhgPqqMXlTgWn83akhoz+508XPirXqXe35vkA
c4w4hQ6+yUUI71tox6Db/Zgo90rcjegyH88Jvxhs8GBYo6xLaWjpFuOFsExwbP0j
HYC9CxiHgYpwY9jae3SUg8dlCsKJscharvGp3E3qu4Trz/SO28JPXOUU/vdzqHom
msLjAY++xsXXa7n9jI9mXix0tNIWvNac9WBHAcqDm/vCIZV9m34AZKmE2FmjNq35
5vWjJPyxln3VSMX7BwtlxizgP9YuKwivcppe/IHEI207zExBpL1E9uqtT0uB6Hl9
rdq9VobTnvyTrC4lR3lgj/Ytaeh604p2OV9kOJEK1JbS08TJeDtD6q2pAQPZvpM6
EJOr8g+RnH6spruhtZSxNaf11EpbRhL5y9rJmEGZBs3v5Ea6HfJbLIGbElyc8VTX
A/iXZ9U5tfwnq2ub3hZ+7aeMlX1mGsIW7RhQQ6C5Leom3dvuvP2/MUCHJqjS8lvR
pP4XwEOfN6z0mEWry/jdSBkKSZz6MCKYcHk/OhCETOHXRR1oRMPSivVWrhf1VRoS
RxBExDfZTmD+yx473Ro9h0kzOiPU2tgQzMzcI3IHcdihyo7AZBnUbu8XKEG9SoXb
Qu6SIPpwPg38orSyfdxqNNebtXO/HwJi74BLBDz5gohh/im7Xjd0vsn0J8D05RqX
8pbqr07daiaf4/91gCWyjZdsfxTHFp5GZ8yqZcVTo1hZw/HdeEpvcXD6+UyBw3RK
K/+mYAvbxdTJKNCWnn/r5hnuXNTKOGiqc0yh4TOuROl+G+CYk0vI/ie2DslVEeIW
Za0itl++4NrcWQt4+YlCJ76rFDyuXPTFw+zobMGY+ZhMjHdce725I2wEJ6c5hyXU
yJBCeqw8k8c0zD+6VxJId9cFkK2aJrMVJ+Be/RRsGOlk74GJs4TQW807tzEYGvWO
tSk2Oyjzop5fRLEok8Pu6PYHlKuTRbycvfDOQ3AElMcLDisV3ov3qz82PWgEn8PM
lox1t+OfrgTEzW872+gcQRNVin0oJ91VqvV8hYwm7k8ME2mf8kwdLineNIYaFGIV
thW0Nkzf/1gmfnAhj7kFTgt17s6ztXyatrjB3NTHTjbAzJ/Op6zgckunoaT77N6x
HlBhujxX8I4Ex9U3CMANRVRmuUkQMJME1vqMiBRk2giDPNK98jRQmjdqX1B7IF9G
FjsvXg0p0tWmYhi8NsYghHCoFF9Ji96Cef9YrgW4/5wTCl6al8jUf7R8UcpQJuwQ
iXSqIcEveFi6BlXpZEUFW7p3jBwEyK1FgLu97yP/tJQ+VKq9MaHGSkEXM78cspEX
IAWJJBgfS2jSLqRyUhUUA8Q2/aCPyWjy15obhuy7SPM8Dtq4WLA9t5LphFakJh1a
L34PbpjSx2MOSyEakhHQH+CR0ahdaUKz3vU/SHZwcuqruMm4y/eAb0GwpjGfaT2y
ovTN3EBUbE0io59AbyR3lB+11XWRyaNc0jKq9t528zrmC/BInek3xFwg102N8P6r
8SOGt3+QnCTcN9gECayno/wkI//YKvJAmshb+CDAuXeV92gf9fAlMl+6Gie9dZhG
JwxMpD4TquVfH60k8KWeNJnZFLrCQP6eM4Gz93nntFyuUd9sZs1fRQMXdGS+A3hx
nyqI9O/4HQYy8JumgPncxBIpS/Tpvzf5SgkvkuPyZ6jKwErn1BJ9B3aIs3IIEEJb
/9y+jSvlvESCIGJkfY4CEWqYeRW7lq9AnKWdo8PKSePGwAerLH89FxcnvbS0GIa5
tV+wLaIfF/4VyQVtG003wkgsy8C02etWtCC9gxHYX2ERrlOeVCwyIEiIhEQCoNau
r5o6ymMeQiNa1eDUa+pxTQdejZQTvnhhIVEpWq1f57OwVI8SNs90Q40B/Pn0lS9Q
cbEtpPtuj64fpiUdGeS2I5P4Y5tlOtAMx21tX0iKeZNj/ZLCDH8b17ieWj9+NJ1/
3YmMpi7E4YlG1wb+hHFkAD3/wRMDUwb2stQGPtgOqqQybwjnavtl194ZmPryQLtg
FcDKu0rzWdoj2uSXgWHMuGdqCSsvqHcmLdqng1aUC9SdSeOkDHYY8sr+ViIAHY7Q
m2QCctoH+syvnmimxlC2XF0hLL3PJIxMCwmYuxtZ1M43MrjeaC1sgcoy46Zoaq6e
XvponFuKHW1S+P8vxzoLkz3wnvnQNcz3HWiRHzNyDmdj3IU1xnl6AtGJH+2gEebG
bE3cN6S7DHMtvhiX6x6stD/EVjmKRt1b/IKXd8XPTJVZgpo5iiS+Ut63qzaium17
o2V2fCx/LQFvTkWDDjz5tAUxopbU2jWhg0zg2B8k0uPi8ARvqxrNNKUQKLkplfv2
yccnxO8Eo5yu4nBKGrm8jRffkY9elsnaNdxKBNxbS3D7LJAGBuDQl1ZMk1waONQY
hqk39GTpWBHTzQwW2L8W97xZeB9g39ZeJ4C1EpFbNvPS4cYqVhxb9Bmwfm++KglW
E7aAESOvNPmNlwwWYuvYrWBxr2satBTbYiQ5cyJMx8jfiFRfinAek2GX3uR7ZEsQ
tFTa1rbaRZZhpF9G108iiZHpzUucYuQVCh5mUrwyViXi02DxWzB0LVLQPcyGBWbQ
gz2/Lo+GWfRH7WJZpgpyRkechiqVE58GUgyfhP/admuzogiZa6gDx7X5AMn10j6s
EihwhK9Y0Hesx3FrUGQ72skOTm8dYCP9daNoxKyxJuThZA15qUyh6XZlcabuf/r6
C3r/m0dOZ4N3veNfu2GwNrPDa0HhSeqtX+ZY0XwJ6NrQplwB12btjgSXZoUZJtH2
JSVBPi+Lcq9kErwYHy0T2xOSzD9Qp/f5mOcIKmXs0Wqqhs0bjIbtrXiiX5MIRQwL
c4XSkam27MsfkfT05K00MD+VTMeFYURZQXhN5p7c7fBS1hcP/F4NJ1cLyLS1aI9X
woxUgHFb1l/3N35b5Dd0xkBFGxGDAJoY1mO9aCZR3xCVzJutWoM5l65V2OBOpUY9
pB9zpdAmPeebUcLQ2CCyk/iLK90Fsj6kysxMq0MzRF9dJ2igP54i2duVDWEzRSc8
Ngh1L8HKXI/vFCwjRf8k2Dr+Qs15DFX7W6nsieajDmXrJCrfKE71cljJH32j+k49
TcL1DERfIzBA0lBXDXEhSPYBaQNRkaP5403Czs/Q/OXRHXlgSVq8AX0NwG8VejbV
5XXZuA2NkDWWJqc9tI2XG20iHdQqSfpV+XZQa4/dj6EenwnrVQ6OPDcvG8DjDqb4
yIX6Hw2cVeJ+5zzBLKu+fUaWdfecfsJroezhfTJh0OaWmyVUwS2czelQMYzkxxd4
MlU5pYhpjODpd00Y+DIK1F8BEgudMz7SaixRXCPzTz74x1DBsVgH+AModpX+TSiH
/RIGg4solSZJa4WvgxgKPDs5vwsRtI8Kn0t+6/Twx4nCu3QbyQ0a2plCDLERGLVE
YcuXRsNWbSNJ5tUmCtXbF1Q5Mta5MGJmOpHnjb/hpf83ObNxY99PCoEpDPJzHklP
XBINk4zjcPNMFkEQ6sU9sQ6q1crTFYwEsRWc7EhTjKrcJ1PZ686PyuhVp3SoXPzZ
NxXRzdEf5kEDv9Oj4viRjysOv/3KLUD7XjNh7QsBjVOCEc1h2UUuFMhQNOermRdr
ofkKS6KfnlBnwgrcfr34P7KWQtsYV011xMkTprku5PpQxJdvt8/GLbJ4Jx7hsZ8P
GOZ7lrAt0+J3u0YWVR7U8wVzcR7hAc6hGxSUXzDpWzlVunqv2yMpwmUaCcWex37i
deBZSQxQ0nhpr2mNvB+tCFbpFo2Zv9Kkz7Yv0gFgRuLfcma0pnXnGeoPvEWrRNJc
Mf3I02u1iR1xq5tKi6kI09Xh6Qp8JNxvuzsOFg7LF0o2qtx1qRTafHLNC1h1+Ih8
Dx+XjsE9u4mnxFC3/ddqsZ7XKjY4BpNiikjFvWsVsXzEdrCSTBHGqP9u/RJAXAiM
EXi76GtVnS4r+wWAmb/UX5lMjvv51wmb02LRNH3zC58M899iwzuYsvQhEjnN4HvC
+1MMWjDdDObL9GA0baGWPWHgO35f6rnlGENd+CZo8NEvA1yfbo8aA0BSnmovRcpF
zAMOihb5fxvY58zmalxUm6AgkpCkbIoilcnuHN4k+lpwCREQd6IYaeXZxmD74Q8f
b07UMQZ9Lj3JJ0ZQ0xvJOxUQMiw/IK8LoobIwRDzHgznFRybW7rtK9KDNefKBPPM
TiDoYBlQLSOeQh4iztZmrMn7wnZRJLkxlguQjAPM6QsB8gPIVvkhUDwTiciLk7K9
kNuhG7MdHOVbdY38q5iLfpSJXgQNLAN2k8PMWwptVA4NbAVDgmNlh07xQIfJZzBl
7ZD/pT4xZM+shna6pf/BRvxg3sSfyIgdDG4AVZRRlcjLJpff5A+mJHBZ/9s77ArT
vNOsbvhZ1ZHjkss4+6zdE2OtqEbABD4l9vjF//eQbJ/Jpl0i6mrRZjSDpjsCi0dN
aUN8ex+tH6l2/9VC7utmnp8F3+pTd/IBgu80UY19UcdSWbzY0po9QZjDhv5TCu2l
Qf2HOi7iH2/jZVGTeUbrwMz2OmHvMO3IBN4i17ZMMFiKeEYXJCF/9c23NzSvA3RG
7K8baz2MCedsOUcvmAX/mFLJqoAwAuo2lwVlrqnEUHMDLO0mxqYUeGVYrp0VdtaC
mU7t1mYE9hk0gFCvg7pTB+Zn+b5pPbDWFYioNMxL3PQaSDJ2MrwGUs8425HXuYTm
qFYJVFj3ZMafZxPztriBnyLnjWR53Uj6tyDWThEB+4hH3t57XpxVIcKLFQJ2BNK0
AxiHS1v0w+9+po6e5ESYgtBlJ2iwGKAQess5Hhw8HI4OkV5tFCD/YA5WiNMfVaJf
ZyJQ6VmE+xnN2LGyINoDWG06/gjsyOfazqJ8D+JV1fRj9rynci4gMiL8zBswN7sn
RaTFpegyxNz18+mIKVqk67fwBPcTd1SMdVZgpCeUmbylty9H3euDyK4yh1PEAFlm
2p27jL6nA41d1gIfZInc2w5z5UWi5542QMjyjocuXCTliux5HOCfx5Tmnk1i/lht
XOm9H55xEalKOLlC4BBATAvtH2DFtljP8a8NqcugCqtNVU4AWV/+wpLDFUcLvpxm
QiRFtOUsYiZTKF8sNgGnkcPY435hpvAHjL9z46rFLYT8h9xGWMICwbb2ehmdC7G0
RZf5W0cEXtZAd8XcdYeAvrZ6s6TRuhgOokC8DPMQrDfLVn+Ef5Of/mVn1DZmD1SX
3GEWkbETjVJMv0f4PWVU8qnp4Ihhg9Ygc6jRA5QGpI9RquqU+GY64spH2LXhz01T
npt9e6TvShsq1ttrG+eKN9iHkoEmPxOWbp4TNtIGYoehU/oI7b8iGxrLn0oUuOJ3
9HWfEJTFmXfFajk97LtZuK1gHtUDkktN51mDaNWG9rdaBMucNR72wqA1pAIkupWr
8JCQquq7KFtifeZ5WWi2CiW93DSMDFSJgcX6lQHVldLT2nJ8RNTeqZbUoaaLO8On
W2gTpu1B/5UmxCEwqR0gNHpdGQuNtcOX37LjcPsa7+H/xbvc0npxV2D0zNEKPbE2
KwcaVm0uIga1LvpsUQKsmhmuApbT4PH5nYcNPWKASnMbUpL/YtB2OxODRK10V1SG
pksgNHpXBKGx9XkLBDQlkWctOHFWoCabk49olcEh+en5/DliAeo7uJHUvfvCdMt8
+5bILZ3psffo2CcdgQmH0Kx55LVFzXpDfUc7Rj57yNsMQoKU7uzRHuYGsb4nmWHM
lj8smpLZ/DDwKDe80/XrqQosZaxXbGK3Q5VVOVWxujkqAHRY19DejDxUF8k4LMvg
87RfQr8U04TDf0r+x70c6OIITU5gw7VL1xzgVg+xeLHEMZClA4lKEvPEsZqMmcJ7
aUEiPr5bHNFAKDFviHKGZTZyifS1Ateru7w1hMaRpz9uaZaLtljmqTsKjFnHpUup
Cd45dSr1C3Fqz05QThlGnRzdo6FxUtqO1HUPGrvBvhVQPza+utY1jk/CNGfKA/Um
dRAerWvnepZSjylKLhzgBz0ZXKvEpNeW6ylUXY4BUF/REi3sYdN+d+rBt+MeYSbS
+Dw4xGfIWNpfXD4bt+lBIg2pFbm/VcrXhlC2XaIOe0DrACiJV4v88ifraSYBFd4W
ilNjP3i/NplK2yNf3T3NuVQ0g3vFhNrzJNjlSXbESpCBMf8Twu6o2sgoe1X87Fv5
UojrVDfUme6rVe72rPm7+7JSq49KETYmkiWGQwBjrURSRo8/PjOUoMArphOPuF9H
i7ysJ8mY+pOKUPWbkTgBzCpxWPZq3enm0S1cdXJq/nz5V6DsyRvTV4QZcOpWWARN
deeSve73CNHRlQ+VCRqShpCau31Wf5+EvSpOF4ZfqCCw+cMiZSSAMUjIA7X8I9Ek
fFNm/EGud3CMD9vPOZFH1dr61IVEeZAWZ6jYqnxSDobhQ0S6WlLZA7pl+vvW7oZc
CfytCL8fClnBmq9wYa6bWW71Sh0zG5f9+B08eK9v22H3bUI2AuJm4jngvTLMKBD1
J4elni7Acg+cLFSVMbpU9KS2E5yHNglkFYb7HNkk92j5q9B7iu1SXK0ftofz8/dv
1LX6rsnesNyuStbTP+ZQ3YtJ5znARk2wEEn4jm3ooOtOn+c7yqpUCvOWlchfYye6
sc4e8k0p5gYxACkappmpF7POmPaAzTI181bwzNxjAmDfisLslAQYUFh4JCmka/OP
oWzdOMlDeMXnIX1c2R8rNu+kWfNDEOHSBArLYHofTSPXdhz0Vt2woeGQyUDg1frV
qE6XMD02QcPH1oRRMSenVQISPQnNIF2zyXuWAuh2oeNCDzCehVU3X86qIoJjwjnV
/Te1dmOfk9mHRJjNchoiyUOJJZTE0xdchSD8aBiHMErEK3qobeBTLQMpDKwUtXT5
fbhohrQ+Pp8sZf/vg+PG/YA/jrfiEOPaPypp6izsR4HhCSWaAh5/ftMs3dUp32lh
ekFksLj6k5Fe01gR0Iq2yj+HHTO+ozdBJwp7j/CPRnAZdxENHJoHx0Wvbyg9Em3n
tjPh1xFmJkI5l3luT0hc6pjobS2klNEl+ozIBDnsOfq+AqXXV2T8fCukpT5BFb2t
B0/7BTmZlvFmhmjBVPHizGJm0AdJg4IJgGVfHp5883BmVclQV7rcB3ByWrTr40Hi
zXKATn/pJgSq+XVdpOJ8FGZfpFwYC2aaA5N2lvxj4HFQAr12Kfw/Ht5VJUEwezX2
VlfqMDPwy8P/ZvWj4k0U1wuA0ZMCZTOv9ufo/VNliz3KWJ64e0BNsrLoxcFw/7c9
RfAktxd2JtylD/Km7npKBY/WCKnybGFmAOoM6SiltdJTKLimPJXW/FYteqF7Rznn
FK5SVYRwPYHlc0kxilJLCWTa5LNzPCKdcn/hHN89ahpkfSfI65pUaZIadOidqHVt
Drdy+sfEsBBwg2FyqSXuRWn4l0yFqSIcaP60xBRe8IWnKWd3D3A8Czcc0Awn00L1
AJ/vfCpYs7ZuhyniD2HVaylWr0RmZEx6Y1siok5HPkBL6D25ESkV+2rScakcQREp
zgQ/pOmuFpr5fT0vp9so1jN0J/ILo/6UPHEt0wBvMSN3QFfZmc6DakCloMtLElsV
P5FHD9QA6wczo41LPRZCyJFZUvcjq3ebGhV7oFbpuGSC7HoDa+62CRCfoe470NS2
jggnkfZgKAEo0FbW33C8vlNYMOMg/DGod29Z+9NhZTrc2qkdl84XYzkUWBn80XhW
Lg3/cwI4LqlJA52lEXhvAuW1EBV80y0hSyh6Kojgx8aTOZxl8TO4q0IU4lL5qTsl
/yEprPEtaUr/ctHdIbz/xloEgbC33jJD/ea7pzSObh4CmEu1lJ0dRLI6WKf/p4nD
dLb/vINS+MzeGkRl4N1HOrQ0mPLTjUUBoF8EGHiLZO64GL98llmqBC1lAm0kHCvy
cJvGxhmBk2FXNHbPpoj8rzzMM3vCTLVOcO62qrVq8pdiQiXL1iQxs63E9z5EsJtk
Fw2bU/uLRtfofFZRMog+JzRpiGnZ+ypR98vHZ6vS4vr+MbyI3KNTY6LI0SBB49yV
eqENKW9GiTjFYoca92nzVZiEg8jhA4bxOAIZ0Qij9erV8z2RQIG0zJ9RXDjpvkdm
qJVpC6/Y8YJCvy5VxxqTe14x6hVajNhNBoos/zslxbPecS9R1RXEbp6L4DuI+bZS
TTjvefj74s22htY8DMLBaikDIIYWbcUvn18oW40gcKDv7GyE3R77yiHr427bbb9d
23wfwy/QO8Joaum7Lo+pfooFXbd8oQ5f7Nu3ndDhhxGBnNnCZ9YHs75cDDgJmnEt
Dao/sWxdZCELgMqvgrF3BcmDU4rPgFfzPJ/0vTW55yfj0oKrIkE2uVRgMnaZjdXX
YlTyBcGiGkBWN7N0cD56wtUzmxjqwafdBdbZI6ZW7R0Q1zX+o3jihIPM4jT8+2b0
4HP314+xKeJVwBhhCuaIUY767dMF4yKKpuPQ8iHyIs67poV5z3EXiCFDDskTveLV
XBdRzAAEayf5C1M0tK4+goXKYryevXpW3VXkkXRhui3NepWa0pNY8eq/HpOv0ymp
BbnZc2+WMPL5jSR0ZusYu12mBAFUAzzMx64OGhPhrJKELg0px3d8ePRY5WrwD6Ol
1Qx8sYbIOhoiZTbe8l3wSMy4WKNBLQPCfFGykw/HAVKQRIWFPBFZT+1VAmsqTD8P
AXIQ+Hc9WakPIuIWs1XryF9Njl5NSOxkFvWQ/qShp7K+zOhLQnzZ0S3Cmjw1P9LX
A9BeFCr6ReVU6XCG44wMHMu+T1m5f6EBdJt6XaGzpjqNnshnEUcqwgKlp44j4Avm
ZZonDD9npoCy+LGR+GmzmqS+p7EzN73Zow8xMXFEdEnkzqHRL7qkFr8vBs4s+Qid
C8fQuJYgjVlA63zVT5cf8PydaLiV10GZdz7vgF+uE1Ug3Rvbgc2QE4Ny5+Xc5qMl
VR62aU6CnK91LF7HacuiuBOTfkf8hcxY2mmlYK9XFiL6NC6J0XOTVTohiLQzJLfs
CKL0Whze2UElDKHxwR7Vv6Ja7WSKnUrp19eagru8CqeO+ClN2el0udXriV/+fTx3
G9vBm6c5yFv4itbf6TjPsxk+tjDgEI6X+QAs4FVpIgLouocVsa9QdVZ7iwcLeazh
WwQV5+A6RxWho6/EM3VZaY+IRqpzrgraUnPitVA3VzvRmXnKNFBwDTR0+fDpGn4a
4Q1zRen1J5Rvpsp8mSzXaVJhRY7JLqY8K1C4zsKEVeNUfK0t0ota9SEcfR7kr2G2
Yct+CQ0dEArWO/vpbwuBH3fnul8TbQsKeSeCB1O4QE629VVm+lzIYKZyQe5yuABy
AClYU5323wcmDaW38rsLySgSgidGQWVya23rwMSO9tBFOIFBMIXVcyPY/CotElr9
4qH5ULgxBaGOGFl5/mo4WnN529w82uwOyzUOiUBZzAWpxjrVOBFBrtHLmToCi5sd
fFAHtvazF/1jeev8Cii/6SXMQaKPBQrlECcrOtcnbsrdrBKi6Dsr0bJ52lJquHuZ
33MkrOCDFKfrKjuheAPooGfzaMbu2aPcgn4egNX0p/z207AVt3WyOqCnmbimeti1
VE6lw3THPuk3vA/Y5yAWD9l/pRUdJEUD+Y1Rkg8zG2r9YauP1owy7rv8h9KQKTOr
595AmWGHVrjES4hxdmVTrWMw8j4bjUeghTgx1X78VEhoIbBPGL349FN8x9x365oF
lmrKcKG++rq/usm3xuasCIKGr3ybxB5Q7x9+RL1CEnUr+HC0mHshScnYoyqL+Hr+
4e+XuH0eCpAsiD4QKVuhm/RZB8vM9yFL+3V05EA6H6ha2QPWaSCzZMebREwcPdCF
i0wokWJumnN8XQOS1p03E8RnpOX2X7Zl06pBJXREOsPOD1UMVVzfh6DA3w46icdN
+dXeYQbWS9WvyTKkbmX21Tx7UM25vwZ0iaC8mmvrX7SYunEwiTt6chCjYkg0x5/A
tgO+Q24L3K9C0/1Q+UCXbGnQGloDKOIbTSFiXWCLsGqO+kU1fMPX2fy4dY7Dwddx
W4ws7lWag5IlJTJ3Vc3fqUX1pDW6/Qc8sSxP/HsVv/vwX136KSbnHJ7MqrbkBtyb
pcjBhE7z0R0a+lvLeutWnakrhqxfy9kFc1x5aRK0z0I5MT0svvXx7XjJOR4v3hR6
CoCrSZfuwvEtOq5oxmkwAl0DhE/Kpt9+O24oozJDfNFiTvkuB+jUZq95W+32ldvU
K73kNXRz/UVVYk8qXXReYiYd+QpAqYhTABBJkg0gSvuW5laN0KUMepuf4ojgg2wL
3hthYKAprDwhRUod5AmoyVXadRhi4Ceg5aB0gkky6AEyEK9R58rF4gATGFVzKHAn
9G4UGnBfBGsco9b9JhJlixx80k1huM+voXylLmU2YLbGxzn9MsJmHnfXsHiIydi/
AY2yNA9ku0r/nvx9sRp3iSvUz83JqkzdoDOw0c6yo7/97eZCpaIx+ilqO6yJUxJC
pfi76S8qy0xtK2TYruPNzpZKX+5xUjqCIDClf4GYf5NInTOjFEbZBFNahHiH9LBI
N4TRkpxdzaC7aT8y6mx9hCgv/FGOy4beTqz0FT3lRZZjb3pzVITVU1XVIhnhUUMW
fmFAMVYOWWFXYr1VnjFPhjspUdR/8QWTRkdQQ+RidN57ILZwhfVo0in6pOhNi15E
jgg87wa4htGrsp1FDQasTf++/4RaIsIsWUoagHX8rbgpbewb7AVD91kbvi1+V5gJ
LFIOH1kE/Ya/WNVfON4J8bRy7wul2l4wXqfV3D7AuFvvYhvKeD6NAs65euuuFH8L
55KDHS5ykrLK0IqmTzrctEKJgAYSL++1z29YjCAco+CXJ/q1qAZ9vj6Qv1A5Iuex
3bXAlpbqrykuEVrx8ZZEY8Ft2oFjyXqqD6nqWLHKzGf/sASdXSREvZ9xR/t58ctR
KK4vOmpzurFEIcAh6KCjsMSMMg+5SqReemycRHcWYPelYlEU52KXPa9PaBQD4KUo
lBp1qS+t1Uw7YJPwIZ1oaMcl3Id9gzGu9LLrFJUvRgb7HtD60osJXyvNO8ktwdfL
2LXDjB/EHN2tgFXqVxJnuHaB5QG1OtKSlVLd48rhN33BtZMGKh8uxHe2hiH4R/wY
/abiA8Op2XshuS1mhmfxIrwXwHGWfr8+TCxrIeCzeIwuihxqmnQeaHzBqX3viMzc
4Y45IPjs6BiO1h6gtS+QWaHL9ubOrqFtEHb0UPpHl/irsyN9/dXL2Bt2Kq15M9fg
BlOYrgxB0PbPEs6fXfKCfQxqNTw/z2Fc1IgVpDFtHJ7SlcoOz3wal0a4pcEintx0
FkfdoSFjFNWT8+hOFmD9TD1afvgLxtB0yIqFmzwoKLOImpi1BQkomGnfp19DTMdq
ILCmbI0Kf6OBPJnWxvGs4Cjh5CVEVwWHwdAjCki5BKzzop+mQWOQkFUAXNSCK9a8
6tDhqidjp6Iv4wYGpxnNE3z/p3gsGmzOGlwo2uTc94kQXCFWBPgUHDgHWOf63dlc
Hd0cmkIdz51R/7ioAzN1MyHJBUs/TRNY44MnnOTAKxHd2rDH9YjFAug28809jTpD
qls2OvGQm5tpGe58BWdFAkELfEbs6pZ8N0AiDgpb4VIto7nzEyd8XVVXPyFM4oNJ
vits4KLQx5KedlNoLUc78J8usqj2Qb+WFTfH9M1PWqBvZAKn/DzxJv4s8HRtwDq4
uwqvAeeOn+jbNNkD0BDfuxRetk36lgwqBEViVKATCb5OiOubXUDr3weN5aQJ6XfY
t8zsYQSl0n9t+zDJxtlP+UbQuNkao+G5jvWAqKEz4o22FKbgoarKVFPDMcnTlGDm
XNVhQGgKDsZ64a4r0gFF2StAxDTy4frwcoZBu40nqohpoQlyM5vwwlB0c58zYrYp
Lg7XMkxO9L60T10g2Wcl5ReNjmJRx/3zuTkLw9ZI8UcgRuUiklShcxpsRBpWCGa7
ppTpspw0v4lsMcDkihIGzmjIEOIJYufczwztOWrEhSHBDZEoffnn2Ft3sq4v0hff
UngkslSlO7TkiBPViObd8IHDthZn72J5WpvAgnirnk4f6vssi7ZpIcXRybeACv8c
cGoHNbvuu4diINX8bryA4SFt+272kCD2dQvTtR3hWmLHfrtBp5TqdW8QIo4FcD9l
rLq4iJfJ0MvV2DmdIGtpQkinr4MCle4rOUYS6PzwokWMS15TxncUEBPHpc5KZO1x
MtWZszHYfNbcXpkO5x3X1UIKroTEt6ecD746fObxNeOjrbgEKR8ERvOH0Vuy2Sq1
oW3vPKzPEE7W5c/7xWGWBLBPKK2iK1zr/GzIc+oE4gg4BMTEX2eTHR9CxMSBSPCd
CFmQRIBVEb2wHXWQeJLN1Qa9NDQjKMUFeTCIIiqarP269ENlhiFGJaJ4XsZpODHO
+4GkGaWou4yxmWOz9UPdMdo2qYKmI0qI4ckyjiG4uEXOXY1zHvGUBe2AXsxvsP3o
QxmMw1MaVVZHIvxWftBE8mQJOoa5lHdb3O5LBHpl6rpB0sWezWrJn+x2E0mLHtmG
KUS0Pmmq6imvSlv8wiZO4E0vYD/Rx99uApdztmVGLlg+pMclg11ALEGqhphgDDmS
ZW2v57o+UddGia+RElZ9v4vxZlKaF6NzJWuaLFpalHEu4XJvyVNZSvTFRE3ATI9S
5eEcu+KKvI44gRgUW9XhEbwCvTMO96oDYl2VIarptbQ1BysDD3IojqnAvU6ajVMS
i91Fp2WzmltK84pf9cgu3hsUSfMMwrQRiSQDMBg/HP8jlFiu9FCNTTrqHzHU+273
htnvZlZRXB9nqE756hEZ50iPr3hRCRcBYeTiJjahGau4nWAOjX3yn19Y6DK8eTc6
zxeHhQqf4/GoWiIAdWfv88DMllJxjh4r98QiLfjxliCUTUCnmUY9U+b2THrX75U+
/EiD4Kss4SfWgjRO2sWu6TH35dGlQkI5fuK8qO+wYWt/ToQamgW8i6oMYOHmowbR
i4K9/tlovEPpH0/Cyc1wecry3OU4ZmbFYsxB6jWXba55ACN7RjDcK87uOdQweU1A
j3UpkLYm+U6m8F+J2t7a6B+avAefpTn85Z8tfgbZoAV7cZsW50gb02Yr2U3KitHH
ZPreHgbtEWD+3C647g/apBSei2vwLxg8zl+M99WxB2aSV7bVN3kn0CID91oUF8XO
A9GKMp4m4cQvxzYGIgjXbOEYGpTdzxEP0WJhcLafnmnJ/QIXewmpgrrMVyp94v7r
U8vW6eZR4lIwFI6O9h86VjdTdy3DeDATstaE/49WT9Lb6jm30VZer6NgOgtOq0eV
iv5NF6dQHLZmVDZ7QNuJRKfrNA+sX8pJqMCoLtSoyY9OfZpU6k8rjWDDsrB8dRQy
1OXffFHTGFPDTRUYouPYd+7pQuVkmLU6N7W1a6F8L1Azie/8TWR8ZktQ3u3TbQc1
cGiUcg4DAVKDcU5Qj/+RYjpshOxNeeTUyl5S8UwikDCtgYFuUUGyfbjF0txBONup
n34F7/25THZDQj0hkcqmw4LboaMLyAl+YsgYAba+R+N4vuyls8UM3LHp7gzv1clF
9qAn4Tr68u2dhMLFXXv9tgBHEDuTcYs0ZHLFxVFh6mzamSvXSAzXHXL9d1QR6tRk
xb/4Va6dniEXpzfKN7NLfMBX+7olh6jo2PxpuoGM2/xXwpufndeoSaii3ZLswbhK
Aqb4tRxF4Sn1+ZR8wr/ACVf/eQxgxyGJREoZCPaaD3ERswPUwQcI71ZeCM9sAP0j
rypXuTCJRN+VqzP3JkreMn6Bvr8zfvBd5ob7HjXBpnBztn679oogMB+3zqsoE9LK
83PP0FOdLrEg5O/AWVnRoDFURFwCelvygfNwUEjtR9774lYIDUh5YnBVHj0SxK5Q
KguVSPJu9fOn0TpB4p7Ud9eCdVnDRCqokEhRd9g0M9foiuxKfwZnF+UsMBf6IpgB
j1a3I+Y5gfL8E1HKi2Hwzjs5frsKKzGGZxyd5KQ/a9QuaeuNUdWBs2cwUMIDDGn8
Dwh3TzMb8R7u0YjPxEBBdsVdG/qQKxBmrvY+NFJQ3NkSCZKC0fjvJPDTx8cOEyp8
vi4yOcYmzMDb7u6v6DTj3BB5jDxnraUCxewC0mBnkcIsyyXAR6HcvqwcmFObCs+0
R8EZDvVjUMMo6RvSG7nuEuE6AHQLFm7mO20AHyjJA612M9gt5rwZLADAUC8vF6d0
LwrnOxBovNVHdOVQt47TICzDjc9BgZ3nUKdPRjICQDb5Eer0/rbuVZzawp6ZuYdW
dG72eWNXyDTzgdBYFKfCOBqCS4Hjtn6hs0UKXDtkqtOAVuhxspWfZHguyVcyKwh/
s1bqGEAat49xR6xqAcIeFOWz+ABw26Ync1l8veTRYWZ3+5pIieaLnvoXRjKRoFvH
cKOfprxu5m62LN/W2GC6dfUdbiT4K1V8KxTiH6ubO8Smbj41R5NDeyj1149QcznK
CwDHTyt+z+3xHrOKDG2+59822EXzD6oZR8bC8eB+GshmPusoh8PTPwrS88n/BvvK
am/FScxSaLCBlVCJjBbu+RZK/ipLIjHnDq0nc7WcT9UfUMwaaqxoj/Y8hTg441ex
ppfR+s4vmnU7jf898+kXTnb77ySffvmxa9guVw/YtXQD67MzXZKiRKFsfPCfm/Jd
prXY+IjS4FN9RgSDytFusDhik3iM9czkx71iozwepNJUQnzgCt7GQfMSEAryhL6N
CflaPhlSVF3XOSyJoQHe0KoavcmY+PwVnqe8a7i7JPBzxOuUb2LZ3VbHZKXWqIlA
276LQ0JXRGWPWNCUfEsfUVJkVcgrQKdvbGuui7A9uqLzTmSwgxcTGUQQLwbtM1QM
p7ZIHwr4sbNrgjFNduwW2RDUp0nEejZgDFsye3SB7MsN/gi4VFzGwislSMYXZmhH
RKeavXkcCewUEwxIli6KbS3tCIRMr22Awj5hlc7wpFLru6RrBw3oi3VLjuChREuc
5Xzv4JsW2yLZDsE1cxz/+Bvaxon389XBOtPWVU5xvOyjRfnTqrAgPaIQkTZoFAUx
9WGYVlkcSfcyxYGEMc4gwjMT3fBU1bpuArpoHxWe79U6I/dhgKxohXNxQBTgkfHV
QbfkuCXa+7ftQcqZmWSh0W87crKwPirlg231Sr0+4vMgCk2nxVJSKH5NRb8U7s/q
6FVHcOp6OgzXyocqFGE2E8q+47XJJMAMpGAeveQQjFUoJSnt0AENyo01reVg6w4Q
yJfOOff66nqDIok3zNZWkpI8gc0/kRcjPlRjCmigSl2qfoeMllCDug3zgLiPn1hK
HoWBc1k2ZvsZaUrFiYp6T7ESongS7W0G07WNOd+uALWQKlTZDNlNRp6vm2ujIlni
lotfqJmRgml6lmXRPUyyZsrSHEJkYi6ivAun/BCsw8GN8CdikLScHS7gdwtpusA6
horzR5jAXrh70ZxhDYAjIBJzFlFJVZoTcDcrpOzzInJzF2HcRk5uNLghJTMPw5u/
vMdhEEmioZM+eZ2+gfIN3R2EMm4j9RSlUAKQk9DEUNNLYiHkLojRUOQt8VhmBbu7
09d6/SsIEbzbqldFMf4cqz6rMsF2XPW6jrZ82nlNXDM7buSoQRJD3mVNUJN5ozpd
j38hDfhK5P6JjiRmenUWvLrQLsti784WMKnPjDGMQIGdBdG3aCO3HNEbYF6A5QTw
S/mH5XIGqN3Xru1DgNYikLBFaRYWE0iD1MZcyLzKZ26awgKSBNn8zWK8NoYCu23a
qMPWSPBuqEnNnnFlLXfUDXgA4exOrxBTkpRRl3b/Cx/y6QUJ9zDDdBGKzZIkZ2if
DqmXkHc6pXtKZEiiiWSSBBOjAt57zO8wquNZ+/ydFlCqE3STm6caZORDL5IXIx/x
bP+avAwvAM7iA4fXv20SNCnkZZFAziYZlHgUiXtzVxxy66js6gk0D6nG7mRpqAAr
NZIFh0zsvxy9u962fBAgbOoJQoPnHzRXAVA4QGf1WwxGQkSTXvtKgOS0lYzaCtpP
VkCi55YUEkv5m4/3TJriAwc8RMo1Q8dcQP1YvgsJSHmsQB5g3tWtpgIBnDLX7xdv
OQyoJS9RtEP2rYgRfr+qY1IAvbjxQ9bSvkqxE+n31azEdLOWaLuHZeMxOGTzfLpD
B/a2YtvI1Z5BT3WOiqD1VT6fs/kpv0wohn2Zqnw5xmHBwPPHYcAkIPWN30+rOZmx
PYor/UagN9BDtwBfXqaHgY3BkZ1PHRnjFcRSSsM/wuMcAWCo2zQqhJ8wtARedfdC
k1BeiNHW3hMuqBvtMFL1dBTjIYNDaUBiHXjlGcEsrGz0BZ6VrRs8WJ/Zw21OpfbQ
rwUTDCLKGZls6rJpRSW1LCKa0iyqcqfRy9RBhTMxgAf9KSVBbRniFpQl8VrJCZeB
AczySv6eqIyw0Z1FRaEIn5+3+7k1tGH8Huybex96urjcYPxZOfdlAvxWFyz0YARF
ynURqxAhy7lRrsgHZqHN82F1lzg3hv0frUVN06NAjO8ViCza8Pq+pIuTxfWD797B
SCARDbF8fUiAg53eL04lMSvTaM++Rlr2lOc/6IAZkFj1U2VV5pQsFUrFyRM9ZtKh
2wMVexONU06uCrLobXMAdE4SHuxesuSCaoxe5lewP73lV4aG9UKjvzD0UvQ8vtGz
1c5K7fzQKLl6Wh9t+G5KdBI+HRf8AraKP1B+ntpGT5mH5vooLkr+hyE3ungkiMPq
VKko8a67NMjkhfnxQwITv2/hdEQLaRgVJjNaBMWiubODsUCeAhm8Rpwp4B5O75f3
N0GKTSotg5gh5pI1i0PMVuXKpYmmftbNBoX7Mwl2qxnRYWl63o6b+GDY5N0vtkI+
23sfxHkvukSnvCkVCbGzcHFTZ3eZon2be4hHS7bnrnbFpm/3DqdY2Id21GVqhKlP
h3B7bvcTyAA5eWCYhaYEjj7k5npnc3z1XlZjl/can+E+sjMPkh/Y6SG9ZBBPa7fP
xNDw8dkU4xB78eyQRE8NUKCKv4v8u3RHAXjnB9bJxsw3SUBgYdH5S4cwVKHGzMG5
uCxGUYVemf+oN5fal/yMrNtuw2fLg1NLCUhLfQNcHbowwcySPOiTueWT33HTTDKc
qZEZgUo/AWYyFqn1arvTlcJkzHxEeqqAFAGTuAx8CNDDY85fIFDGdHUtltoskJz2
aHT2odLzvF8O3wpxuM8L9XD6WihCzxbX40PXf2Wx+QYugk1cjzDSBPH0HJv3RMBh
sznOQeWCmDCJWj1v6n+WyFprAQ1tLLJtwyimnSmSIsXf91APY9kDgAULbJbBmMTN
jhSzxOOuDkXgwhqcgNlnalLUkHTu2f/bLNGuhGSBpQWleVVsb4iJ4+Gh3GuAKaCY
+wUG29/DlSbvsLLo0fPnd/yYYR0nHoZ+NMfbCGrT2XssVtBUOE7v8CcJn7XY3/CA
Hr5r1tJuRykJvoIr8I8ltUp/lUMGoORGeEPjSguXN8TZQj8OkR8XgsBkxBRCr6i2
Ujri5HOao6XwM1qcUQtovCniuV0EJi5S4ur7McxPRaABN/ioZJdn2ARfVTpwwCKx
BfRBHpOgqB5Vlp0DU3C3qp9gTo89OAK7TlDHd3iX8NBu0APLoi4asMKWLpPG98NR
xQyrUh8yP+B0FiP1roOZm4+v1v+SKUw3guwtBCIksRJ30YB9E8ObxtxLn1Z8Tve5
8kYJDQ2crZwesokAhAvrbX1a5PfARK4zdEQu7cba7G1xSOZrrrlU+zNIigPg8/UJ
NZG7IzLis+cmiaEinw1Iz/LIcSmSLooAzom5PeZvlx/i9eIBvV9ZHl6uBp4t7obJ
mCvf+SVA+uJUbS4CEko5oLcbpz4qz4vt6d1CpFpGcxt9Jdhko9ZOa8RnJOs7Cj+m
jHntC62KdUj5hWqS0cmESqrz8sDTJf3++bNw4tdsdUGbGg7fh0j0HAzMDqkNz8SH
hG/GUAH3+WNMqdJhckdyBsxHjfkhSDHQ1/xd0G+0RIEI7fQRlr3GsGOZNmRutXPq
Uy69p127hO3hq1wOsQ+Ja0+7Yu0hSLEPAohZRaGWjnVPnRR25IvDtDM4jtb56x34
MBzgd0xILIJRBKZ8M2+0Nruy/I7a49Hev/ApjqxLkFwdeF59LzU43YyQ04jKe55T
Bj/O6O0L9kJI7fSew19XDHMySpdObMCN4EFxq2MZqjovGY/mYzAYPEqVHuoQhKgw
IbctK/pqFKdub0OikNAKO6c1K7ttwgQndU4SGXrcQdDbKYxEGA5ghKukHZGtiHLN
nRlGEsDvT3C6YAOOjUfZU4cqpKJIajAd6Oq5KUuYreX+tgSUVe8qLRhmGCnf9TdV
DPnNvXsdY+n9EBWMHa4IHCI+iJRIxE/ohua+c9xxuNHUBcFVEKspZPmeK/F5yHEB
vA4yaxmV6TunwnQM2zwMe+mQ02b20cZmLBkmRo6+7jqRYvjAsR0Denny611GNl4z
u/9SeSVRDvJa5lKGvREgi8pwICYBg4dst46zszs0dnkTFBuSXw0DdnLlJFsbF+Hi
648amO+YC3VripRq1U07rP9cIKCdHDqKz2wddrGxV+KhegZkOSd0LCLxn3qJPVwp
+MFeMUfqbGjhi1BKHwNub3InZmCxy7rvRyp5T1AapJLOxfklTWnAxeQS/wYcZ25d
Ul2b4dq5MatAqVWY2CENvq3ZUD3/9Ies6c7XEySmQxf0fWsWRetmw8MFnLgtryTT
pvdIZs1bIeto//dGqn00cgfXpZ0ut62wrfknNWKKHF+63+r73AGH12gjZ+VigkCj
XnWN9HBqszMak6XNg8ezMp+kzZ5tRtp5e5xsNVt9BoRv7JaawxFKy7AZno/VSDFV
kthDk18Q8F6yplrgp7SQB3uEHuQ/GsiD0TcSfxdidS4ZVC7qiWrELVgErtwL4kVm
hzNkGmaKkGxcH7PpOpCGmAyu2Kfp9pjf/WyRSvH66KH5ZcrR4o2fEMDXEW300jK9
BjlttE1BfkI1Yr/mkezSuShA37PvMHzi0XrPERwnWuckCLaOjuf62utz6BdO9AMh
LLALzYuyAU1Ju8WV5z+Ye2YnRtz5B+C1K0887vFdQQfs/vK+OsaW45vqm8xlWsmF
0y7NiNbgK3g0n4XoD2lmRvENMRpkUH2QaanapCNODYJIJNzZ0zoxX/u3NFpkl6Tj
6AC/5I1+nrKr1KFOWyy4sUTSZOrYIp0lb+Sk9rsN0lfFxGmYfuynFSnqvCC2msqz
ATURkcTKd7hv18nDT4z12POtJmHfs4Egh9lzlVeM9w5pCbZac7eWSdzhOgJto4cv
qs58cK9fP+jxtnxwYdUIWQeCfXTA4Fosjfc3S2xGDzUJOOs0AcpHZ/EgVIZbVczV
EYWGjAVtU2shBbZS464o2vPByx2H4kK/RcXdgTsq45IkXHgKOIWdKRWF7tFgbS6Y
vH8ddjbfaEIEzmebe9Y/PcKohSDOfY5Po4Zpq+7VsUvSYs2GAk8ivDOOu8cV6zbO
o/A1JYkC3J6Jx93azAkuREJwRxfSleLTMn8XJdA4U19mz4/0Nubunzf6pyZc7c1+
4sGGZh2+WkWH46d21PKo7MbsRcEN3JChfB4MWskqMq/aA2yu53Ck4ItQ9Ql7mOaG
8aAk/Olwkso1RIi123zcJZ4ynHD+ud4qiKMwl72tm16GDnXlahko417Yk8I4wWNC
88qVknM4zjju+tvZI4Ot9kJmurRZ1VjAh+a+jCUU0ymZcrP37OLt4bjFX0CKr2GH
uhPj0+7eDiALEsYpdfvVZneBCVkuja6UG2LsbuTb//Y/BCbkQEL1ZE11et3vi82L
XIS0y0rySkis8RaQQlnftQFs1ZwkxniRDvDMrLHVCaiJvI07JXe4LXF8kre/BsTU
poM9lIfOouqm3m/GLH11LASHbT2BQ0MoluXQNmMVcvvV1H1FzBWcMtFpC/Mm7Oh4
SJ5cHQ5sWhZPA+nEvuOxjqIhtwk0VlKl13yhTUWXfBbCHoEb0ARdoTYTQpbrX4Wl
2LeIi25LPEjVw2XllIkTP0Y57BP001kZR8RFo3QpwwWwl/3qrkQYuxaHEGWvW4mE
Eo52fKInKGp8KH2od5gnqatqYikM7tcI2S6Y4zHjaFuQmABloqe1TW1OjMxwHmHl
CNzdi2/nJjRp3aaSahspFgG6nJt+GSASI6q2+NW/KSWnygWBNbg7tWAXv+LP803n
nuIAYCXKcICrM1ReoB3pUD8DLEMjUHYtJ5ev1qCDQMTX0VcQAEXjsuTB3c+c4P5B
t9en7+EgcMHJVeEYYqN3b9bp+vDGT+u+sVd7gIw159S8MT/SqibtpYisTcCrTyw5
tyNbFQr8dkTlUvNUO5trxE5Il8MzffeYtMw2Bh3aWx6BAU0znxD6S+bRF1omw+Ew
TO7KCUjXA5EM4IaCYbRmDTNk+HT+JdFpps2NM1gVwa66sifgz7mkGWszZsrr9+jA
UwjAbIvMeOC0N02TAFF4kDUhV1JafC69ICyRk4BU0Wy6ngi2Liy+ttJfSs7pPebU
tmhGTGClduCFJ5rmPcE1Qo67YbnLHBbneryi4XpR1MiBauC/w2QL5SYJ27MswRbU
k3HlBH+6GvYSzJlRCU8L/9A68kAYfVhKTxelzIPh4C3fwvIZmbI9ypOQ6mVsVBls
qJtBi1tNoO9EuqfPAsAxM3T160Ys4E6R9qL7iq0pMOC4l0uWiOWzwoYZdsuX43+e
rp6Q+1keP0uWANVWzREJUtRhhvqSWZPbwl9BkH1OlAvovDvsiG0HVyeqiGknpV/M
KjI7XZYp3X7OIoHl5Ojb/hyyjuZhjwPkc+eIueVpbv7HqTVQcdzxVTe9fCTkPVXJ
yMnrD2oEpW+UvTGSpJo1Z5yYII0RzrE1Tz2De1UFHpPuyBDQ65VSTn8UOh60A1vj
hr1M5wM5FJ7WYcSfUBiwDgIRC5Tqb43/Jb1Ii68d+3JeF2LZK6D4/C6dEki9/Y1D
GI6rgBYNy8D8W7OBU7avPUvFwrs6rJNCHHKRZOlARP3t4xvXBwOPjc4AQ1l8WPO6
ztly27PlwTZ/eeFlgqyr01iFdF9NT1AKsWNv5tDn7vYwxdGThT3PkcALSN/6vDjA
Me9hXpJSICWg8Xn02ubUB+QZCuSwjoNzN0dzz/bBcfr9N2VVxu51Mxiq3Ouq7Ju7
SHdQLGjftq48ZaW9U9dVd5Dvm8iSMnNsFCrOGgVNHNDmU5U47VMFJBZlGSaI8n5/
I2Iqnus6+uGkTLwguyRPCRuJ8pARCLQlxDJLTogavl8y8y9dOzyG5j8FNBUp6buB
+yMriqr8tyaWm08/Qju+GHg7No++2KCdE+kiWAYrNcGpGSWvXQ5WAso11PH/ohLU
eBiw20j7SnlIv9+hk5Gi/tGgpTTv3zyfgG3p8bumlMbL7O9Al8bT9S+XXIC7a7/7
nsqXc+1Jr/EFwj+SOQG7szmPFaulpvQ7Xmd7U7brlT3da7beZHmp6fj7Mx/EaDCT
WwCnVnqcGpplboC7tD6LwBLLOETqq2nSAxYr5YS1GxM+GIlnVwt/h61vpGM7Orz8
ilNAuerQzmSRcOdfZjqi70CG6CLr7Keq1CHnXKPUdav6EZ1jq2BFer4b21PIRLmq
6GdbEkjF8DWlvDaNamZ6dlEVhtfGiGgjA9VpY4FkHAwSkYGMcycWvoq+2rhdK/l5
5Gl6M711J7AWCcPwwvmSiBo6VZKSirxF+rqU4HdYN0rA0jhvk5EMlL/OtTvbf4CO
fdmlPlU9uxfzDEdHzw+IOG/Q9hFmnXJG5kC1RWKNdzDJJqEfyzpkhQbKTYUIYeT0
2dLxO9KAQ4s596wg5LwY41gMJL+RGFwWwzqOuG6DLV36/HwmC29gAkrZPssBfsvJ
IAXqohrKmb+5OpPT+KRtYraj5ERFF51sgrd4ieVsN7oAgTZsQhpu9MBiLXQu2aqv
pMa8Dg0htGSQit8y2I6iKh4lbuL4mujynB0kT39e+P+2d+JTU3Ue1anuLnYdbVQP
F9dHNsZm+0FUQpD4OKfWc9j8FTGXteKwslMCpMVQv3kohczi8bBChEbwpGDwdZZ/
HXStEOkwWvcxLmCEmDQ30aHRzAOlgzHBfIRgcUl18j2oNmbSP7RInrH1RjXzLSdz
SQ3Ns1kqb8jIkeptipm3EUPFVoWSlc42pB4x3y9R5WL5kjTf/TVqQWqpwKZV0DDI
6KFfbJPjeX6MrTfszL4UdktenOMOMrxc2B6NIWyvmjzN/c31+Xn/MKTRx/OKow02
/iORVeXuxHKh+bN3xtRa942RnyIKsp5FvUVQzVp8Un89SoCuA7TJm/1/2Av21/ye
Ha1FeEfsirnHb6XEMJeWJm0W50CnT17u38UrVsZyXq+COOyDLu7ztPp4cyAfkdKo
OthHP3WY8F/U/2V0l9XDM3nUFF1LwaenC7P6O5QRhv6rCu6lbe8fKAH5vYdtePdJ
mkzPltX3ZoASD8wc6X65S6z97+GI57eiLyQHhfeZ32MchvNK6a6C+bWqe2dI3x7b
xvRdVar9w/GwPmhraLudqqjjyG26sLfZ/HKnxVyt/bk5UgfyyxHM1MGCQPLNSpMv
y67+YxNXDHL4dENN7nKVBc79FV37hg6vtQY89OzJF2M6z/0gBCTHxAUyqll/yFlU
djE+Bqi5Em5MZ5Roh+fn6i9JTZjou+HbW8G1LW8GgBP/aFDO1Ytj5kqh+/l1D3Db
Q7OO4Ch2G+E0p9mBJx02ZFQmfSEkbiJzeGmu7sgft9thA2Z4C8rVy8Jd0VlWFd2Z
lTIzuFkGMmCAoKxDTAwmnglvyVP/N8UCm1bG0XrK+4cd7ViRZezSISAcrPDmcN6L
6F7pu6q+9aCaxUvIdwgPK2VuwYdVT92m/wHRe12F5n0jie+qWxGPsDEgzRd2ZGGr
WVxGxBKWKZu86huAPUx80QsySeHRsfz2M3AV+Ntp0oDKgWW0qCYRFm4YYNuyOHLD
1OZ/SlwcH3ZGIi4wgSuhcIGhWl4snKHpGayvdiLdU5k5uR3DjNM7PuD5CSotrhYP
BzQ3DI56Bk02W+dCvdSIMIMWq0RhUCcrPgvFJUaOAIM4jlsvuBbrU1tLwxaXGC6g
k3WAqyR/TeS9MuKrySAK3h+uhZbHJzvnqGBYCipw6pqRPJWpJeha8DUdVCZEWjw+
Ios3rB+4W5Xu4fZCIVn6y3ewncA5n41LF/VllBIgRmNsZbC/GH8iJfWxW78VRoZz
fyjD0xj4RhkF/LZ6wrkFYUac3VMiwrZJ3r92h/WWUzgy2pgP9msckdQkHltKNvBc
CVEWAnPPEvMuRoJgR43/a8PuHfc14GPvEz+tjy2oBlSSZnfsYKV4jjqvcE6xbVNn
CXqFHnxDN0UZOiE2Cfh7Y8wgVR6tqBxXvuEHY3RbVPbhURH06cisPw7Pbgdr5YA8
KxSErsBURWqYWc9BtdX5+dK0i+4aWdSKmlcB8+2vNsAdu71UYrKwxbojj59ZaeLy
c3CGGeTAcTksyWDJQI4BtbU+q0jxmWE3YCQQEEEHUHklR4LsrVshd5tRwghKJeAB
2ScGvzcpMAnOdxdVNTFxalUJMQwif4jOPHJREX/RFjbGFR5bZ8NOqgq0r27XVUJI
M+cPiMIp8OiGioE+aKdQEy510vN9MSioLtrmcjnEJ2W9yRn1Pen+9u+9WZ8yONfq
/Kvn6uD1gRI+7PQNImdmilGN+WnBYqB/q0IxZkgLL3sfdkmBJJvwWhpO9FxU1pdu
QsEktIYEC5sp1rI+PS1FtCdOZ0wHx+c/78eag61aS8pxeyAtTHGJEDINhm6XNmnb
9PcISyK2cz3pYlfGZVVawRZ/QoEmN9tBAMI29AeBa2dDs016fiGZf3Gsidwh7wrg
NuCJXXpwPz5qXlBZZzSLKxpE9o8gZYuoyTVm66xw9n4BUS+DSiWbTX3tTgry86YF
GA3ya1pnVFZoY0NodSp/64P5DV60G2N4fze4Svj3LkxQxK4TMlu4Jve7HKpvVcrd
Mvi5LpI6j9TqmjRf3IGNtcLwhKaLQ24UI6QvYKyVlHpEvwjZReSFExWFbdo7BDlH
Y0GCyUSG2djYqbub2DP6JY8EbUVVHweM2/7154Gc8ANzdMSxRc3f3mc3gLfNr50t
nt1GfIiW7ry3ECyYED7TjN/OcApsrIaGA6YB4j1r15ZikoTe/0VO2iH/kkmM55Q1
Is7U9+oCQdcXlyGm+PPnJV20NRw0YdfErV+NOMEw6nU/8ZgAUBnu0dJd3w6pVv+R
fPDZ7WEzeKIJ/TsDzrWUQ5SD8GBrRQOuLbQKn8uyGy06wNvXIIZNbiyLuf4HBsdo
ku2O8VTfV4ea89QmJLxWUX9DmHH5dWLcbJXW6ow5/rbd1a0OvtD0U4Tx1n64lJZN
ch3gw0etF6UZNCaKQBHqszxL+Mg/ynjIdOyZvvTPelY8zEgs8LwGKImNSskcrcMY
ybXcOxAd6fefvGNHDfpVe7nj9zpMSApxHTGLPM1ugv2PPok90IA54ZBovSPcJh1h
kN2azJaflTaVIdcY99/8LanaLP+zeNh9/HXqUpAXTrlcb297tJ86plppFR1SqLgk
D9PS6ru/ni/RshAmvSDTdEYCNYF0yQBCisN6CBmj5uKwdUuOiAG/Nr1jzwwNVHOp
NjOJqji/9lQZPhDzODlZ8BK+eo4ZqFDS3MJ6B35VaWtTqKs5vIVa/p9V1pxrmnDE
sRguSVtabTqPG7dYfTcKdIYS150q/FcwzD1rlwseQq9PvRhZHM7cmCSGuPlNNPw1
E7Q8Upx/Y/kJmqLuG8J0t36bhngu+cV4C9ZDxpsR6iby0Xv1AJq1wMnAlxZfYSOb
q4n5sIIgdnda2WJoz/jk5CxruHpcp/gwzvQkkUPTpxpNir/LgYiwWIws4K1MANvh
mtTWh1ChozAp+bJOKA1sXywjG6vMjM+4nEU0cP5wg8qyjB5hXn1BzcFmbZ/C8aMG
FZRUu+MgjkbpaAftymno9kMt2PSIThmiRSGasmEiTfb1qA5y/e1gB84761aEMHJM
3LwlTe1zMMy17ibHbPExv07fayrbzoGP+O1d48YuzOEg5fSICeD1LNRmyMierYeP
2bsBna8MwHwNA8+NNTfLFO17Y2HvOvEZeEEBs7/QuDlmIQXlpHzEJ8cjKCwNneCt
QNQqjc8dDqiJeffWliwhXyAmA/+hFiq6y3h2popT0iLcouz2vg/mSRAZVOEWa4Dr
9E9xQINGZs9xyAsMG8UpVI69Zww0rYNNWaG2vh0fBNC/rRwmvHzorSLqiIm9JrXP
+mFzmL+VUCGwBSMuLTuoaF/C/JONCnXQWG4wv2X/QihIhQdQWm7eJvxS8B12MwyE
FrkG4imO5y080EBqGvio+6n/gd+V5tggyG2MJwatQAnFpE20h/rNmvCp8u3BRdiq
fuQXl217a5Lw6EIcrvXOv6VmtYmNMg1nkrcNciXcHhUDPejLQ9cZ0oksop3Xl64X
dU9AFZ75CDvxmDkB4p+ahdyZMgELwTHRXmjqZ7+FklENy086bCGuZ+xHYDkJVvG7
WB0mV8dD7Lz3r1UghZeHYuXok97Fcxf+5j7qRaiQbFC6fiMd4JGi2A7U6B1scLPW
V7cODbyHiweIyO4jjxVLwnBC0bjiRkE+RbF/GnimRepCcGeU8kgho0FlQQLOh81C
EcgYnascb4lU8j5YkpfqZftgPeyA2D9IVs8uGz7Cz6Nu2d3xyb4JuGEXhz6uTPQ0
j88GEMPd+xKhPBEJJl6QOKej0jZEqsSl8MNz0ORVv3uvOVZ1+CiC85HPtYE+kV8r
XiD+2ZFR2aPoqp5v++QGuF1NvjE8sL0kSoPhgiaWA6YvkjB6CkyklN6CJ6H4fUTy
KeBhkrOj3WCxz8yKf8uWw20JaoCRHQXFIu6iCdeKg18MF9s68Iz9tDLfPOT+SmcF
uQhrUQoG6NUV1+yErSLarAjoLdS2I2pVMWWnfhsrMD33lA8HCF+mhNF0ZfFiBf5t
vRG0QmNuz6ZYpzkmzsdcb6nRvm4Ur87zpp/8ht/9PbEgMUThjMdGtyZ5ErZGZTvL
qLwfS27eQtGI6cEIQasz+9SxlHum8KXEfUsvFfvBIWHxXpZn9vlib9ArIFl1fKJc
k9ha/e8a7riKif6O2qpuDjngq3i4+dHk/67SlMPKHiyHSPxmCpPUSvOqH8Ycbpa0
gGYkE0IJat2sx5ocApwRROuzk2+7cgQGrPqTz138eeaWXlUzV4xvjo/oXBeYpZEA
QR0GY+2Xky23VkHmmgUauGfeiGqjj3z7v7nVIjPDfCVi8H4Rw9MBAWziMz/e8DN8
y5CP96IUphhbrA0qTztBrJmpCtNb0lXwTvibiTrUoaQDP+oEbLYTJ3mxLcaBsVb1
DoteeazlmQmo8GrLEsETtxlMR7CGFtdKWA3ApOVfS0qqpP5dqup/wnXnxC1pZ9ci
M94Sb8x/n0+zaiYASSGOY2ongYpSwVXAjVfyKSlZXT+hCskH9AmKYuUtIFLzoSDE
VM6sHB9QwSU6D18HBDtOAjsaYZA9d1rAi/Jtswh9Zd2NhowYI7UARY67ufWwWR4G
cXIfIDiX49FgFiugpfc5OQu9dVXjAFu4Syu6oO7VyS1ubJJUD45XSfBxZ0RmEj8h
gTurcaocIeTZGBSllOWcVhxvddBu1CQS9N2rcQI4nGRrqZZD2P6X6CN8+QWRYKkf
k4HDHfTS/ouMYHfE+SMohr1bThKh99HqFuTSBEg2ovdV2BFz5CN4EIFohAsGOpWd
K6ecqjVvJvn8Uym9gpRpe5GsYU0YA1VRznI2+jVrhE/fTav2HRexvJiOe7wWUC5R
hqYrMoxw/AQv7w2UoKQA+ZzOzXSY6wPD3CRu44WmRENnG6LvUhNQ/1UFGp/R2U+2
slKUvSDZXOHEtxNPORigcJDee5yjoqZ1tb8uCmYD89Stos/LdP7iwn3DImuNxxQ3
vX/lPyqd4hlaOgKSX4tNZsjtfdaUY+DNmGUt9Vtod3U5imVxSLWSQQxdae+MUb7l
AtXTNseAW3ZWwlV33MZjecCOGSvPt+EiUSarPN/PUDTNvGqT4nDtbR78oRhywRqT
eDmpi6P7Vd6KgUjxD2htSaBczUkblSo2DhLJsI5s1YkTPiaQdtX4aL6q6QtMnIfw
8QYSDaqcAKWm+CaftJk4l1resy5Vho114XtX5dT96QvVvLRrpRPXg7KUFV85mbFD
h0osDmykm8OK5LjDvSATu2YbTV7HosZ1XTHiaqBRX2jCCs/1OqAple7B2RkSyqT9
6dqp6ZJoxUotC1qqHifELLm9Pd589Ffa7QEbOZYkKvcQTNEFDonhEhTz7nM7/Vtd
9zyWZoQ+leUb7N6k0gfGzzhjTKuf/C2mJlFEtQMZKd2Nr2G99Da7SJEMTZKGEyPX
SVC8/xzefYsps56nm4kHC6QzqgxLBrs/hHlhyCoW4Mez5ZRW917Zom3IpqDA6aLN
Ia17ZOtb89u2dwnR5tu0KQBkNVy8suZ6sYxjMFnhj6yuO8m+IOJv/Rlu6b/TF9MF
qUKweAUWBfde7h9MVWpg+h/oHzwHA06TTCgvgtkhaidYP0ejyIkg/wS6cPpSP/yp
PZAl+C53bm6FHeMTAT8upRz/k7IQUfBsWuEAWxvEoyU/MQqJ3gtpU7j3zKJgUfo0
5RHoanSkChDTUiDwTlo5FUhLW3K4UdvLyayfQi4klDhSc2cL43GDBDPgv111cDc0
CJjY3kFK+rVbZLiHY+bPTbpCm6u7GUdDLcFpoetgGvafDK+Bw332Q5/lazmTnKvr
CFi+nXwd1PRnRPjlIDYqbgtHoaQ9UQz3HlVgSLGRsLBKk+nqZyJmOSvhswj5unHG
AAx5sERwYiCtae0uhTwt4kSSa5ry4+8QbBsflly7pZbVEMaN1De3W4PheEdxEiOh
rvfnGxG8ADMBswHSHTo2GGLn4dNTQTlvseUYE0P1Y/AViA8opRe6vs+f6UfF1w1c
3G/hTKO05HPcgECgKp5q5LNwLV7QlOHNTlEplDHFAaV0uAcrBDUg6ewEuYjR/AOB
SEFPw2SqlG72/9XVKlp8zOGWE0dj3kQ/p6qJZN8IEFyMety21LlATcSccQVGrcvA
en6u+KdqeQCkmrQazRlx4l/aFjt6CbTuS568cM6QLU5N13C5PCHxQ1cyLGQycuRo
WDolUHsbgt0fM05w2a8Y2Wme1CT5FN45b1I+GRZPyVGNyjm26JlKlAkwSeiTzfES
i1nyfBwJLw2oZfh/Tw3/Xch2fh/dOz5cJh1NRBNpv6y5e1iTN7f7vueseLvRayKC
L6ott5yKw+G/Puef8QwKUzTF/8x9mFFP9cauv9pX4yaagxZX59G4YIPZ/PfAvUQ6
HeYC9GDUfxafdXHdQBhYO3/11QzKQafInf8jE8h96qbtdjBRcMVHy9kIPSZ4JudH
O72m8YZXdrMxoGXCiRR5m2zHLuXqLnb6Xb1fxIW8TRhPggfpiE1Uid3lOCo8q9Iq
YMa2vdY8nwIpZfxPWzilNglL83aDdxKRxERHbql8T+rxqnIksKa00ZZOVAK7Wnm6
gsf+livQd4kItARdmA4DL61+GGbdY3mZqhpgl+HMwW/2lfgnrSjerFDVoBrunrm1
A8mgCZDFdB0tO1Dy4VsHYY92i1yS3KgYrLJwW+acn9dNLQgFnAqZOzNZnczq5/OU
s5u+wsytm3p2rjGsrappNlICINB2b0tet83L6x3SKErW7pqkWMKvrq6/11sxsA2K
aIQCGyvfnUu3h/Em6Po0rKaxrrgklbXZ/ZTeQWS7Nm74ZptIXdERfFZg1VRORfGd
maIZ22x95N8tvstjmqeyvfH72U1VxhL9F1jC9ckJxDzFxG9etYljz+YQp9SwjQTk
jb+BxiTlGuA/nRCAIjBBEYfxEHdu88QDQl/2y4mLXlE1zjnqfpcYY0NoSccEO9MX
5MYNeOo1/mPXdxPMBHDCjD2Zf120zsc2PANQxEJ/jso4DWYl+iVqCcD2XsU53uX8
SW5niNtUpL1bX1N57ANfFQXfvcmvX8b7OwuMyBGk3LOnKH+qhthLJ8/t6qt9AZvk
2kaviMaakAhKBOtTgskfasooH0GkOT4o5LsKgPcsG6Nfl0osAWmznsImwe/j+Zgl
VJXKDiIPGbtRBSdUlowQ1PO5IxWFFQMuPP91YBv6+P1/4b5YGZmKIrfEYtxKxzRb
QVu2OjsXMUn965xIPTiroqsihYEnYhoWjTWKdCEvwVd2JmyIQzabyi2TajB0BtIn
617wqPuRV5aU3ERgnk20Vkduv1RtNSkjxj4gA82xCvHdhNVLxSfnctVQeGnSQ5g2
ETWJvoSnAdDQL9BaWugvaFlLhQWeZz8coODa+dYyGzaAlRmYQe7GR+An9VYOupeu
QIpSRoyCZb4rDwF+XJVQey4uymCoYfxEkds+6jFSPNQMV8mZPSbD5hYt/Tppr7iW
joGXm1xSSaHXwIrdStmpPSf5zBbDnSAk5OAE52dF4IRtvCV4Fpaz6r3p0wlu6kbW
xgqTmX0syRNz97/f8UiBKqCUMccBkZ6dl66B+T0jdKYlVtd0D24fqPYsgveCYnBM
sHx9f9VuvfZDHcQrbHNJn13FgRUXFmtL8Cyp/3jeaEM1L0lF5I51k4xi/2ug4DGI
0JzESq04+s9aGMMByWhHlzUv9SlVfLI956HJKdJ5+feO4E8riu+NkemnHTNpgvXq
nLFNjapbIbgh9HUB/gs8WG3Uk37feSx7nKJ6uZK3r9+MVVGmJJIwacBxpRYyShRt
UIydvvROowc3oowdPGS74/1FuALj0BPWKV7UjSfEG5w2Gx5ah2/HKQK7AHFw59LJ
iZcD33L2gy/6F3q1JMFKCZF8gS6/JZs8i2dcACgR+Rs4k042LVJ6MaIH80n60SqB
Dd90DNyAWb0hoAp9ZN8ZdmhIfao/I3PdXY6RpziWZDYvUFLW35FwyF+ncCl7NSgw
4NGhE2Qw4+jOKqpy/LU8lNgK06tTk5bYIVNm9EMabnKfeAWAHIijvHj+j21+pi+X
jEdHTKtWQ8th3G6rUprFhLMxz4zsUH/PKGn8PqgiJUNCSgBftzXl8x7hiWwYYpBg
QBZQ+I2QuR4CefaYdiA37STD6t6ZyxYqw+snVAlY6ZXmr8eO1Umpwf+Zt7YoSGDR
HlufErgN9peWMs8YDLS/gi9MvS/pn0AdvBnG/zVIr8pB0eYGN+pUk0jXKW2e+bPC
SDfz3yVNJ91uNVToO6Yr61XeZgCQJ07uCmixRn1zXKp3t0HnpBq6wtZpObyd9UsG
AUIkmdbox31UYOYdwH907od9Bs4ay0zfTKaV1NV8hYYKiSM7s5zuZxOH2gRtPBUc
ElrUBh9BApVpjyiRKDjKGk1+bIGuHRj+i57ocM+T0e42PRarl8QlMalyta7oiPK/
732L09x+vOKQ2Lpl4m2pbObOlI8iXgFvsh257y9JSAN+UGD6WTVc2qC1jXhIjhph
C4CBjfrmFNeVPW0317bX70eseYw3iC7DW3NbiJW07iHoETnnBsATR2WnE48LBkp4
nzVaPCTzvTW5Z+NuFL4XJGLpWc52G4+IU0T+kenSaac6h7zk1dA9mACj5yJeagLz
rzR6Yb30+O47ttNqiSCse8YSy9rZ1J/m34+lLwts7vXlrvBjOPssk9bvBFNDqIAL
X5lwiF09J9vsXvPbl6W6sBfG0Wmgj2h1baeAuYVp0hcsW+oPXGfRrcVAm9d7Jc6H
6P3j4MuS/63VTCyWHP9amAzTmII48PA0PWQrY0IZsePfsv90+mUUsMkw+iGgOPHu
yyRSe3o0Mfa4car3UPH5iwAmyVnTBFhA7Mr2Y6NJRwCQWONJP9dUjiRvatHo7HkL
HntpWtgokPq+MUXRgLaG/IEPUDHkOxTeub8SCr+KHAU+p5WHJht31oLgixEC4wg4
QMF31PTYYw8dy7Q0bkZaHI2wax38KZ98LmXBuuGRUzlVrhPy70jyN1rAuks7vAtW
+/H2Q5IWX49AGuFeDONkN6nDmgXExzQXYrXHJf0+3EEwDIKCErtM1bvMclhqKwR9
M6rKtgwI9p47d+gO2gzPhUYhEfZVzf8Fzwx6qi8kZBQfrFKKWZNFCLcx9PjzvnzW
o6LWsDDCMTEOECIcQA1jEp7e+/429EQJ0vW9HMdJMifdvvp+2w1KlH0koJEzjf86
nAPwYWNxw7+k2pL2N5uIejsNxM+c4tlp66CP0myC94rGLPxJ1Ws4IhfqzjjHrMcL
eBHW8PvHDq7kUQ/3qjeoLA7Qjr4ENLIWpTZlfWi02JVivAkcbJRzqZJFDdCnWcWE
5Rcmna0JYYt4apgmPIipCsBkhmr+zl9bfPDm+rXDfKjn0aj95lEJffAVr7IvpSrr
rLt/SlE9DUfM+lhDIvxCcF8Je9azu26TLKxaKufr0UXw++QytSKC3rL/rd63SvIj
KOOGov7twIUtL45MrCV9+Cn1ZvmGaiEMDJjrs8oFuMMIseAIWSHlB34+m51XDm8C
03MhyIkOKi3d2H7rgCcPYpn9D+1Y5TYoS5ffGnfgS5XL45WKJbwdqdDkSAugh+BN
eFOmk1Pd8NyX94z6TRSXELk5LSQ2vlXodvOGsIqrBN8CeWYXGctl7QVHnSJBE0IU
jIstCRzY23YArpeJ634lZk/yg70mjbMz34byImJB2vfuFsQuSTdO9TZMyEj+/7ty
ztPFaVDcXMUSt1Z9po76gWeWvRYQpfPnThJ4ENiYdXcAP1pl2fcrCFsqDbQ1PuW+
R44It9RkLJIfL7aQxlk8+jdPPnyKtLhSqTwYkVDJ1LtCg6tAad5b357jVrswKTtE
qwkmtI8N29KAlB35svwqStttaRi5Zh7X1h+xUR+yJ3mrLnBGnPe0lI5r5s62V4Om
hXTO2erBMCn9fizanKckJmBvmM7z7SV6SI0hkVjJo3fvRWAMzFwt/3HYv3RlwFrV
A5JvWP/yJqrP2xw5nXLUfC4xHRL7SDzLiki4bWBdjUQd87JEylCGMGzZ52A5Bz0X
4T9c2xTtWY82qhOHfV5hn6+fRfDH18bUGwX7eZ27HxXXP5/NYhsV8t3ParqFjdBX
QjIPSAHcHLYRjooYhR+WNq2R9Lg24JvjSvCcj1jB6417mao3xcHmUQKayZBOgPnm
Vy0C46dCMNoPvQMjYAKqMaGrpoQ0F2OfkdeaUqTDBQiz8Uw3Xw0OJBVxkLuInIR0
QcVOJabSPQTsQzjlnR5SaDk/7tE9csQruSmas7cJgqTTQPz1P0+CW1+tM5w3MIJ0
7tn83vs40iC9YOCmBKNjy50YmuTB1ACH1ilRIDwkGUvgrc0DgByJWZlcIZ1IUgOS
Pld1Xy96wPYcMqOTANCxDzewTOONG6SBINh3YydmHDviQc0tJYeEvafNAiwsq5Fd
bLr2RwvHwL0+ZgNjqF0fHwUaafseDPKSaaRc7kjewThLYb8YUzZZrexBsDwB3tvv
jv7qP8bqLnz9SkJPqShhcJn19cL4N+KWtLjCZijTBRtmFGY/zC1LsPoUebe5oTw7
ofOKL+1x7NkaM0qm5nxfi20stHRHgLKty/pNSDJGUtaLPckzqdQlServGTqBoc1K
c9GENcKJvdCPJjqTCU7nq7lPhnRMX9YdpysNDplhIzHJzNslHna4yhiIYKJYKqAM
dUG93Dp60kNU0LOmirNzhqDnpnA/3IoYYyGS4kiYjmRCAG6AHddo8iuSZcXia7gx
RcpWBv1x5I2TsEPklTRlKJDPoeLbxbpT1k7brQlUw3NLuH9FP5WYkXDVSfLxDqnw
MqEoFW4GuD00GQmv5sS7BOj/OayhGNH4N0O2fJ/Xm3Ts9Xv1zG+p56Ea/PidHiq5
9oUlzJSVBIXFCBrY3H7rKX/GBvUpLrW392pB4G/2OQNAw5V6jZJxbscNvcMVzGzE
bGVzyIp2cxyVREw4OwCaDwdxAg4VVMpqoKIww69H37tfzzAdbndmri8B6Vc5tij6
zzN0jxQEDDpKTEsUaFJcOJjSPjKaRGtvQ1bfVuGWWk1MhFeNxQofpAgA4M5DWAOa
2Ih0izNBfQOZKGwDf125lACd1EXw75jARPTRYGwUGHcS92JhFIGcovdXnH4ryIXr
pYFTI4QC+OlFQg7s+x0cANI4tfqJWOk+3WN5aQJbI0l6auIHmQDa+bsaIyNrMJc6
nRq+h/pxvWwgOqc/6AbAQKP8J/mqvY5WRhsIMxUXGL/oTyvtT9UrWNXCfVIb9ISY
Rz/VvHCa10SzV6Cj9gYORs9dXQ215YAGVgauIqE64m4TUfMbyC6oHVtkCT+48/yN
kNflpnjCsBh3/gD6Zkvqcril1ITj5s52WwoPmExKI0MigqtTiDgYHn4taJhnG3yd
+EJ5yPWDic+Ql0BqxaTdYmGCQ3WO4uqjJBCpj+WE7ZEp9MFB3/Er90Vf4TA+Jmg/
3XFWBf73GDvDEdhveV/hB5CUDKdM7mzmIVF3iibOQZK1Pfbh4CXnfapDKA/3Tikc
YYcKaJOEs8TGbJCp2OWAdCwNgdrbTDuWni+G+IBhDNDzHKBHHsB4MsjYHS2Q1WPg
nnGETIrvzT+GTNyDo0PiQ3Mlp9KXUJP8nJZ42p0KTztK88NPKqI6lT/AsuBcVCIY
FPfjkJKg4lqpgvnfsZoXcl/2bbCAsT30rIMJwDVujWMtpL22cFCe6hvbhLGin6Q5
pvj2fX8SFo4OeGuir1u9P8luM1+r7RwrqXti+NkjBqHQ1N9LHv66qydjAtw7Gmw8
ZK4F2qOiq6XPSWPMBivNSg91kuBnYE1vILYesmiNAfpqnIVTU8Ue2YNtnyyAmW2K
MWGIgyofCA4sthnJsGvdEQ+d/IuBroMtp2BOs7dqO7F+U1J6l1DRAh3sTio+YYCc
XkrwcP8/MWheT/qtieU+Oj0Zpgt7A9TFBqmb+30D00aASIP4n6J4+kgNH4a6Tvvu
M8G/d3CqXLIr1D5oyOAVFjnkg967FZbVzWmH3PaVYMmlvV8iW7W5nO06Uy+D7i2i
yBdTrX0qtGBCQrQGspAuvCemrVvFS16CJLeyKp0QeG100gIl8VaHLEJu2wrsr7Gn
OBzE9lfvvX5ChUf5YU0QECaGWCfX0kPTEcZshijdjf7z/d2cnnU8eUzXk91FtwrI
Sf6VOMFtdd6ev5gEWGgq+6S2WdWtGLRTK6lQx2idvHHmjpyRQuAVuR1NXqJDK+Jc
9EW7wAgxLyZVvytcQOyN/D/Lwvng5+KXOy2pXtt+Xna7XHKHuYQvof9ecB8M2YRA
+brgXPYKiwAkwbKjWqyAT0e1XFBt77VSL1kWBVHCkMw47s3InyBYRMnjQIeGg+dg
7BzrB9pfeVS0mQcBkGwYbOYKVNsc2Hc2FanjV1ivWDG8KQ/BCuoHytGJkgl91QC8
XjpqkdjC+V7B7Q6TEhQlXj06C2Vp1OT9ETvPvyD2kng7N0oAh7vXHsSUfg5SgsMt
0Ws+GtSiGElCDu6DU/cbk7+38ymuvqX+vcMDIRZlJWP67QDEVMhfxummKC2q0u8s
UvM12WzNvw1TJq7eytHqiuRLKjvxLxlAD1y4HzQX4tWO2MmyjlK3MCbL6+33ardm
7kiFIGRsaelJ/dvxNLkVj6QVBoZ4xrB/XNISUO8bMgQ83RJeyMGPgJXZ0sR+UFz8
xDtRLS7STJyUq5YQb2Jqamm9C11+8B6o6dqkVc81uSTZEagiYLkZWLf962UqHuNg
BU9mpb3DgEDBJn1d0qROBtV34uT3cOfmNA1FJsGmbVZYkPstdfrYIQk9gD1Ulpub
kLgamsak/ilM3FnI5NAsaCc6u4Q6qzkqQGnofetV2tKD4BpsjD3ZBOe1v6uNtQHu
W1qweLHcOoFo82vHI/I+39zCgsI61nAIc/MLh/kMx52ziXSAHVLSfdoGnFYz/A8V
2iycIWiICstGhELnirXa3b6p7DshSaTNlnhq+7M++FgdOEgZLDW2iRzBIh6/JWRk
VIfKB4mk6Xcfl5kwjyYt3UyJgzavcf2Fu/BVc3wCfZjSYAw7Tdf9RlQgeJLF094y
UZZsb01wy2bU4t0U13y/M5iEyIjXAnoifYtr9Sxpn/yBOEl/YfJ3+bSwOLfAu4UZ
QnmgC8aMY0dscpUPiW9JGODNZqxxUrpLmHYxhihI9TZT+kjv4T/9dGCefwPhIC+q
5N6gXLb4OayB9F/RpOoKlPRVfhGvuatPT6AUgg/+yJLKyQ0k913rF8cd9KYEo/rQ
tIafyONV1nRhRW81eWw81JBhEzvb15QfpsIg+5qOtcn+L6e0+7s2Xrg68dZHgmB+
xODmZghsRiaYwkJ08xqFfFhTCA/aALVp9jveQMRGBxyVcKfca84q3gHDU7qIV/uO
AIsTpOP+3t+wOTkeonL6UVFJicYPmmgLzNV+vNTVgdJvTiBrfIUj5BMRXpy3wMre
1WEsQf0YiJcMR0/E9JyaT/lj+zOerpcf+padeINxn1G87//sLmhKXbK2f3PFe3HU
wl1+2zaodluT1m/KmnMza3XF+VHgYBqiTtztesN9C0SpCV2okEQ1ubxbs/1Rm8rV
O+z/C1Gdz18zquXuXoAch2eeE7IqPy4KP/NguxLTqYlJ3XKGJ5leUw8wHqEXFSn5
HTA+yIxbmFjDn1y3WXzxX3FTxTbA32jhzm9aQlKw7irvxRv0kTGTGxFEUOIqZK5M
BVrTUTn7aCrcIaL1Yqsa61GkJN+v7FIUC+AS6JpWRwjJG2fpeGTyw+PmQ6OAblYr
VMA+uF02JQpSDHioQXzYlq8rAenizmfaPy5MBbxzceTUtCnFYyiZV3jGI41MSP9g
/kC4V4dddJBkuRjWamNmviHKzTHKWkS94d+KMZuXGRphJZ08QxaieiFY/1sLk8pn
7ASV6jPP209MRKvzF8qU80l3cu2aLPXQp7d/GFHITndCxnQwWEpIawJTRDKnCnCZ
JEFQxf1BrE4PBCMOW9yqIS8N+IYwIZWSPnb/xBVO0CDsC8igf19kAjZQYsNENI+l
ugcSCHhFVqpbX5QA9QYoqmx0DmCyqfnQX6m+01iDwVD1fK7Ld2/tGVASvGrtDFMR
8Ds1pfk2Uw2kf/G2D9Uj/J3Ey9wwNlQQLkyLh/W8S5lD2ghdDM4UPlZfh7n1kzZa
FpLXKnuiXF0jPvnm0iWedQ8EnxP6Imzz0f8KnskgzLTjL6SAYOnCER/va7JassuJ
d+C21HS1/jiU1A8jEsAJK2f4l2yt7uJBkkB3+bkBWIiWNEKY85QIjsHZn17lJEl3
1Kt3aSPs8g+UjOwyQcuqp9doRlv7ZQr0SVyJzYnM1wVwThQ/4nXI9TK7JkuEGy9t
ABQuEYE3S0Xr59sGJNWzZWtWN5+JmPsH3y1mHkPRC1+Y08L/fqyHxwJsnlvKlHzQ
FXC9CX9WRj6NKE3L3L9IfFaJMR/1H4GaqzUjlo2QqFD9q3WzI789splhe3YjBbDa
x/nepadaZ+76nY6XsDeiRYrBxaiYLLJrD/OlIK+Db97U832kqEveBjDfFBstem2b
hGtq1tOPKvIZeZ+gEsOtBO1U4iiP5Si4TE5KMVnBW88bIacrOVZnRTeD6sru/Kuz
79lVzylazQ7VDo4IRXelV9r4LhljCUNw2hdAp8FER0NysZfAdRsr8rXv+3LwTyBA
0vSYdsTvB1ilV+5W3EdT2717ygX7T+DFNz3w7c1p3IT6ChHBIWFN24fVRCzeF4mW
5h3b7p0ApHNWNnj+8ntTKxTKzvSf1tZ7XeoJs//dpqHTwVLKyJNyY0fjisy+7hpW
Zc/wEsgnx7aNWhYZmAVP67NSe7qfrw4bPSmuZy+oNqi+yhD4N4NkPDWIUXSwB6Xm
2fcCuj56itJTDGe2VBlVB8bzUU9tVASE0v0q1I/1urvx+IgAOWm0vL+HlPDTCDuO
dTd6wAqvqQkOemlvbmbkLi3Wji4pcpBtWaHdvmmcr2971DR5OQAvxHhljzCKV15e
LKm5juvFSLxJBKl1SErnaz6f6Zb5kYhVScD8uJjg8aD7+puYG0kmUiAWEMYLyVVu
4ZtlNnxwnHFb9s1db3Evy5wCcDH7kpvtbzEhFzdd8AniKJcOIsy2F/24QV5Wpaaa
Zt1j9un9fWxg770sPQEifil91+ChghzkSYnW+Yco7dVvq+LatrR9ZTAvnaE2tI75
24Bp31xSbS4WA3tiPUbZ67sAclx6qOkD/m4CAUwp7xI7Xha7xvUrOg/AKdCJ4FVD
WJGY8vMIdD1ZovzR4ObOyG1tGbiuxi2Im010HWvkHlDPkQwRn0EiEWAFXTOSKkQ7
KdzSsYugFcK71UJV6vaXu6OUHPsegcf02fgCkckowGuluQeukS/z80pvfFhI1I7S
KPh4XsL1mwS4uafaCyzMhQvt5pcZGCMvyvsSi45vMCyli2/RYzMi8SeFkPSITedZ
oBRIlJZkDp/XB5boplquDr8nemFEZuOJARB0h1MAJTUi9W1YRWwG0dLp6xXCPmdq
9aeM77XHxEf+6+934Ay/YyKRnePOrwsVW8Z68O/8sKhKx9qjRflANn3CAS/szu/1
BX3ZLTnPZ2s5ohahFnlaIzIMia92mdBSbYBQlGcTbbyFaML/C9UVEpvxK2TLbtgU
gNcK00zylOK5hVyXPPi2dKdOb6RVrI+sfj5wq+e3pDuvozddEuPfEoHyRs1kwww/
5ewKFyaLtDZByvxtc0xM+W5/RCS6clwTKL1sbXfdmX0TLqazO7/DrYIupITiKwF8
ySsI2DqrlAZWbtBfiO7IjvrfO96AEN119h3LHl1gNOFhw0fY3fuiOCa98CGLuUDI
jsPVlOPcJ75hgrrjxCIWspd90HJpZ/ihKXVmyYnUYpw3aq+7wOeYO7aWdSNh+wZc
PGTq6Aw3WM7YiYEmVb5E5FrW7mqCrWCU0TQms8JZVkZuZALmaQ7qiXNh86GgWybr
0HBeBISqt3w9YKqqHQdK24Oifj10n60voqeE6sarVTSwKrKPnCiyeDJ/6MQYZg52
Bw8StE/EzlDo545sjjDknzoHLOhA6S5mn8ZxhGC/f9M0SV5g5UIFno1W28fdZkSc
k4x0GIw7IUuzcUWMcxNz47b0f5p9ldqbqFhEvqwoXG73VOD63E/OPkMnzIBpft/G
J4OgIAU7IiVmCX5zBAoiXf9RKIDLI8lTFiMb71edYLNmluDzI9D2s3apiGXJnmAi
T/DjqczvaGLjgzbQjly/hlDo0zSS3kKoqYwx6/uFwuRCOTIasKRxjMdFjofgMFBZ
E2rE8d/FIMXX4ZrVgGmwMREEztRIICX7LDRgajYXxx0YwXnk71ptwKFXzvPLAZ74
cQVFODe0NANnkvDHl3FAnp5ZseM2RAOPyrWbKfgxraJJH1dl4EhggOEJdo5zpZdN
wZRIVRyij9SlUSgrrFnz8Bee81irtoLlfaF8kqBDHG2YC6P1JGRTWOZ2u11Ez3Cn
fU68o0+le3hq7HOi/abtrNWt4CcTDI2NSH7Dfwy4rVWeFG5Zhv0FwzdcRe0G+pha
63Z9hjfDy8WWjDlyehtaKBg1q93ZNwi9WBos4TKGZtLpczhvOPWFo+FuGYoQJC5j
W5UNQUoz/gG2Mlwlm0Or/p5HUsiMnx8BEvjhPnBwNChnt8XluyAaDXhqNYEJIRD0
uGhijNu4EWj7yTM63MJK2+X1pyforbDfMoWQWm6duRsrO3t3USjK4Kb1r5jIIcbf
PFsOUc/ViU8TVWJR+gfSkc+JBvUDoFEz8u6mPwSBHHJzXQGoT2oEJn8JJfGbfr8o
O8WXS5i2JXvv3/Ii+ENLTD2YPKGzbYB3PzCBZwgQwplVGPHsJmdi/b5nRK2eSSMP
1aF9ANVlBAy2QNdSwe7GTrHnpZxtQUp7XC/nfBxHi1Mkcjh05fJdk7uvibm1u4et
7ZfVTqfesazePixgIZCef3d9YQp+aKySbRreKuCqKY0QTYDd09Fk4k7ZYrlaP6qb
r7VtEd9lwUZxbml9RiIOy2rGl7GfjB//wZDZ/1q/aTsuL7LNh+56MB0VH7qMqzI6
FZ/QTf6MvfW6hSb8H89tjSxXd2SS3fwJvTK5HQKvYr5f2a6s6WpwB/zV/o0ua4+P
NO/xp6OeI+tapnSzL8gQXEUcitMYDAk6jcoSVqYT/QIto96z78NF89anRtyjgm74
FUZJDWVVrPIzOaFOzYcm9wse35pJhkMEH7jN9X48aICt7DHW5Jh9RDpWI0kMInBn
EUDfp7ysm3IHSKWwq6+5AhNuRFIOgcG90ny8sp0HRf2QDR6BT73vxkgQSr2IDbe1
ed39RBj9AveRSfPvIW4Y3KVGIgpzOnZTQ+VNFE0zKlUglcadc1EEQuj6mKLAMNF/
8hSIkAq1LMAl1tCUhUSpdgWK1x6RJ3RIjyNxjdoiJn8muefDc6u1GhddD4jIC31J
2d/8MXfBu0m7FjR9NxtRSVRHDepkCEfgCdpj8yLlRT/tldyXrszKuCEy/+TGbfBg
ov5J8Sd8mvplQoVX8180E3ABIJeOhdj32Bm25ejZbXi29/UGa0DdyD2gnZkoFsNy
oJUfchKNtmxVn3TGHg1YSlCPH7G2+jIz0CTQwKfIWH0GvTgkabKMpsuX5vcgQnER
DbQHk4J3S6mNi22QW+WIkcP0EWSOZYxqCS4fWQKE1yOx17ymY+AOxSOQBX/aUT1f
GGh8dos9wIlaEtMrZ68LvW8r6nRAfzhj//jy0GhYYTCjAgL6ZqcpvTC3GO9aDZSY
H7+nWVzyBcWd78qh7PFXPYFtKpjMGS+VwscrzWwmkPzlAa9D/KKcOyx3cJnqAIDy
cweT3Ul2ayJ5fMHnnJLZCfGIbT1fOaIwqTqCiu7njq0G2JjIYTZQdyJu9lAaqS77
hM3bqj+uUdYqu1Lq3keknUqp6lePxVR6NGdHU6jmSzz5XX8wrfwrhLjaNUmeCAJ7
t6z105vT5p2o3rmAp2FJperRW/qBlMUgp905gJGdToaioVD8P8glej7lSolpstH2
E/1UHAJLbrroeJyofbZiEN0y1MBMODrar+9Ihc8ypUcoHjRjswcpXtYdFqjYenMm
5hEUw1BIAX0EwVMSsfm6Ng4Avqnhq2qD0CyQEDIK3p9RoeHIQveRPmgAm/6lcNBZ
61w79S87T7WenmF+TFN69+zkIHtyXY960OCu8jQ6pAR4pF/iKlSd4cFsALy+0xPF
ipSZUVFA95SmM6uYQtqLsHECIQHSc95cJRFjr8KI0DlkFXjFNMNbHZg/xmBXHSrP
YrCWzVxMVndQLWvSRLGlXfs//KkcmgkPdNbwkmgSyWGzrFgKHzl8C6fEnpms/3+E
QTP90t8bEjeg7zF73c3OhRPK1TrvbHgmCFe17/bylprIRBWUKgJMzGc/dESCxceR
bJKWD4WAkE3rE8q1qkTJIrGc1uvvURXHxV9Eqa6/kdJQZUnvWr68b7buyWm32SP5
nuvhf+tS67pVDClS4XD0T2DStFSadHLsG8z0QF/TT1ZHry8DQG1KcN51l3ERkTn3
4OBDPqd09ZJyiJvjXBFC/lkcgGWsP9y+HP3KtQaEfbUO2AgOKdV1IhLEvpnNm6+o
Xk4MKqFsw/+JaSBePWLsPo845ILqC9uC4XWlK+FagsKBuTK9OjZd9/Olgl3V4Ur6
wuVIUAyFu4eHmihhTNAiaSvmPh4quwrEw+K6FnAgV+HFIuP4LLClLLytavLH6P19
1rv0hUtR3iAHz9q9GdA512kjsxVt3l572BNWsjIM3wT7acvKGcmO26FOn3lw/pd6
gmwamIQtwZtVlhuYp3FvgW/pmYSXoUeEmLZRWtqv65foNhsUnYGbftcGCFGEo3Ah
CGTR9yVi1aqXBm5NygmxGuABJJIcUF17KvZMCrg77cdNGYNl3dRTMVnqz7k/3sic
NkhIVYEe+mzUdx9W6F4JfHoB251PD7/J3yYU4RQs4d/qnki1l4Nw1/QgDe+AKJDu
4T5htl0Vp1YvZEQkSRl/M/RYIkXT8h5mrY2N6fJoX8SWkFGL5PDCrEP28frIM6ez
C41H4c3QQ/MZ540IsCX//bDgAM8P/q+eUWle5kw0YgLEmLjKmKlEROEFLD/goGjC
Vekw+hs5FY9R2VMlvXwPR0Rkul8BgJuV2DixkONrsa2ZUn02BxETEyh4ySt9VYY9
FMQj0inxIhUNXdlSbh6LVys9uVzirXVJVcQmjv4OrBrEjAjweDb1ot24rxq4Mh+J
AAeg19ZNNeO3DLfIdGsI0l3GitivJOyRyjNs8K8Nh7oXdT6x2RyXOFBa7qStjs4+
6nBaucMDSoXDm0RH/rqS1HiP+jXnte41MXEzNEf5GD1fjQ2P9XJ0qbuxoHBzuXiS
idTMP5uKFAeOilzBMC0JJnAFQVJQjIInO+/IwsnrVEFIjxA2jePgA5pFpkncIGtu
3VdOMQKixEEfkaPtt2g2AdAoQNFz+CT1+l51JUJ2Vj0+BHwhvayyUZdO4p6l+O0S
HEnvfQdwx0kENeq8+bL/Kw5rnwVufH/PCGWVjUwzDGXPqjzXWBH5kAcFqYHS6NIu
ag+ErxNLJm3us7oE3wBZmLxRc/jmsCRJiBteuHbmfZbYvT3CPnxNfjvidrUueWir
dZJ0TAQmak2rsYvEY0wlTSdnW/Tm2ZLjYj90aa4DFyUUeFFYnOG+uuHHM8L+Nuxj
0yotko/dyErZHeoj6siQyyCOQvsrmA/kbS99GH309FMF5bfWOxOeppwJ8CyBvTGE
yL07m1YyUATNhDOUB6A2B0aWQNkYssX0p4wzXwumV5XvhSOy6FNflKbmOykzm7SC
JhR+W4fYRS9nE6eXYuHc9p3to+uUPnSP/9xv++f5H3nnkL3M27/YFe2nJ34ss++b
c2VtZTdqz3HEmjcgu+nQMvh1iffcHRmFqDamUJaPNvlOMcZBOXBgPw02jjyYyaIG
y4pzVFQ54EPe3obtOKIeSC+Wy/L9m+0xpnto7IMkma0kk5r6LwZzNdibx+M213qh
4WwkvpyJlL5eQUvlybKYXLqkz2kbOSLq0dpJDE5qblSpK2tadG8iKy6cUJckTsrV
DwPZSnaV6zDifb7lU3nKzh6pz6lF+Y/FW/bfawvUnyqVD3PhCL5P4pF4NrMcPIre
MuDIvXpKbeXg6jr7S797wHdiNun3PBfQYMqKGX9ifiiP5uNaC6qt8gjTarsNHpPy
uMZct2bV58myyT4RBfd5Ak7NGgY8Jhj4j4yZLA5C6Tmbbb8PUmcr22EqVtgxSiVM
iRB62QxLlURW1FubP0eYvb+vJJ2lVp/V5QbhgQPJBm85TpROLDb6V5ZqF+mlIpF0
k5JpQw1E0lHy/Zhtbh4DfjqwXDNh9J8IS3X24Aipn5Nph8O6cTpEeRLCaI9CBti8
ACQ7UBP+jF5gEUsikQnIJo+PTikurw8W+j5U0jYHPaDhqrJNVf9o6bVEyheI8XSm
YcNNBPs8LAExiCBmiSzPDEwD9J+EPgV72w7VZR0W9AcYyjnNufj8elEprx5fWnYY
PBldwSzVGWxZUBVOMSHTU86DdzCCpxqoCT/b2tJESa6QrOzkfnUDQTDsWXqvt7Ss
87fmLYA4IBbpbyFKZ417anOZKlP48ZX/BwVZ9CSPYksEONNtqcUwa8VKSFOCQMJy
DuzAuRTKo6rxzLO5EoMSiYA/m2G/63ogWgfvfS7nzhruL33k0fR+DhYZkXpineK6
l47zmQNTgiQlX4hFECpzCsVJMDXfDZcN38kf1OuACQgITGe+6Da/XGn+Tn2/YInn
FukpTd0W/h8pWrxBf996Ou+4K53jg9SZYTCKrGvlq+zHUna9DHl5KPJi4sv5UgKk
I8vlDm11y1MkCZRYK6uuQJZfdVs4Cbsl/VHM8d2rzbVEiVUIpJx1Xt/8dMi4mFa0
ILhcGo0mGH7t+cyR+s27PtSmrjeVRJycEWXHJdReD6yB2ZSHxp22861DVKg971vj
ddCYJoqiEgpnuYEEl/XJBdzmMfRLeDf4uTNsXVgynrkzGmaQW2Ik75GREJcoth+0
o+ydo53EWgx14+jJ9LDahSBcS01IWD7HAqetXOxWXSmur39YVgZAARK5yj6XVApU
yK9RTQcXOwVUMBCJ1/v3T+Y08lqQwQDFrMi1J/LfkrwarBuJoTcRjL2JaoxiEkjG
SRYnGH8y0ctgUClxIT7n8kreofmdFjTiJPl0bLdrWSep4b2qbSi2Wx7VxgZvNpFo
wK2J220GQU1L5STEUu0DkZXlKxqncXJ0+exkJRs+NXOkS56UfYm/fh7IWF9SssNm
kkAKzkQiR5USPkE9aagp/Q8J8726g0IL3Wn38yeoAXKN0t6eR1J/LNwgDH9KyN92
gOBcSNGvE/7928w2Jgw9bAYXAZTvxD3ua+5PcR8z/bQiJUAjWbmvSq8D7NtGXkGu
899C0V0+hbTAgQ/4ujXo4cC1dCHp3tvsBNyPzhODy8Xvg9UpyPenNhKPujeywuh9
7+WM9sZwATTv5t77Svdc8B/C7F6MneSd4lFbUH3XtDAkCGMla/lI8iSnhUZlFO/6
qtRUfHXh+aoI59p2Z6b/SjYvqb7L2ki1b/8uol0odmhdeYwyRLsMAmJMVaK9/a05
oKrwQN+feHdPJgFn5t8PyIg4WJu2c6I/LekPRSQYSe25DGfJWuuOXcf6Q4z61jXB
SaNRDJy9An+f/hjZ+SXnL93KnM8YR1KAsPVkLN7DQGkJ4ytsy1Ke4+WdHselvpOO
JwiOz7SdqZIKt8WCC/SUf0+M+AluU9COiv4zpPJCGuAa4IY31+/YKe12kV0EmCYC
7zOUla/1UmzQjRKlXC++q03hdNZp/gk+8KmO1GJ5rbJMsAVMr1l0zLUNGpHqzYmo
y1NWv90fsEv3VHwMJORJW6sR5/ZZlz5r6x7HCCY6yeXnHnexcQ4PNRIgyMtvJh+A
R9k978JCZryD+gDcCfKX7ad1EVHLHuQwUDk3e3JzE2J519g96SkWzows+dCCANrp
uDBjiO3yN8KygHKvL5EAqUmvb7w7p0fANxwGa5l1SDKrCEbiSD0ZBVs8f846av6c
nBOitD9yb/kJgPv2UAHwGm3BDV0hH+KRS4rIa0XKpKMWurXQi9oHviiaaIPb8laS
VZmztWI0UcgooOAn8jXLmY2pGGW3bzcmcHymUgN9JmYaCpXhpaHUhLUctqPXATnQ
7MfcPRqTNWxxy653AFCAhBRY9Ezv7qJkGvOife9sQ1xrHEvoso7QUSHUCWX4bgIU
ek525oKMhGYQdTF9GfaFlR81Olefnlv+EpLL6yQ9WH7UdHhwFQCPv+EPxr3AFfdc
6C/BXVbOiI12cy8uSjkl5Z4jbnBk0Mw05xAE/Q1WP4AOp2TJ4sACTOkRhFV26pBU
y1rGlAqrQgkYy1FhuJu6vzh5cdT1pHFBTRKjX+fVtg5C3nrb3xeUbd8fXap0LA8e
CV0DKUN7f9KSQ4nbjNMYM/JJv+/tQWksvW/PjWIaye3D9Dve3f6lLOJXWYX3pl+t
+QCE03T5ruuRX6hhREmeISk9gJiXf3F0n2KfgXq/tEUYafaIU9fny3MYAh9rSLP7
wdw2pYqeZxVB7rlkCD9f+vhz7cfdJyGKjfFzcfw93CMe/TfvcpIZGnQRe6hpL6Uz
SaS2BJE7a0yLXZ6E6EmmI3lMlQVpjxMp71zWNEjbRG6hhs1VrgjpgXD7Py9r2FiT
vb67Gtyg6xRHLdut/4UTqNztXnnjR3/TbgxBMPO3TkwXxyEoCYPsrhiprxnseaDi
/7DLTaxXoxyn3Zonww6j5iX1MDivKPE6+NMWsDKbMKE6SKhuWTyMXYfjrcEM8CWC
oCjs3plP6uJQU4PbXx98HdnHdiPqiuNikJ9rQLYU2LzU7AZXWncc6j/ZSxq15OLm
rX68q5VyQ71J9X5BMpGdyJNurGThG2N3LJS+wzVyWgixao/iI0XjxP4hU0wtSgZt
A8FBrRDjuAWrWMl2K8ysE6WiyghqS7vp5mHk2E4P7za1nVWqc+X1C60eKuc7X+6f
8kteibTW8bUNwJO9voQERYqytlN4VTCIzwmiNC+vQJFBn+2rHm6/YbymTGVKPEXW
CmT/yogdWor1i0UwyQfZvFWyegSL+FJHqM9X0Bw1tdos2YqXVsPmSCtNGkGpCoOy
915bSZmmO8sL4VZiuOoMMoOKZdHoMZkq8IFBANiwQ+BY8EOA2WfC6bidTnmqpbt7
aqczwIQVgB+Q0h8ht0398bKnae/dQo3rH5ZUtATCI+QXs3h+XzB63954Xffh4AvP
1qurV9sGkpNLRxuKAckNO2oucx2tZ1z+U/fVciOqnxQHJU7av+XNwmk2HPs6maN1
7+TeYKByfMa0+JCCVuocJqS/EjkGKFvUwu4+65L2oHjFDlqn9qsiMTx22WLMiqG0
Pd18Wq+8LXJNIjV3E4wDPYU1T6iLskMUlg3F/HTgVdCGq8RyFpo2x0SpwM4hXbMI
I4vJvpHk7FzXwz/I1FqAonEzFMMexCUuzYEDolEVguTX3xIJCSSx4Eeu7m2WPc86
WPy/EO29honwq6F6VSDR+bqFbsysUyqHbCsqyhswz3daBQz1OkOAfxgaVImKQJ7W
etQc8ijN+UfZDoFj1bmoYZk33vMj2gOOTQEGWClgRu3nozIhuvt/UYCursVkIqNC
bvXf6twa5FXoM2i5/rWCSgfwcC5Y/QeeHcAIw/iBkxuRKLQEiYFbrLNRpEwgyws+
/6Z2JCn4UmXcgiOR22xFhoIQz5g1A13g7eZsBfnBQhQEvt9cgMQc9cqju6AWFzjE
1+3tkvoSqfgOvOvpNmoHwV2fGQWDq7htINXeC3DBXaTdchaXRaLMJ09X4CLnS3+d
bUn6mgToXVfcANvvm4zyu9KI5uUduwrChDYO5ARLUrplOrLNL+kbCgAI1rVUgrIy
7TnyFrQxkOwV/xOxNZt0WEwrdbNnyQTBX9Kqh93SbcXQJktKQLkSCuWlXvYzWkAi
o0JieFy2T6vGZaw5qNkSxJ0jz/+Tp7sMlTrKECBkPzZARCRTPNqfn0yd8BGnwchc
4WMhP3B9/Kh9nZP0ngM5acLUNWZTnDX0T1BViclpnyLfCHKHpZ1TAxFmFXLDTgdJ
RCcYiBrCh1sS6sXqMuLmF1BYijMh4TRP3JfBDJGMqZlIEMt+IVcsmuUuKusLdLK4
8xrDi3f+/DqBfIoLROm8pMaHz2jgRddVPMwL/uInLhODqcExsJjHVynbbhI1ykuE
ln11psuQIGdv9Cs1C+27bwH5+2EJ/xgEbVuGXtHO+tVwk0udiFIML0w3XMmWSsJD
DTY5KbRCBhhBBJkqtetJ4dO281Fp3KjNrbbjhseXQ4HgAESeK71ldog9bEYCZReN
qQcPLVo2zf9/ljfgLMFZYaaZmW3c49CUSCVKEMrsgnvJosra82du+mv4zceJQPIF
/hjt8EVcoRUVhbnvi5uMlzJseBkbP2AiULV8N3C9UZV6HDUZ+4HhNEIgBGfJakOv
jy7JybbsXoimkB9O36b6T03vcbJzrH2i4Nx5Vv0LGlL6FA0h1/GgJkGdLLeZx4RA
WSyKqxCaJwRdGrDAADrV1uXCyf5RJ7233kAc/aWmtKWG295Jl0jEVQdGbjAxKhKA
x+H3mU9bHZG7vEKZh9l81jwhmMr0gpLeoWhk5jaQevlbPqFXwGm1mBfo7XoPqi7f
wB9kK4nTpvVUsV0C9D8DIpOMZMMLof3HxgK6jLt24KEGz+G0m+DVNKaEzyo8KKox
RiLiu83Fscs3Ck/tvbh62EzEF0DD6Sj2hudmthafa7YYxakmgony70XxhhBg1Mx5
WtVvqfDBTzFQOZ0O0PFQyRRmS4kULlKJE+mq3/Jaa7ydgt1K1QfjFVAf1/nWR8SV
XbmABPjuIkNkzvicQXsyjPm4f/tXjfTWWh4SF8QNBfkEC0U7ZETszhodgp3rhRRD
atOnmF9RFBTZRHn/qOA1Usd0TJ2hHD2l1AEssZSKAQZRpUKY/Rzo/0UyibyjHPj/
QY+6yXGIE7qAy7/ABoFDzNJYXB6rLNrU2VprPkjYXP7rUSJfuEpTqSCEcZ3BrMu9
kdYXgaWw3rHJNTXVNvYYuK6ibu3ORtQ1j/Mp+ZcF40+7ktB64XkAqKn4THQzo08T
y8FoDF9Hu050lzbGDbnPB7bhmTPaZPIbtYOB6OF2NatbzJp/pQnmlImFYs6+tY9N
65tyEqMdf4gsRNlj0OUL8SYj545+Zw870dznFa3a35+CnShb8S8Exfp2tk93hyig
65EjU13u8tTLUaiXomy3NZD4X+M59aR0NEplojFW7DFz4mm/Xen9Fraey2qAURbN
YQpYbwOrcMX74pBlzkn0SUZ8ceVeCakgB+W7XOFgM9zW4AYsXWJCBTKJ6eSgoDot
sQIjU6iepo+QnrtGRKxww3JC/llcBo7tPrOiBXHBBLH9QsFM5T6ap+3j1BS3Vmyk
VtKPxYKphy8XoEUnAb3RZAJ6DpPsh6tuzY+9PL6OHb/gr7kqKX6Fw9stfI3jDv4x
Ljg9cjPqR/yi2zoWOd1ang7KZrN5wgA7RpT7eQnq09tE3/hbfyz568YHttloabu6
zTkGZif10bFGoJhkpZTHvWeZnBXf/c7gsCdILF2slWwhYa1LlQjs8mzROAcIivAe
rh468QKWt+50x193DZjAISoTKFz+qyTyTeL0RClaRVRV+TCqUK8IYm3zEAQJIcsv
46kaTrAkyyftv04zvkXlcFmEbf83RyOGmTWjKvltxEop5x1yxcCy++eIa4hkxX6c
flnNBoOX0FmIHIVSPW26eKYMk2A8Hid7kIvg2AIARm75OBh0JeiY3XgLUFwZpMs4
+yZ9bTTwVujZu8E1R3AZR1QQejv5O3Yf1Bv8q33uzz/ighLtEbyb4Gh/6CBEAerN
9a1bixdvVvkUdiYn/h551pVhmf9OrwyTssk3gdXWVU6WiksFAw6w0zjRJ8m3Nnfa
VmJObYYqNrC+KqCnUc6+qEhQOvo1LihiZPmXH9a/ukrfUP+gY42RS/teWQyCxOHY
vD99SjfO6zr2NwqcWo6ZVyGZoTd+DPlX/XUpK0WeKQlfNUEhh2syqYCHiA/4aan3
6T2FgAP9OpyDuoHs/2R5Fq/dik6lDTAAruMlptK2oACwEp0BDkaouBePsGNnUnod
tVsveYwjVwtxdhjBU/puwCOfHV7RmqcFGiJw0adWPisVQ2Bh0mrON0njhWq+7gdo
g3Ib8b3JagemD9VxUqbJAf2tFyzDGTelTk2fva6t1egkDQ13ZuBfBWlE5DO1+zcr
qB0yPl9a8oW2rDdtwtPgHiCA2bWG81AzF7Xu5khYUuruRIDnTOp+7DVjSz5B6OIR
c9L8pizhiGEpZ3AzAq4+wDvLgGXSuzGrmu3tp1T3zIApwBX/lT3gD9BqaRSF+ObQ
NqmGNy+CoPtQngfPAeJTN2yZjPWzxHuT7LH0BycAGNPfohrzUEXmv+QJWw4Uga49
SAdlSFT7t9TYr/pCYFK6mJF1jRI4hgaoYWOkaVgsJl0aEltHpO+Fxy8Lndv0hGrZ
BSnv+MkFRQw8kTvo6uDXWZ1M+I5WiNR+kzH0SJhG4/7nVfYPsQen7cQBTpApN+M/
04FG8WQ+Gb3m6ggmhjafmtyCJQcbUiLWrjR+XKoWBmleA3UaqPa9UCQafV5srBkA
1dTRhljsmmFEicIZEurze9Dw0/x8FrXjPOExlNO5sLgfGXWSwX4Wk/OuQsF+FBMt
/SFApkn/Fg/6ERk3RT4jsdTaVwcPbQ9hFtNBJdn5QhoK5F4+3cVql8au2+Y1ZdDY
WrllQ2k0XwrT6oVurddRRrsQu87/fyhVL9qKyM6/wWnwXmJMdJ+XRRVDlDaB+whp
xRZyA8zIt2ako8OnTqERA6Hruawe/SWSAavrhfQdjpKUWkbW32eIVnJ5dhadvBgF
+Bd4/F0PTzn1lymIN4MLe6PY/uX4HMYEbFB9Q/QF0oq4FaKX7Ax+BWBdBNCGnDWS
ZPIoMjLaeG38Z3uNIB0aKNU1ONd5Wsl1KeNN4wfaBi7Urf2czR5xLKZeZu6uAE4v
gtkIt0Wuagd7I2X76183h/nTeqW5pJqXRFOKe55CixgOKDpexxWH1JWhFKBJhfmJ
s93plmBevgBRJOoP90fIDfd3q/aJCAKCE0etRGKvb1odQCHwMQk3I3bju2SIxK+a
i541SWOdyleZ7X9NIpIKCgSGwumJEuI+1+jbc2aTCKFvdoAL2pPC28IvWqNJm5Bg
cBIG6NTwGgz1gd9CwvGvQzdgJMDl9KXlXz0CnVb08knsmVTg9PAt1ZEXLKFXmbqX
+cDfyxsjlqugYY2ZofVuQgQaxZBykwyjaAbDtmqv1tbtIHijThjjrUrv795i4DE1
n1vAZ0xqKYlkz4OYjgLMruyG/HnNa/V/OpiEtRct/AVLpJpgt0nuuxQZByM686xs
DCRFqA54AY/VJEHj1Tf8TXpQJt3wU8U0cG+5X2isolvHk9ruSqPMdZh6mL7UWDKI
47oBs29bApKvHhYsppgvP9oWvkOX9SffeL9o1DAlRm2wMoYtQQyEGT3rB1wOuUnq
Hl3PpSsdqis3hcYZrYoXG/JpKzAmPuseBEk7WhOzkVeD1+hgghVvjCcvkfKDUqAr
opslX32QaRF2d+/V9uxt3ID0pTV8GvMMgwR0lFU1OQsGjxj6TgSYazthCWNOrQ1n
LhsHAFYgMDmPuIUbXFz1ZCnTgFrdMHKYiBCpVTm83f3gPvWK6uPuC2+6peE4pEY+
nKRylEB3zxHxXicPBcsKM/TUAASvRnlAR23E8RfUS/tROnxQIKcA4vadvIEmcXYd
ESDeeVOeBTQht82Ow1qLDRw6xG2syJGM8Om5IRUUztm8EVcaAL5RoXsHOTA83uuO
krR1dVSCDMzi7hSR820iJXmqIs8T7Fl8YkVAKv8Ka8NRKBt9YaaZF0WJinyFqBGn
0jkVpiQbUddwd45aXrgx986H46HtaIQX8ddbvmcs9oEixh3Nzd41stS2r6Idhl3s
NfwU5Q5NK5dArlBvYt0C/URBeqBkTmdnetiEjxCwgBcwBoiNqvwf98HnFSnCYFXQ
HvWDg5/0Sn4YTpqFirN5tEnNlnh/UBlI+eQshZf7If1EWzEsMHMdhd00ti0CsBKR
F19kykosFgM4LsseBOcJ63zDpmUDBV5bTfvImvV8yW8EPyv0OulBWDeyVYse0HzH
MiYXweUwzv4naQZ+8nUXJ+Q7P9fPVfl5fVl4dqTrm/VDKpXPx2UDlQfRZQ3xJAkS
7LqyQyNjl6NCTbezj1iX6EDkiL9lj25O+FCpY6ZuwGDU8hFJbG4fVXr2ilvPhokw
LmtSzzLPlNjvnhOQXwG7X/Yy1IauHCfSQEbO4khfpEzGHbBmjOBN5IB6Cc7Y5fva
d2zyLJl6V/lBcSBPEnzTcAm4Rnrsy2w1uQrpNhtPGeKUUami8G1zfgRCMthK6/AE
378O7RG1dwYZ5YCxV8NA5M4A4PpvC9XxCpuXs4fkG/lgg7lboUwmzw916M2PLXnO
g+lo2vHetEtbUn+0I8Fo3Jbw5QK8b6w/RFPuQ3b8zvJPrwDmkSl5H4tZHU3bsI7+
Z4esLOjUK1yuwo4tgM4a5XxGohq7Zo71rWd/IceUUE3gTEF+tntlndIyx6bm9WgP
Cy/cHcdn6AtGGUBNv8n5lcwkgOcUOJHGh5PWoRDK7/Nai4bf3LJNhKqujE6sfCYT
VqTgAqZIT8UCWjHzHaD5SwKR8l+QmxPUfK89HSjoiS0EB4bLZLtLfz9wHykpPBPs
T37T4rWA1HnK/xRAUQSQSSTDaKxpkH3rRwByFOqTKWX2yQrMdUjgswQYlSZwU1w/
ehc3yq8HHnD0qU+m3AYAWFNDQclKr1i8lH6Z95wBwsterzJxY5FSpf2Qlj/jPm3E
pI1SwvACHhNOVgNs7sj1SvYom4ydLWUkreRcA3DPX+Zrmh+dJ69hmF5HL8qj/rze
bE4YeP2FKbCgOm+nbBXdmKIaeh53AX1hg3XkTdWLpGOQVvyTt5da8RABg13kVfGN
nltmUj1bN7qffbJBzEHbhkIlGUpQW47qmg5DyK0bNuJTQ3T8m2lh0cXTIjEGbeHg
CZk1ePtmIBJ9UOFy06zKBiGaap1+K5weG4HEhyh+YoJlTGqTfJ+mZ0i9XfGAKD9W
ZAgFCRqSgBlLIblVpU7WZFumJRRqXqXilmSINUoI01ziF7DxrWOTaVEYysKgzaB+
hAlgnjczBgmSeE8SrjoV0QO3fKLmm7to6/0g1WSrTN3RcD/kFv1kiRfzP7VC3zWV
ku32l2qLIoBi2ojE7lfL7FYvwGYOUZ5k+vvmSmV5RmK5MieXH7TRYq3gsJFJ4HAl
Lz7XPNGFR+AI/uddBeA3AmvSd/Narb/BB3u2TVxiGkMcAlY3iJrMiTznbsXJW/kR
UtBkMuFh10lmuKhN4gKURisLIea9QCIq4ul049oFCwgFuCPj8HV5cXKCPDdOxvN5
NccxCkaYfd5EcdNqgG4BP6WKppYNS5B/sHumrvIRbSHiKicWiTwzxb8w25yBY+ec
66gFYGFZK7pd1LPSGYS4uHCGNpPizvW+3ouOUbOLjkvunLtWakdPqTUBt+SxJ4XT
8GGJ4/IfCFjb+ay7M9+WaBonJEZJ6qGKkK99u6ETepD7BbgxI2YqNK6+wha3Ixi8
IdxUqx76lTDDFkdBCzbExNOKQyMoC5dH9BQyeARk8JV8k/Ah/RKdKLbIC7GIuJS3
wyXV1/u92A33cYejg7q9ZpZ6bL0u6LGSzw/e8ROUXKtoNLIGuVBwS+dOWxJpuagJ
Lw1nQNScGm+e5PWFCPj/kLH9XbJrKuKzMezMQHyscCIU14+QLkeg+P1Hw48cyr92
o3sRJQ2WcQotNdlRKzQ0sV0TWGuG+xSYJTnkH0jj1ApjLdEZCLudB80WfmuU6KlP
aIlyEbXUKlqv7UNyX95ThEAPCP3LvzQDsH5EA3snYiJ/PbXJJiZMDQ/SCubRLfqa
U6yZmlIkwqdqVoTnr5yYOPFajkcm7q0lsr2YR+2heYggwmDYGQ0+LPRMtlVhRWSQ
YvWvI8cpkw9UP3OCGZ5+w08WJaUnktjUhmG3XOA3MmB6ckkSqrNrrN5+DtBUs5uL
8bhzMacS66m9meV2fhA0CpW3rD/+uFIxfVg2Cqo81lyNPPetFIYRsNQ5L1luNl3E
weK5E7JbdY7Nma3/JqU+ALKhezL4Ugv7t1OBlLdDJ88UvB7ROTFcqEl35Gt1ZkoQ
jlZLtRXkCiSyux2TraTkmuVQQ9/a5Z4ACjTrMf8TPexDiNoW2IzcGsxzUjjBErs5
6VjHuN9XoljJWjBxZDPFZfJgJXlk004Czp+03IDrE/Tm5amVp3uBFyZfiWIbo073
2W5dcTIGkkBBBX5a/FzISvLBWGtsmrNP513Z5BtgQBnhwAJ9EFr9X2kjeo/T30CW
v/CcEFCs+I9C1Ru9K33yBWLKZzTqft5VyxzG9PWagUiRv4Otp7JO7TpU8e7V8Jy/
yv5MFLHQiSgzMTYr4Sw9Dv66FbYTptFkw4PdsgpSF8t1f1heYwXmmqwNiwY+9Rxb
ow3jHaD4oA8gC/JXphXcq3uz/VHCoH9yKgYzvx/LvESaWTe+3VYoL5NppS4o8qWy
iw7mx0lsktFcGs6RVUivmL/x+fkw6lcEu5wIrH8Pp1qHAVtxL3jUtVSkYeN65YM3
k6pz4v2d8BA0QXho+QJSueROfrDtmu5PQmMuoPaK/IW1ajLR9F/EHdyJDETZB4or
klx6UU+UxsS0jHQWnUBlsMzyxaMqVOQgg5qDISIEA/y7+Hv/nCCIZfZvIdX0T0GF
J9/+TXVUWw/Ha8lUB8QcMLigS1o+6YP6AhK/dkc5MHB/G6+Ly7fddKVDttJxGbEQ
J/m5Ua6P3TjntCkkILzxq7Ko4Gj0UjThLH8snTraNg8SkRtmkCxOaCgNFXz9GRfD
7apvWXNHWdXCFNjKxPcKMdVAYSFu78oWl0eTlWDRbu1UtTePprUNa/idFkcmNOeM
fE4ENQi7+pLNxLNrhnlKXjAqg+IEienSHrCYrp/RCg168F/yQlo1RGCajGnuKtk+
jed80jevz8f+yPg3VZSmMeakB8pFRxQZLPI7upWSUanp5XdPTbmQ+HE9yB0l4ZMs
LVAv7KzARLjXRxGUBu0MAhsjlH5WGAlEaXnUsGPvoJzFovjWH6+m6oAAYcj8A5lV
KJ2OMsMS3c+tSSBH0UWtY/QTYgTiPoWx6P49CgcpxkuDrK87GXQJGEtr5dK8cD1s
jJDVagcff43HI5Jgk2kqYsW0BSm6lqBaG8a5RTCmFtNTTwtrKpuqTWn6efesLuep
wYwiVWjQhKiBFrBMOUFq/Rt/OxD6OOknzpXxITqBy1e5Ap+5ece6Nbv77KzgK6iQ
qQYLr6sFW/brnNT7SDi5DrnfH0Q8GMxdX/qT4sic7MpIA/EoN/tq4yJBMX01eh4y
NRMu3U11rIXB82jrhnykg8tnO0aoCH/cmy4fBKQEZo8kttfvpLgnC1IbIR6yD963
nW+ADAzmvXVeeq2jdOjmBMOuvxw69/av+riniAHkbSqXeu1kVE1KOHu5ZWyxj1X+
gaZydqybbAYzkgCr2HKpgovPDeXuzlRe3dXDfzU/5SaxRl+f++td/sLdfXIC+XEH
9Ew8TKhCktY78VoH1jaDqRh2ag86qCfTYyFOAcYPrBDGwzL6nd5EzLXt/6SefRk+
AWGebiC0hPw9cyIfIW7c7JewRoEt8W4cGWH39/o95dQM5HvBsj6e17ors2xH7y+N
tf7jKwFFzX5gR5I0x9TdzcWv7IgxhKY60hnx/h7kiUK0EPwL18vtK8/8Qb8TH9Do
MI5XaDX00rIToW+jLTj87AkfSN4TCAZ+71XXLGbIyqt/50X3VRwNqGZykvjtjdEX
jNfKSTNxTTpKN2EDj0qsXqtvj1kj/RcZ6IE7bRkOaMXlwng7cLyFkIc2CoR2oLpk
oePNBpNWV2ezE22miYfzDNAzzHd/n1/nqlONKbDrANPOHDkxAJGsfB7SWlnqo+xt
1ktFjzfibaTfzNa8+lQZEZhjOI7dxj95F7t1p6MUR6E02goZbDdeWy8KwYFQ8YWU
MpbcB/cbqBIk6mPUsDR4ZZPll+efmEF2g3g/1/mlIm2IUsoaJZjxB67WHohga33s
wMb3LBNct/a+qS8Ecd7kJmV5vR9Pcv0cHSvMSEc/33PYKNggekTmsD2gyUKmP/7G
hU07Dqcu3tj6/aWCN0z33Pxm9BVWsXATgsNT2f8iHkiobv0BP/xzLcQ6sFIlC6Mm
QVtriZ70YSDCCHq0Jp6exyeZ7nwU9Uy4tQxlHTCRqjx/tJceY6cx2XZDjaF38lhj
5Zy8K5nGhiqiQVdRBnD9D/8s4wtxVq9vsjJH8fIqC4Ia5PUAZP7d7iEzmJd5z5sY
hzgj3ubWHaG1e2JobXsSXc9AFZiY4hSXv3XuZEVYJYpQfHziQhwUxG4rUqF393tb
j3WFgPO36nRz2vEGMNKZcqfa6OEuoFPLSZPaQK878LgodeCpgAVigQKBDAGArgTa
vp/rORfH/bHxIiatzVROP611rCygaEfrF8amYz7Z71vdDY8gchKGt7hTCY25Qse2
LuysPyhh4jFj5zh0j6yCP8c7gKKfx/HEcvtwNKkopL2tq8bFViU7gaOdnitaXY6R
eY50uiU2HglxNeWhZrINoin/yopefl/+90kz4CTOmIIN67dGkKOC/RI+lJOrlUpU
SPMAzCx8Llq5BpcaLxtVyaoaUoEjQ6SZyMXirW8Xpay5PmIyC8ZQYoS6kLxwcfDr
ZUxHO1OvRS1sRcc7dHpbfecY/3NX4LLX1QRcUIbnXthNZ/rhMBfJjlhj9yEynJry
+rssRQNPkt554K2oXulJ96wSLcESIwHY30XLzkfVf/UU47PEmRu2jTOjw/0hjWSy
W1doClndLEi3EmjQQK1q7oI0eYij4hVXTWOevATndL9oFmQ4V/2+fe6nUZ7uu+0L
fQdRChtSsT8A8alyJPDCpocIghbgSlmKLqx7TcrqqAD6OIScHLWith5EnJy1CNyq
f1oK0nhpe+DTfoDxCU9IJOljq3aGYsSiIe18ja+7HDmT0gc6xoI4tRslu/YJCjLj
XH91B1MfIQd60GIJTLx35t9kFspOKrxduOA7Uim0/udMHogw+di6rhJ0yNNyO4e7
F7RNdaZTNMdV2P7XJ6ylkhabVnPulIX1qqqPjFysxPb1doExMAL/9Lg7nNELrZaU
aLabk1MywLs061i/FS/T6Dlf7sE9COGV0a2Y2n67x38Qw4kQQi2qmXHVguY07AV0
N6OvRl7f+hblj2UvKIVlBtBS8PfOQqMe8NixC+hBYl2aYFUEoRVR0unEXrj+U/ps
ssRmZYCO92VhwiS1DeuldhCrdYLpv1YTQu5WZ/nysxVRZ6tdZse3KHDjlRDkY7tC
JkWL56Y6RlwumuVjWjnGRu7Q8tnUHp2gCOyFiUTKkdy47hsVZ8jGpE7Tb8m/JAul
P7LktAZ+xENYg0YAlJj/d8hioGg+yMa+5uzBzV7uWkVcu0dpq7OC/yD+38bXv2Gi
hdwVNxzaQdPNeAueeDJym0baRyNWnXh2OCqsK40ILWAA9Snw0sFCYF7or/cYsDB5
cxx7nARXfBZFzaIgrW+jvuzkxpJz9LpPwiy15JJb3hN+fSUO2IA8wUev0tJz0E/e
06Z/iiI27ksRXnSK3Iw3DKgcWcNkd6qDA3ecXNl2prnFya6nBkV3bDmlfh4rqDnf
Bb/ihmEArTcmkWVZe4GH6nvwO9q+HR/o4clxFspqex1gmbaiSWB3aSaNxGCCd0c0
F+yOlZWMsjirxfn63pxBP1lcSHg/7kyYHCE07m3PGTycaX8KowGKSiFthRVgVSZ3
diH+NwtIFO3oSJ149eWkLd+pjvyblQh9Hcejstj4QSB/OhT/088nVTvXujyuHDEn
n0fbQ0YBM1l6UHv1jqnj4WFSN76/OrLXQ3Z3E7CxdXkq6Mk5MVfRCqxhOWQDKRiQ
iCQ54hWDFl3yD6bsOzAyD/5npl3Mc5CTRIzJwRY6TW0LtRsHkPmpkT/LGIihROWt
f9llyEPeA+QpxiKzwKaHfBRdK3bedh52PwxvRG5heA2G8Gf60gLWEQpXrPldtRbD
O2Al7wEwr7wSqdyZHJu0u/HVngSrEMuTZ3zaYw1bj6vtK5bzZQfERfHlMuZ2bpaT
8vIxVZV9fNAXOg57NgwtrEUX+9AMj3qh5tP9SDsrnNPNRg3/eyR2ljvZ4IyiTOVl
cDF04YEq9VZZjQLLOTjvwEqiTus6EdLAs2x/GHWehelaWotsokb3s5pram9VxzRg
CAxxDW4VwhhF5qJ3AKNhMuFqXlfMGz/LF1ks3cwYFEixZ5TZjnUWrxXGfpuZyu0J
Aqp6/roMEZQOwoJwarjSmcI38YcSjB6JQEDgdYvUNNqZwkdNX1uJOB/UmjymXVUc
dESEGqCrQtcfhSckwUwqoa/lhD3aN6CEnEmm7Kn70fvvixQ5REUCS+rJ7CeADzlS
BF/DC3eG2rx2iCZOELxKPSY5CdSjZ1GpyW7lSiRiO0wVFSyGmFpuTIwuTST0/2Y3
EN1apx5CDV7RQutzKYyfyT+A/g/ive0nV+d6VMRSgykLau7b0dT8dM1yRGB8+Bla
LoioWZdJwdb506gAjOOp8dE78koOjWU2YXsVV4TdRmiR74w/RxO1jI9ifVWg+V3U
xvX47aWlzTJC244YeK2WNKAYjGemywxZ5zIHVGI0+tpT08XxAmFRH4jg/PgCvS8G
Yd+dGXl4Bs55e8SHXrOQ2f+Aw/eaPxZxnr8wIc/3VQQli2x7ehM8XJ3PeErZ6g5R
bpdP5WZ0BI9ZxyKulwoi2xz4hpzJ/KNy6lTS1MR15CgsZzVbG68jBijbAnV68RB6
yH/t5datOMtMMv9f+RUGHJlpMTCRY3QzFvPz6Ax78W35Vm95xn2+gwi/yA2ykgl8
Wk0Z8x9FKy9uz5BjGPnfxsuhUCLPhlsynZvPL+Z6LqxLYzTclw/Z8jymRZJYR6/U
xQLn5UtqMjHYExWl+D9lcJC02RGTQhpWEWMu2N4tPgIYjBGRQIIgYfnBoGLY9Up2
GVm/EztxlzQG2ESUQuba1ZcWQsZ+5XrXUlm6AEV7Wqa5UYhWeno3oG+ITVCWH6Vg
ZwJChzjfxaxw+wI0+MAY6aWPKzzADHvDMUPpmWw1hyfp4HcOuCk/TlhmA8u9hL6X
/Vws40dc3CqD24BU3sbMNpd87j3ePKNzgaBqHGVq9o0QPvGcBlye9tHt7rpEi8NT
PQrmARTFBLPYLx9tpuIgmxvL6KpGwNTVyKX3YCLMCeqnP1mjZR4niD7jAVMSIJiM
N1fZ73KXI8DlZIHq2NKrWNUj8c1Y/Oxnw4WzXVvqHer15S4GG9kG7rmhpFAHF5fW
q1a5hcR6c87EhFhbPjEscUJBdNqjS8+6AowEjQkILNYidsTPEstSijq1rhu/hOor
4eJ6OLIIorOU2LBFPjCXm6n2rO9Yqe2CvOodWRBqyotQC6D6mz2dM8VXZsbKShw9
k8iOYh3rcLVSHAvErpneDRTuh8pV22GOwY9FrrcKJXWP8uQKVPsoAyn7Jc5UuAvT
yZJGAnIGUPBIVqH23qEvf9eVCkyEVtO4FRGBzWWFceYF5Xr0JnHIVNdM80iIV7B0
NAJV6bzxKI0kSn0K26msgJyzCqPUqqAKpCXVoXnV5MuCbU5PA/vGNysMs8Y4j3+a
cKXlAhQjcoXPw1s2KJCvIIxsamTJL7HtUvdRhwogdCLouR/Ut3QowEEsENuJvx7J
XVq2mykCKNMKBiGnmfGoEIuAtzCZAPN3B+ucKNOlDkVZjcgesnCJuv+kBzngJp1E
Xs7C4UxmZQh2a2C0oruCfoqv7Ywhb6evCFzhCiteKQDaEwAHujLbngxWbzoJaoSS
7RWNuJmh0wO2/AJKcF3oJBqczOhpmH7j1HDsUEBzFwo7CwLN/qi4ofD1M5J4MfOV
ZLr2cRjU09k8BTWA7aayAP9XULZrFD7Q4NdS4Yf5XeUWLiTQvZGV1RSHR1aWDXfx
FvMTTM4CIJXv3IDirWa9X0A4wlDp3/5kpvN49vv6l/K6xV84YjPqJxY8p6XJkiTA
wZI3Tg5Tw9QUoCUpzp9f1yW4DWORdahmmTfFbLKckU+hsghvddjvyMJOVuBjVbb3
YD4LPnNM7aHWNYEZTHGfYSp+HY5JYrJ62gLWElFmrFg2yqEKKYf6GyqP5LUIH6W5
EWc3uX+B0ufmYjRURgxyIY1l00KDzzD6RmAL615rQbB2d6FmQFbsTcnhXybFsxqh
tl+RtYe689LMFOeqEU44sCfadD5Wu/MwyE3CrLYS0sShDELKm6OmPpmIuZVHiXos
KfvFqKmmgjEpSNkEQoGNLHcJvN5tGYAsFFCdCvKTLUfidv6XaSBN+vGSTaeEzVdh
bb0dvlF8DVfAnQeAA3EFnl+JF3kksflconbN66KiIWgUyOL6U6qaB9wzBPfHGDcl
k6kKrX6LCpP4Se7uqgt33uO3/YACeKDMVNylG15tQ1zlPBh2cqhcgMy4jB1IFBzd
kI6N6PmcRctzarPxTci802cNUlakJuEsJNfXaQ6uc2GCXv29b8GKGl02tQGPPCVI
VFma+fdH/bibRMfzK6jPnVTarzfh+TqUurwpDCNr7nOLiShP9o3rqKsS3CuaLFKH
n6iKh4mkRn7wlygwV50xRfZezcRM9eyF//gFSC9PjXjfDDj8ICMA9pVguL8s9m/E
RCDvz4Stv1aq+7JYMvVqvPkq4Wo5loTUX2SJGRYgzlcRGt3BNaHX0rPnCpaHBc2e
yVRPHQHW3NHNTcMTICIrh+79EUjm2cpDFFM3hi9Rt3bJfim5IQOh5sxE8xNJ0A57
y6m89/ek9JVSRIrzB4c3CwgIfE0eg/FcRLyMidfT9+VqLfik9aRC5hxrIpjFG5sM
Tcf6m6+bVIb2IYheiWfa32n8LOrGaLj31e4FXtqnW/H953bFRtDfGnc0M+oOSTdU
vG5MSPdY4C415Of5D7K0CF+lm5BItg6AGOoj28DiClkkg271SlHFfhu+SV060wcs
6wWgr3FvncwtS37vSnR6jzfznbmFDcWAWE+YdmfP2xi7Zsw+vCyyPgE03K61S3AQ
YR/QLw//z9a/mpEPp3dVuzoZCHn0H9I0vxzUxMQHvpMb14+eWQjT0Vu0E/6A9dE6
TowzLFAz+AtZjf/7cp14NPbKdCcpe7pz+fcxpAI1ay/o/Ajj9JPoLFMxHSaf+4gr
0FkWZMl46qwXPFcg99uZV6PYG+5mS0pb4IbNt/2HjLIExDil8jqCYpeld6mPIpcq
1UK+CCRIdZibmeHFMvcsJYi4EoCRdZfb9IyRNeorV7RXTWn6lH3K9Yol1jEKUu+N
3ZTrWwyQCwZ8kzcNQHaus/b8hVduHL9qGCb73sv4gR9QBXkJJsC2Rf0djw45q1mj
c0SBUvxaQQmuINjRvDo5WSwt2kp86mb1fXDlHaQDpWu8CN+efsRGhDTBcbg1h8X0
Mkb8lo6Qs3nrdvpmstaWforhXVSaAIRgjY8KbeAaUNYiHBQR1c7AKlwHvJ/Kp1IM
cQl2at5lmFaG64WzTyYV0QRqdEvhfQfsNo0gWO8EBLKxhE8dCEl0Xb6fISZUOzT3
anR2fz3CGma60CrYx1efJKjakFXzcnmApH2/BaH7o1Hj79+5wXXaio3pEgZKUprw
xADES9p1pdBJMmfoK6uwl85mvy+32XSLhSN8DsjW/JfnEniJbCVLXqlBYMChYCVW
Vhb+fOlx122u2Njvd6nR3pkV7ZpJ9OBX68dWnPDs4xz/sD9ycgV+dVXXJ8uoPmVN
gmXEIZ/uM6GevoS+i4kQB1++jGJDn/oH4rj/9je4Lb+Q9vYDkItxTpve9Cd7J056
fogQlznkMK7x8BxCveDW4L2LvwSighBEi5ms5TYyXWqNl1Lf2aB4XZbEI6cpaNDH
i92hNHdVa/puSTvAnVje4CL10xj4fvYqCLYi785+iJVh/TqFPrG76M7hKCNJaqhJ
f1tHIC5q7ONNJJAeCU6H7jN1KUhrK2YoC07mWEyrAUjBJfbgJXokAbQhzQpETOvG
ANgDnRLRniWrpZlrXl5pZoSskk8uzYe8KqpOHgmXCMM0o1U5EuJ24FaADrSFEWnV
6zcpPwePWr0MpKA1w+JMJN6yBKi2+lebFXRi+3V5wVHBD3lmGKwFsCiWQgcQzEnS
aFG4jyRVk2iuZE4HK3NxSlsO7+dVyl1tDy4WL72K4ojWgzs42MS4X0iSRJncfk+I
o65cCrckasMaunB0zWYWSyeGz8in9/YuW2amFi1GJfVoZ7oMYH9ds0nr/V7rYmT6
JOr1oldFp99i+4ljJmaQqHPsPueDAu7LqXsTIu8ToMFYikQAH9E3T0yxH0/aF7oZ
f25j7+adY5D/l9Hd3KTMYrfLfye1y6BnKdOT2hSNTSUlViQ/leTT/BDeOiuZL79d
Lk3RXSw0rkkrEjk3G4sOKs0kHFll8XBbE5Tyz8jI81NLJOPWtxnpbLW6+lewdPg7
7pcolW7K6RzdgEcmH1iwWGmSQCYyleZcuGCFZcmxo913QEpAr2SWGqx7d3O0PO+O
IQXqbSj3cGTSx5zbgLx5VlXt9cWsrHlmDgAjpWIZ+cc48Du37riM9TJ9EOSeRtGB
QiNq/oiKpKzzf3av1K1BrG841/jp0dCzPbNa1VkhpcvaghO+r1ne+nUCWzYP3gw2
VG+JX8KKCjdxnUJlaoxeDzF3vWZZ76nHizupfohHrQCgXbb6tp60YArnwHp55ouQ
NZgF1CvUgYod+nwyPliNyX4BqrqjCj9bPOpXFdlMUSy1G7RZt/hgGA3Vbc4eZizM
DacZ/mbuXxwY0LD0i5Yhkc4t1xoGjHspO73jDCala6aaD0j34Wt2oJ4ozgvV3yyP
ZhKH7GTevY19AoywuzDvgT33vZKNu7tEwp6El7oFB1ymdwP4944GfsBf5hOrClQx
wT/dFKlO2gNoMjw8AcTHzKHXGPV7Ha/W5Kk/vc4KzFXtpJ2qLNUDobX/mL6NsJe9
GaPEq5BO2sZl9q6PUJR974Wy3VTA5DuoMjqXOCJ7Vx8eABK0FY3dHY8G05wypRrK
ZW11Q9h6IHpq2Fyl71H6K+oGzRX5Y0tVBJ4785VwuLbz0J/nzOXRP+OsuPAO5lzL
wX4WH/X1aFxtVsVvXaTFnH3rZ+F+pRW3+BHMzz01Fmp//2lOTxN9F1PM7E4o1Pu5
Zosp0O+n+AKa7uENuiLkk2Uxu7vxDGkIdMpteomtAsp3GKF+Gw9cb9XKEKboS3Sy
268ox3Js65NxZ81l9Y7Tgxn5tL3jmQOeUp7tKccRvgi3zmJT5ymZyt8co51mHSJP
iTPIO9Up5+xRYmzx+SrGUf3f1+xx3RgbVRvpZ7bOpBkrbQ280kbOGQmwg4aCu3HI
fuDxF8WIG6glI33dmYkT7OgZ/BMg9t4QWTtiMFxOZW/XvVbCvWOrMIiTMEdR29nT
5JdpCLo+77l8sGs1c1Mx++C9I1iZk6PaPs+eJOMRVk/miymrHCaYBeLJihX7C2p8
xdwcGpfpuKye2gCWu0kSLI7p8RgDpZmasIzj2zX6K/1AQbfLuCYrRlFd7Wl1hTBl
c/4/Hxvfzjs3WaPiQmqf/6c7PhFbNQGYgXX6EGkEMFiuegZ3Jqrccf0EEa85/8XL
01egA+ao/fwXf1ZG8CykpVkxgwYArWy0zBF2P/UHBgPdXNtqJZdvdfawE3+7OUye
hTd6U/jHow3ScWveywkineDLCz3oH2Qs41j+vAumPbi6N56nwY3L2hMteMeuIywD
t5KFx5egispvnzLY+3716gK1V4vFh7OJHR62/sJsZPJ+JiuN4TEJPqhmMNMQ/vIR
2qbQku8Bj72UxJYcdJt1hYlX/k89qSFKuBExjNC3K0IcNjLHeQ3OlhvroRsvrkuY
WsICBKm7VLLxcB18YUxWvbZsJg0Z4SB6aytwHEISal5YiD/UnieH2liBRWGmtc25
/XVOmQHnnBADwh4nJDKJ69QkWv/owdK6H5r1WiCG8MuFtApDm7b0RxRzO4LHdHeK
ctiC1xSsaRZeZrcMDFdSTuq91hWnegK7NHrwRMPvW2/eTnvMC921NhYB7LUvjSnD
WOHKYVM35SMgmORMwJjUfKPZ6hdk9ZbOHmAgzfa784Mg7vJwRII0bfm0+UGxZ9x3
26v1Pi4ia69Ke5gx3gbfXq81hJKKyOvLQyv9V7iKi8aAD+fPadG91J2OQ/ye3oQt
F8AgtuqypaeD2dtz+M5oI6xvamDpWr6g2j1ZQVEu3fg8/9KHXS3guggCGxUpNQ6D
1ZEj+ATwuCTV+i2A5oOJmJbqJOvvHoNns1pu/l390qmjcR93YyrjZvjguAEfuxaR
YR6IQ8UgfVs4l5aJud7v5CNlrf9tcxinC7KSSDYgUlK2zUJ3guz2R/yJbznkD5bP
VcbXxP9vGDT4/VsqEP+UE/tEjfJg+x/iaAeyruRPjNoVAzvtzh7fTtrldNOIN3g1
m+NFeKtKsHGtCRutFixCsr9yFfBRB/4gY5rYVwJRdL9SU1WqBDkLIMgRySUCSXxl
WB2CgqxojhTcAOk+zARkNUsTmPfjTc7O25nuZ9FvD3s9aPPfHwihybuxVRPHLwnn
/W686OoRgfPYur4mWkfxE4I4rgVbyWYIXAYncoDwWwujl5kou5GjUpsx8/bfFFXp
FzQRo1ONGwf16l2aL4ieB64eMLNvyNEV1BPbMNo9N6qDK0XmyRVXEbVirSJrzcnL
xcEJA8mJKT6bD5AdgZYlvAfe5SurJAiqd0GjFnz+MLFxfzX2/9ZVLIg0ObJ+uRBB
LRNcZ1Prrxw9TOMj32ta0w9Gs/h09Ka1NYgosQ+Y2hUBLAxaMyIgFx/Ebf0qhY2o
HDMsm7pRua5HhC5PXHiYrl1MT4USilOnIV8qYFtUQHqbcz8FAJRk7T8ClEUhJirc
Lr7NT3JRlgGDms5anffxeMhgxD8Nc8fRQX2Me+SkusnZn9fK2TjoDFbdkJ5mNftf
t0dJBiE1+h3BNtZ+pPSgf2Dz2Zkg0647JIOxKPDByN/u/q+Gm7U32fZGy/fhgJQM
CMqVmzfk1oXvg0HsH/eCuFEbfiuTkmhPdqYnaQGjL6gNOvf7xuDCwE9pSYpX+SoS
YhWeU/dNcNWBrjQoXcrll9VZ5iRojjISfC13oMzmrsBwA8QkuL51UkMUcqcsKA3S
CPAyg5033de1GORIzErl4vr05yRR30woodEDMtckJyOqCfw+VG2pTBHgPrHLcm+q
F4gGB3jIqk79heXRbVLhogufAb6vL2Y8Ao+8SvKqFSVs04K5wehyuLiVPHFvb5Ni
aw3TzcK22d1V1p/O3a7H1HS8iiqs9k1PaFunvh1OWCshlLDk/qOobLb/prixkH6x
WAWsD9R6yNLW3BhnBmfHzTOhjGKjP3j6vSWJcvMcwZd14a8hIrODmEqqM5ZHClZa
Ms9c1vkZjaxJmUHWGxMHwhO6sFCCKJpsQVwRRDhc/2NUEW8pr7gU6Rx0RAk3EylH
zVLKySKhebargnt4KTywNW9jx4wyViUTAg6sGsKub8nUkV+7eRF2jQK/XsDzQyDN
Vxdh/iuy173QC6bArn5q5g4V0sYqyDlFQu2XIxXMZxbRqHIb1L/k19IE3rlkNY7Z
Q7nRy5fAoQodj55FDuTsYqV2GmyvMbIR1FB8MDxiy3NGGyaQ9OBOwCNSj2SMKZUu
ih6WxSFvyE8WpOpmP8C4pqR2bz1UJzzjcG2fkA0ml8ZrWSnF1TUIKFlEOJdRmR0S
8HcINW6ZUSL39G90pQEuQuQt0GsUlnI4zg5Fu55+Hh/NIVtFmXekORjpxbp693aH
PMbsfmF/CkIJrJS1sFc3k9o+IZzQpoH2lAYubxLc5WslyzqsNM3z1yw1b320WuUc
Ujd14s+Hsvw+2U/RIfmkKQL039X2aIFdmIIIJWWTAJpvARER6TtzwaJgLqQMKfLA
y4Z8ZHZV4xLJCmXxuOLrvHCl3VchIrORwq/G0iOXVgo8mnDv8b+bhnJkYN7MbP6p
H8Iy0moiOLMCZ60tcu+3yRshD0xU+fAIcX+jSIQE43Hfl4OhYW5z9W2TGbiP8eDC
GCxD2ZWqUrb0fvAjLhPRx/OTotw7WsngVqLGqX5jVpZX9vG4ZDvBmqH/1/i/6UQ2
ogiY7ybfCWj0eGSUU/egxifz+0i0hDMU4j42dPIbA4YPxqX56y46JFiV2MrRRUtq
1y1X+KS+hPreWmT9+Z18EGodol44SXoHr21JNtyNli0npimjXjTdez7HYDo1jeqH
yjTKwuuV0h4oyB7X52XNttspLL/ntB5nxZcT773HU+VGpqTyx9zY/U70KXTyMt/b
Khq7CMowLRn5TKqy6dQ22xw8VW3Vgt/RKjbqQcF8Esi6WN5nnKOdX6/CijUGb9XQ
g1r14TsnA1YdU8lC6dZf7jr7BX/yzysfB8iSXTRlAxHPkuEYiiRn0601mmIgTNdM
afoSvll9sefLJbi2y6dqogmSbEFCz8TGUIZ5D5uVGBQvlUadJJIkqU13s+r02RSt
8BWz+wnT16zPHiq0Y0FBT0QYPa9GgCfUGyrA6TTJDEeitFHN76qvC514P9BmhcA9
uUbflRq2rdlg6IJMU109SL3kKocWc/e1bejkmQ/SFBwk4CWKa1Ult3MKpI0iFRJM
5pA68i7Jr1KXnrhvM0FS7GXrnFMnW8MVJ7cVaGyRJndWomlY0j8pa2Ll9tK0rvt2
C9vR43E8KyZxWAjVaIUDsIw7UBvY201bR5LqujQVgKBvSa5qfYQR8npm8aSf9nKz
/yfUpbobaDxMkljyKJwPi/CuJ0e3FS0Vg4G1lA2364t5VcCAn6KDcg8LuFwfy3mF
r72mmfdr0PZwGkIeXrXYXxwbDy2LfBBFkVcsAjk99JhsvZpciN1S2A5QWChmXepE
Ay2SxHxepZvX7K2AsVBJqOCnbQ7f3Vi2ZxVUg6+KBZVwR6X4qp97XDn6urfNJTU2
Cu0ivivXsAJHL3jWKLyGPB+FycVL9ZvhPwQBaTtG6aOa4EszyUyP+CWtt1W3tmLw
tNrcJBdCb0U4+IuLs92DNy0U8T88SQa1/Je6lTfkEBwwzJA3QbEPuPCxgEnou7Xd
3ROSNcpkN3H+vAomiTr8MesKBsqosJwiL7uYcJso/iKdnSwM5K13tG7w6msi3+IL
EQ7uG6yhhKjiGMr3xHI835rh9ubrnJ8VQp0CaD9NK5sD3MxTY3cXi8IwRFP7c3mX
UaQw1jBbnGz0IFAgZQ9t1V2+t8oIViN/+KFRQV4PWEvjUPF46aPUd5F0xCdgrUkM
qmbaHo/zq0vWESatBd2SEMJ0vdZnHOD0tFc5IBt+vdRJBOQ6b2qlvO5enAgQRJTd
U5en5oeHvJUHaniWrEIsx+3NC5abURZQLxi2fHNsgU53YJkGKFX54Gy4nvT5Ho/L
v2BoTX54xClQdgCTb9gOKmQGGk4EUhC9eBozdmx67HqkyjL/7bYQGOmOaNEUOIka
e6IRhQkS/dwQklqd1lqcmha7VPC716kGXD7cE31oTk44+SEPIBMURSa7jzI5s1pi
c7uRUt2GwgRtRkxKRKR+f3bhjnRH17P7DTvLc2NBBRbrt6c97pbGQCsxw72RqKHG
aKp/ZjkiE0Rdwv17k6MFQ2HtIcaQlXCJy/uvk8S4TV8t0p39oUkV9KJAqNP/CUtu
R9HMmKwLPpDwkY21Qf8PF2qfwMIW8t7H+sJXpOqeEcDzTrBFRRjeLqq4z61eaXRV
Gt5+pSYk+9lw+7c3b0m6EQB5lO9Jz/WLqVSQtdaiKDzpC5iQUA8Ib20P7sJQr5N+
vI897UKI57++SrEdQMf8z55wF0KB4f6NY4HtBXbGoIE5Rr3mNhxcIrgDwb/AuBgu
K28XukEpx1Pai+ZpB8p7VpbxXVw/c/rk0e4+e43LI16Hs00gofN5711v7R5VGBZN
k4CLQjT5yFhkuliGg/IUd/M3DfnDzMxfd0LQNiEGCoI3rwFYH8L0dNcewraeQTY8
IZH1A/4WKfnhg34/Lo/7HhVfIrC07J5n/X5aQvkzgshFySq507WReDDX3tP3Nq4L
i4nVPJwR4YtdoIWO0+kjOygwIAqYQUmh/V0TVnzEYaESXVPXlBRXH6lvAeqsVlcP
aAdJArpANb1Ql6vOTegHavxTorEErWXPdCMsnnTTR+QSiKFv6xyEO85yzkVKdlZF
EmXfWN7iV2GVrNvqw2PsAjrIb4kZ2shf7tpm3yB8iM+q+vxC/kvvwbgEARz2PDSg
RCZ7fQqPUxpDP92h+63G8nseNmqSDOc8w9zCc6hJWp+9nfkZPaYIkUf8d2l5kuUC
UAk+QAgPFNrQuvRZVNXEQt0UUZwKdfHr4korwYw4IpEzb4M34AlzbKUz5R7W04Ul
unCWdQCT4/Lr+Ek9EPE4MT0NYY3KysBPwM504EWV6mUKGtTOvocl4Wr+NhJdAm9s
VxNDgREGllOGfjfxILca7HuBKg5ZeYhsCjno+2RCl9hhM7F9XIDHFe1n+wxV4zR2
KsCYp1YofYvyfi1uNK/coHZRnTAFvPpiF/RoWXqAPX8RqUW/37/dRghVjKgSKJpu
RFyi0E3U94luq1bvFwCevW1WZTSrllWvi4GA/RRoWWHobmbL00EwAFFpQUmwdSiN
gSjMLP7+kkBs2zFOwLXKFl6OK80kMb0j8BQtJ1vBJpDKbEUgew/m5WgLM3DvWGJx
DGYFTAWOPmTBD+8bt4AmdFKEpQkZoKFuMsE9aH8Cz5nd+8eo3osOY8A2kxaXWpBN
7FLHOuZqwg0uI3NlbQI6oJ4HnlIHzc4JQoDfQkHbPyPeNqY8ZpLMIrHhKuLo/rBA
vBUdD8HzV3Cp5CevpMGL50bQ1HhJZC7wkF3UpXpNRFQX+fRIyksCESKCHwqClZ/k
MQWBjPAX6YC3LDHUiNbIboq974rvlufTC8qy8K9u4ODKwaZ2LeqKNOfRmsa6iMk4
QM9bBhlAx1NZBcHohMHEtMej/w7PwnXVL8d0noxXNWpeyzQ6vvqNthueoJZOFApD
NePXpQpRAXbWxdBZYqoDXwGgO+pUqPwe95IyN7Eut/ppSZ/Y8v7t+nIJS9LRs58n
0Y3gpUHokYpeUy0uvlGj2NVJUa/CFHc0cO6eTYYrpRjjtcmlHdkRmhtCJ98IGTxT
j+KIJy4rESCtKuKD7tYm5jQfM7vrCq5UCtxEtvsZzC+tyF7znzOjL6XXCVW6LK99
A+0rv8vqYFQMC7id6uKdY+BYHZAJgjBKOpj/kQj3KjGAEAusMn/0vkDs0/UDZ0FE
7PERqim7WTjf9XD5X88rtWhV95zBYAf/Ucz/iXxt7kjLt4O3E1pwh8ma2hItEmzb
9bJePz1/cPIozcBStLNU9p2cTAlX09hZqb4fd+rLsmqXq1BMRoqWDfpLkYYfd1cu
quWwWiMnUzCntpF1Q4L221rdarUeQKrGVwzjb0P3yugI7KLpjJLiasKB9d/z+KFR
jQBvMqYXNNc5/TeN2qoNn5Fq5OgBPZmXd4TXmXWM8I6Wd+Zu4m3jDsgSHTpxZHYo
j7gUO7f6A1po2jJ6XlVc+3qZWFNa+htekN0MGdinwDkYFcsAWIR9N9k+NF6In95E
Z5GMlTPF+MmOMgvoKxBmqa3GeJGuieAjECctGdJ3P6yYtHbfH6TNh28Yav4RBtiN
ArOCikVbuhegIpREe2WjlFYcG5WXCdG8ZI80nAASRNneWDI4FDskE8nuOPIDYFUZ
m4y8OKFqciaQe+UQXSdNJkBIYjoZL9i0rQvRs//uTFbHDiujTBe/p8LgJpypcrFD
d+Z8cbwFNzEOXVTH/xTfCXwffJT5WqSvoJalXDnMtp125xQ8rTTCaVgWeM9W9yL8
jLmmXhq1ASJ5eFjbwiFEbv0jhGHJvhBHIhTeUEJjSW0mnlUSiXIHKApaHHKTuqpV
77LqYsGUIhdE6b73qiu1qOgeF2YLWzPXf18FyGYpoF4X9enc4nSyeKIUZPCNI8ny
9IoS5R7bPpKQENHZ/UFJwLx61o6UyqAxKu7krrCUsyGttWl4E8RmcUTvQxsh5dvR
9X8STXqmEl9Z7CAXpHWDnINWDVK44Wqw6zTTQpmAZEuJCPJijKgf4faQEL4ei87c
YjqzUFgpAG/SpA3ViKLQA4EbCR+1sQeod03lKIqp/2hHGiCF1zq86yCBu5fZ09qT
bIBXBxksXvi0kml3mMdti7CVspdCVDnhviLJtbMysuG+HwiN/sIJ31ljQu/xZVQz
eDhnIp0JT9fSQImE7gbV4CJvEUZiFAmGXjGzlbLmxp3pzglXk82PL0Dsv3gYf5Za
Kxj6uubi75CBysumwFcoCVVZdOZenbwYoI+VDgH1pKv3WCgrcpdprhtosV9PchGY
EQc82SLDP3FH8tD5oxehYeyGdCZhdWpcxmUbHKZ87ZV1mJ2m2kkrC6p5gt9r15BJ
g2USNHDuxBrQ2Nhi8ydpThnj93nX2JrRwT+ygrf+6cL6JtasCghO5ZwiZsUbl1i4
N/gRbpLGT7dZIcSL4Nl6CVdzVe7TRKSdG3NRwSjoSu3Mgl5FdevC5YWVbWbTqQN1
MAX5h8LbpdJpnXLCPdwhcm6+JlDqzm10cRSyrKpfVaUQIu4onEJi3Wnhonx1BzPT
kVzL57n7H4VXBDIFolYyTOap6HFNt0OEa/mevAGUUDW+WU9CZ/HcETmdapTXD2Kg
RSt7e9CiLSyI8CpQTi3Jr0fnOI5TLBO26OOA0tNpA4DtbX8qvEeqXr+C7ECzaeIC
T5JEegjgYt0ZQ7gJRsX9axu8hhDDyVIeaku7LsioKpD8gPu4AnlvPxRzpidWi1gn
rAGVFLcT7SwsbEKd6EyyvFXMudHKMZBWo963YEBV3pq89LRTeHrNXDMC1gadq9DO
kDMH+5xq0oosY7F6GQJYS4+DHHyEQ/8kSNvjk8d7n9aNFpTaxk735xQIxMudOpQ6
zn775v5j9yvGjuXR3hddbm7DaenSjOdAoVFj11WXEN15tYf8f6Z9x2vsKdGq7rt1
oJZLMdj2AnSzIEFRh82STRSsTV9Qxu5dXnaeFNYys2TLHApQL0oqkRYVX+xSuIzx
Q+QA7cLXyzalKCH7DKuEHI6VS4ysRPxljc8iqGQJX19Ax2N7L26fcQfBX85AL5gE
V1yulGWcV45lPUNiUGD+kPMqEoO40/n3zFjMXTDqznJJv9JD7b7M+/W+qT9Zebsv
HN70m3JJgN6LyKQniKZG4+Bmgi5F1mY06ybQCbRqM3T9Z2vsmisUuU55N2ovlg8k
4W6W0TGaho3tXfJ2yNao9n1aNSuXG2iGLcvuumzPfN5AhLLuiJL3DALAR/7Ws/Ye
Z2X28N9wKYScRg3tZWf71C0ImxOfKKTPkiz8/O47olyYH2XyvWKqvOONeJzixjfV
LYXRrSXF/FnePfMpw5kkVHM6td5Br56Ch5qUr8a2lYVcBeEMyzOE55yMso+/9FcH
biDqlsV3KVrdRxBCRsL/SiQYYzidUPB7I8V0yzZE73x6osNFH7lZUBnAKjaPZh9f
RqGIEDc9j2d4oTtCx77FJXYWWcQbpj7ku7/r9ZEXwgXPp/g2vJ2ak3aWjpO+qqOd
SscEuc+hIiD79oM3kykb5v6J5IjUOWTmKPkpwUiaA3TLcKHYwkLj12hw44tOH3zV
tyBocIaSqQo+thW88wLMoRbQnRcTREvxMIiRrWXTd3bJ9CU0eBjoUcs7AJIR5u9n
OOFxryQqEy1fpHMx7sGp6KwnTRc6fmxp3IOupiiG2Xm6HFR9pA8ZcLe7lkGRKUmw
kg25+nLNQ2J9ptpzHsuc/IX9Lc2I0tYLf71+z2Ho3xDAoW/KZOE8Ap7PAVt5kMha
y10QvW2TTMzP/NKpXvrg/AqM5dIHdSeuJPcutM3FvXCVhuOKY2vuBSyfPTOIF0xX
+ZtVZgV/K1l1jgiAX7KwlZe4L9vFe4+UBxugSwJwDK8hFraNlqRM2fLl5euuRZ76
qDST0cFE2FcGx/cHhBFLBDGEsIpP5tBt9CafExL4aoXJWf+kBN4NAmvIfrEzhNB8
QKQbnSitDeTOwOjRvgx6GZdUWiITRUqJEnPZ0JS6jPreoE8U3km7n20C74tUoHjr
Moux5d98NmBx0RpcL9SCrLMmN0iZ5YeYkX1gFrDcymrjKBdYgifEKokxInlxpbxO
RVmNNi9m+7Nv3i6gW6fUt17ipIWtn+Jng7w+oK1Slb6PVZidWMiLTCJANxlO4qy2
V6L4/CSmL+C1e7qASiTKyufWhX9fe0K8EUOItViiUAtS01j4oEbpsC55FJD+dLmo
/5aQ+1mCAjHH2+ez+bggVPxCSFkvkIvlINnnstl2xuAc2YQ71sdqByxFEndb9qlu
6ThmKfWqKLgRl6Kf9yeMOWTftuU8CiSRK1DR7tF3YU12Zmngv8aOthYURho4NOX3
83o4O2Z6Wv5HewHC3DdMeEGwJ3v78JsfAoZtSZ4eRThupvCAsLGrpUtZb1bTS9av
PHcmE6QJ1o3gaWxXQbyeA0wqAISNzlTz9OoCNqcepj819fMvTGQAw7ZYeNVriJ6l
2/3U2SUWx/GbvdFoFfoLIsDPrlWhl92lnSod6liV1OR2qo+bUaoRrvOxhiY5lT18
jqcq2Zs+WJ6A7vjI0bhdpg+gGCSeUlVB10NqBWn0CsS4b2DKAPxEH8FYwTkZyjMZ
6PF7Mz8AzKzrnvldp3QfN7stVP+EbYl3JvRuTDX63u+YS7AO3vHKwGqu/yztdZS3
/yHD3Imk2P05S+4mND94zqy9LtiG9eSJg3G+JOjURdvSPYTrabHnk8eaTPDzhAzu
J/7/CvPEwmnAt6pmXuOrTKNwYNcbv8eanAoGj1+9P5dz/6r4Zyq++GvboDpTfBW/
jUvO4WDBfJh3VE6BMmVOhQYFmT/MtcDgQvqE07iIg841SCHz4/PKRQS6D7wBAyfb
iAs/KXY32oQcaa0x9qKIAvrchbg8riuVnAxdrt7W9wkEjdG4hs/jZ+64iQjkAhzD
5OTMNENCY0mq6QyHzqeqdvWbWKDo5O+xb9vaYIOO3lFPPvBbtvkutFKMsAY8TwCX
GVgQ1IfyC7ZIF7joSC3j/bC0kNDzPFqGlSmn642goxhWZxG9Prkf6+fOTWVn6V3z
2f0ycoYgzFLgnx/UtcHOz4YooKkG8fkwIcvDymkNDLVGnM9CM4q98aJW0QicFWHr
Z+VprNogVmlUHRHhXmNgur8uRYOldK5ubMNl1SFd6wFgHzKbA9aZwfr3gmx8VBD+
jLfqqatbJ+qqfVydaJojYAvx6qxQ/E0o52c8WQ0EToyh7vy+m0SP6Vs6DF4XPs+r
mZcrEORElL7+MLjQz2qG+GlHY4k2dhOBSVsJ+ZzcCcHfATPTLc0cpSk+mCeCWwl6
BX4bzlCRHotj0r4LYmlJmw+orX8z7cd5XV2nsb1jvTl+BYDwvQH5MGPLzhoiu78C
FUDIJNLryDMTeawe25MHPSaDRm0gQgS9KwOmzSKBCeCIIy97H/MhUxNFjn8eLLqQ
183DG6ITK95Wp1wzIjcnOP5lWo3MhZ+klXnmZ2q5Wa5AM1G8JsWfvH5xSfzyQUYJ
Tu3Vw1sK2vqaRKaRgS+qOcgM7jT7BbXaTMROtqBqvxnfe+tY2TGAbssHHwMjsAUn
HkkYtp1g/Bu97+AI9ffO4xBrHxe5GGR1sH4havv6ETnocIKhcYgZlsWKDEF88axG
nqDRkDYGoSLco++IAMAeZ/7ERTaGgDG+eLDgSyfMTKJ7ohw+3/M7/8aMEk5lupy6
jdJsk4FpT8pQj2ELOEGHL+Q2Fmtl9RenS4uo8g8iXwtofzL2/HbaeD9LfbwA5RyV
NF44dVvlxOiLfdZL9J+F6aYoZ4n00qq219BY8TGBtq9NuZtuXNla/YCMvJXMyMoT
WBDsqdYpAiL4A8UpuJt1gXaba82IIjtpSz+hw+7ugzvcag8LQA1fWSpnMkSPmahM
7qkA7p6bbzBcFzhSwbk/+6sVrwzRNUF9Rt6rTFddzTK2eL4lYEhC4hZyuA+8vwxW
Mb2mOWRcgoo5JWx1FSriUtx/De393n5XUkcKbjyv6Z3H+NZxeqf1pTVrqmx0z/ZY
FrUuDic0SkSC7W5PC1o7kC7ERXWwMsQcNQfcJ4wmzUpmvRQQ4jklzi87ouV42gd4
RkSFNUyGgd1uJ1YkP51azGdpxJ+CydddK1G4lJ3xllOeBVtTFPlEXX6KTGvWEndg
7A/16CgnKD5O0sSxmwT+6HqEuGOLGc5PjLtr1Y+q2e425HgY3z0bdW9RwM5TUguB
3H+YvGP0lcfW6JPU3NTD8qcB3rbqdpBaNytRSR3oFBut8kBjWuVQ+kIKUUjnbwvc
WX2W1+Cf7YQgY6Q25w15ezGJiDEGxmChW5kZ57QzhyLkN/CLJ1EInRjjl6eBYIes
U4tgQiXQx+S/2LX/hbOngBNntOvHxmjtzSOxWdw1e3NnjJFHhF7qzNNMzCUL8acg
CO6u9cJa8rESZVVZ7/n8Ajm9G+6D5+Uh0nZ0IbMFW1EKiDQqGYytYYmGnMV6zeIm
+g9VAX9o+ADGYlz4xTmJQAhGC6dqLJqsH3r6nnWXicILmhoSNj1XncimdssXR1zU
gRQuDlu9v9M/hGYmAZp/wv5RL//b8/AsOcIYJFx+QJ83zqSR1M2xucIqjQSNLztF
adtnQ7HmshgKx7iJp4TPkPWG2GSiL/edoIoFIAVSrVbXaxAq8KgWyaLjkARWve5m
7J03RezZzeSHPnk3g6muTuAo/ueerHKUQhQnvB+iJv7JB8zLpmKhxqLa+ecYr5Xe
wpYfp6ljiq51WzpQay74iu1pJD2TXj43lmxrraGzLfSKLjgg26JnnUxnyuOdyGw3
nP8RbNaOqDAgtf/e8G79IM4w4yYibQT0+TmbbML6uJhranlDBW6PCRK73iAHAhRp
gg+MrV4KVnSmwOTH1/0yV1FGwBvtPQ2ynqWFnrmK3dcDNERmoV4f+5+nbGyXcrI3
JGF4nVwU2F5koKQ3HJXisNZUH5eNRx9YTV5NGrXAs6BR/1oTNrJfJhsayaZS///Q
aQVmbTwXfs0yYlAvhYS1Cx0d8RJSFj1zkBH3HL+W37rLxdqWGTd7SkhWelLNpTmJ
Pz+ftrDnwQhz35liCVvywdlBwvIM8AhWfgWylbeO/CleqvOGe/KpX/6B6IgCts/f
5W6diFeLi52z0quTfeAMyvAw6IdEJTCNy6/b4iIylQqSlGP3o5Bw25KoJJOFXxpi
V2R8q+PN3fEaNOMNC01UviIqVTiZ6iVjb26N0YoDOHZyHjvkQrbKSn1UN+Ja3BfZ
hVFO9ZsuIblTjzFUZCospcK9nbr7u692etuidHMJF+8nUpe2Tn1PbmOkkfUOruR/
mDPNU16zebGkGSBipwSIdWk3CEO25K9dR73wY27zgu5AWQyv4Z2UFRTw1cQCIOWN
zEr/C7rQtM5tXYj2Kc2eQarL7Y/s+CZZz9M3phTDxgCqhgP+Omr2BFBuabB2Tp82
GUXge+C/x4pS0D3/bmB7CDz+lYQ/JEfu6Jwcm3H9dv86yWettHa3Sq7QEgA+DOTf
43njNq/hliYWGEU4B5hJo2fr28s/A2beXTkxlKEcL3Mqm2HF4kRZ4mR57DphMttp
OfZKaYmH9p9KdST1cnOtWPu0ILF2SoVGDEMXhDxelvhBsv3a/rL3T79mqqpZYRCr
//pzQvzJ+X/XWcGOfB08E3nU5Goh1Guneiv7XnNhXSrjLn4snGGyy53prdzBfU+T
0DNJz/NFa1aMEDy+Az7g1lKJTpqYqjD+wxCkNxvxdnXiCWWSO4BT9Ohz8/Juhl7Y
RIvT86UFySx7kLmsUX78CAatD0rqO5CNU26taqo09zNPeMpuri7xYJDLepmC8EIi
CGUImoHs7LS8MfVCQe/SEKHC7DuJgxJuPj5uhi8E6S0IO8UhYEuTlAwZmNW6Ks/Y
Stai67PSGoIxwVNOhUE/hYmo5tG9d6lesNu85UJ/8QzakZlPRbXZeRiR5hBj1YB0
7nJ8kRTz5Vi1drp5LTnYIWXWO5HZ0iijXI54rYCK8W/S3jjf88WAZ6nnMKv1tZNi
x9LVKJ1wAz4Y9rWUz4/4kJ1IeqIiRQ36DqPm1Yia4ROnuCVhKw72FoHRNFFfUKfI
fM0WOYbr4iQ6CIXlN0uHyL5d7ri9cKv28aJEzEy7mz04c9+MzRf5KdkbS5eFpLIL
rIP8SwWYk1EjzwsgZD4wKs9mr81rDebTImIzuAsok3FvJFvj2I7Y8DuNatSFZp2U
YDFsp+mmDhcm2B9u64pNlUDFE4NyrLYHmy8e8/W0fz+nCIhYYLCtIHKqUSb0vn+F
rHLw6V+5IaDlItFIzujdaBtNBy94GRBCXVkbsfQuR42z/pvNXwwSc0F5XCq1gbi9
h6E6+4xuh34kEwlzC19DmEAk4DFWzpT7XFDH/ynwfXEwotZkRMWQLCvT5S8Ym/aY
UQPDBGTI0WCgqBISJOEh5teqv5sTTsO9oB4PX4XU3gTZf/egrO+EKY7jiyCGRU47
YIiwmk0Pkk9x1NtgQBZodj5EkIZmsEZgv35gBJTPQ6Seve8NfwAyh/5cdCnRpdyw
zArwlB1azg+0rg4Alzc3zUeBtLEnFN/nXBaIVEJx+PNkesAjkCITBBefLFz5LnR1
gXtYglP8JI/drhOSB48Oq31/q9MrmJOvWKwYp3yVFarxlsMmiO6qWzpWt8NtuiyJ
bxQOixCxzBkVjFwCeu2JEF5n4QRJu/e6vThCac/8fBH3jZDhZky26H4GdSIvlHBt
yqtbRqhgdes8S6zTmXo4LheASPsDjo9m00XDtD5+N/UDWrYISLy5zS33AsohC15Y
/f1xLX+s39nitO98cvNHMLbGr6pf51Ww8DblXzRaymqv1kcNkFxJevntRWet7KyI
rdtbRzw680sC+mjsjiHaxMr44bv1BmLwzZZoIDnbDtH/K87M900gDrTF3GsjqSkT
GN4/foUMwk7TuASB6EXcMNrrs3SCI8RKWjVKN/j4x9vs2MS81NbXm6Og9Aea7fOS
bqDpeGkdH2lcx2bhZ7OWAQdm2giV2tpWTEiCke1vCvzD9aWrvuDphlzyH7WFp+bZ
4SJSueLmplqdQY4MArmR0lAO8Ynfewxq52G5SIpcg2yA6ucPodPJ9LXb6ZH1BMy5
gnn71wtlRoGTgk/5VDIJkCbKAPAaH2Ao3gZSR6jmHbHcMCX8k7UELTXwq0/Kftnz
rvVmL5VqwIhpH8k62bh/WB2Bn3l5C1xkT4ToJNpJR3eRKvrR6PQUBAvzt1M695fA
oF9RltfrUyHDXow+2x/wO7Ck4GyKYDXQRktkDgAbFe6PWYoeYFToLddHL712N6Gl
kAqmqvqOUbeboVJAGPHC8DWp+rpPXwDXUum2TOd0FPsOa7SbEYsz70tHTf+yg9wa
lojvbUzgh+mGHaSRsZa+ZdgfQmPpoJ56Sn5HkMxwaNamup6ZXLaaSyLsQkBspJXu
EoGmluwD8lLAcduRjgIt1TTMwfUC7Ze/6CL3PzGxoZeP7M4Crc7OXQtYQHaaq4ej
2ItDn9Sg5GL16Kdkb3ZLypdaAlzudfkKOE2ZAf/mHFmQ1CkBqWcjLISpiqH53O/I
s62lop/abiI45r4LtR6aUmPISengpvbQKzwFZ+SSJCIt+8huleF64k48T8HPri5k
11YfJZJM9uJz3FtUwk23LUMVTrntzEOHmQlabCyyhpH33dc6u3rBSGq3ZR5F659T
cyFOUKSr+FTqHREfYUoagJGK9aB38T/iKx0QeiZZda3RmRKfYctHMyxCjeD1Hjlk
yb9+MDKAQgAwEn3y48WN0lYCCEUpegWERfWdlBxsuRB7sItRr8kAKVSw9zUV2+dk
xdRchmjNIn8VCmXBAkLGjG3cDrXt0WPciJAqlxSDqieBb1+ff7Zo0Sbruo7B8giw
HR6RGrcGe9OQW0yeKJhrisriB6pV+DpAgr15kumUhUaP1pvc/Kd+sXRyuDgqWaUd
qkN6/sx8WrljVUFzYzLTbVOqoaBB2VyFxt71cDGDNQVQW6L3bzLSCJXDqxBqZWIe
QBTvAB9Agmn9ojQQkeDpJyIlx/yufJ9CN1oArDPfJ0FJGfgr+vbP02yGD+YKQgRm
R8NTVEctV6b6rZzCLUfl/oMp+FuJY+VOmYOs0AQLuBKmwZRZv8lDLY1hUqT7nMaG
KH5qa7vKiiWWmrQFnt+8mA9JoFnt4luBz9QH+9Mxao5M0j+3AC6yiV0rGdUQNZAI
4y1dqKNSfqJcDp5BYxb8pgYj6RRTga6Ppb2MLYmQbe2W9dc27Z7ZfQQ9J78rvzVB
/5jnIb7+shSKuqvmo+/tH1nT4tWT/bEGmp9WiDqsyc6V0/DNCXLBYFJA/ZMXOOe5
QpUOuL2E8lMGBEupSOxRAFHCAbmagEaShf+XciyCxzRYoVhXcc1iPbzGRvbvurFj
aELIb1fKCJtx8hnkLhkF+XOklE4GNXwpX7VK46L7Bxi8g8YFb8umkD+ENhFL1lIP
CK4Kjw1t2F7cQF4JR05D6NIlWIZlzkWJLUkdu0VANn7+2zhnhtcyRZGJdVWMsxK1
lCmzZjphQIkzvFGvSdMY+NEuE1b89dIVn2lJcbpN67jTEEnHoxJRdmQ6SdgzDZlM
hHpkjRuioyCJUTyLPTZm9iXU14Xg8uxOZrGz3KO3ODwFW1TjhbVfAmq16/fJEzC/
xhWSFmeqec9hPPQRd8xVGtMsUmC84Ui3vBuu69BsKLssGIrNxnLr27vOqUgNsNdt
JINBk7oIOxQkMCzOhsqIkB1I048LnYSFGdbhWRG9b5JGopUJbdrmVDfaJpq/mbxn
f3dC0QPlYDmHHnMxgwGBarXfM4hT4xjThhvyvCkwTR2Iiafmvzr9SXVKFcrRppm6
zNdfQ0BIfvxmtXxs2NSm1kNkAJQEP4xy1Q7Kv9NXk91+0n9F6moQ3rhvJEJwS755
HvqSPctsr7/3bhaXJbD9Ebl5clVrKGMFCt7L6ZM3OANCyg6+QYSPPcTUu0HuoGNM
kIDOjcAd4hbvWpYWwRT88lgILtsed7BGjI55GhSt2Znw4Ch8RyuToaTCEPqyHkHx
cRvEIG78R7+JnXTMF5Caht9PUaJgyG1bBu4REZbsIF7qFvdktR+aqSHbTUJ23xwb
MmSoDBhaJwHoQMxZrtqryPHQz6qINEi0q2DiHQ6fLGzT8YHfpahhyArSLStA3EUa
ZQPsDQhdcHslwGOjoRsKD//lUUK1hhVkGjymTXP+Yz61DHAHm7+3O9QjRwFv6kP8
LQKRrgcY7X0sUesr/dJ9ffXIquTcVD6fN1Lx+RndTQShdl9Ejvoo5NHeMwrMUG99
L3XIEjN0Mg0v5IWu62chzboqQPaPW4mQUfaS0so3eRvrv4wnc0xrbdZQXp0nDGFr
cVeoJbe6m7UTkeH8ubuSasuA57nBmwK5otMOucZPv3S+/WhIUotPV19vXH2vzR5v
EhzaqWoxARIZjC+hND3cIyj7bmW7fdVplMJPAoZPC3c1Tb3AzxuD1lgLvkoFKt8H
/Gii70Axrj0pjDY9e5pEdZSrp7zwbWT90m110HwhF+DnTKrunY37tEYJHXyOxZii
I6n2Mx00p0pwlGb3XmIzUzVLvMxhnZ8Y5KfLuxPm1dN7RLuvBPIKoQWp9NXUxg5u
gGZ8o8GzUedwhQRnVcBbxoHxH5HuJpslfP+XxWE7N4N0112vzvOJTxFf6ayFx14h
Isr9ZXiVzwnzP91QrkgLQCFFKWdNeD2hmqCFEVdgQXU7sC1p1BLuoHZ3xNwelZf8
4qhdOxTG0RxL/+g20CJa3nbuyCRc5T6Iq0qjLLRTbIJyzdKg3sgDM7WIUo/iSS96
D0jmcWxh7D6cIlqoDgnlLZSNbLZO2sLsb9dc5EPGR1k5PFr1GLOFOWOk2sFiJ/CR
DTKTY6s9OleYhr9Mzxf/E59/a4H0DmPVhenKS1OBW1WIeUc4/Do7dMGXrs11wOJs
dd2JQXhPapnDDKz26wSI50Y5R6sewH/WF4f5v7HMD6vxHqAB6wW1m6U9Wkmsg4+H
+LUgA6pXBFrVVsamuM1SYNIVe69amG8tMdJ/EgxWT5ToYHvYwTF3L0nt/4pCcsrB
rlsSwPa973gjzcqIScxSpXgVdEQu6/7a9nyBp2dXyybUzMKeqXYF3rmeUKFJxXhP
m1dZs3POZaELJQ1ZD5Q64eXbdWmYn3hX41GvQyKcD+WAKepsb4wk5xqeGyk2f4Sd
i6Tnx4dluxzgRYIkYRjHoY4MZL9Olv37N2RCiP/wwZVmNaxrllWOhOsAga3fdboN
EhZztD2etZBk4YL9CUAbOFtsF1bcjqF+gd/rQbo3Fibk066rJGddNKD6wJ/sQMtA
JHTV7z6Lq8qb+EWLq8qA8zy8o3j68ghfUowQ09IG3195+b5j4gQX8X7738pxE1Dy
5JCL3O9V/aBmfHAVvNXA6l3hwFt638/+cM5PgH7kPKQSbGGXFFrxgXceO22/iHEg
0jOAI/eOBJfK6BqIMZjhSr16QykzqJLO+HDXQCb0XAHzGDvHFSxqmyh5b7+SiVkw
hpSMmHj/7TqZt/HpVV18+Hh4A0IahPGeP/2mQqt2LwtSQoTT/BSXXfxDEB9uiAaR
EOJo1V6cuDNxEcLpUVtfrc2qeQCsApceQdvnZEjlFed2JEvNDsvAof7A/zDwlf+B
jfuDKGT/dcKvucobPOscHLGps0OV9GrOI5RhFAluWzgMzhtxsRPOJJD91ybnGLlr
ibwT9h2p8olPyrb+Uwa5/4k5O5S7qp9NqL08neojqDh9yIQcJWDvrI/x3fEdsHSR
ruMsq/KDjV/ipmQMg9bhUoe8VqaWNYpGs0nCYBS8HB8uJ9CxEWr0kt6brkQw4gk5
iDISSpsahT4amWTg6wVjSSglI7lEDXCQW2tILfmnku9XJMIQAWOlgln09lpThMmW
Dk3qeK3FP0diP3E8Mdyf77pdg8TPt3c+nUQRtKXLVS2VaQLrUa0mAQE2pTj+1UEE
sA/NyufwpSClkY4q5JN1SVLG4Co1VNIsL4fXIBIEV8NusnaxXjIWfkQAG89vih7n
7bz1GSbanCGrEeETZTXL5zs+CBJ+aBsousaothERa8ui6/32k075pfejiCqHNQFu
yUhhIy6eQWGYGquU+KqFmiFzprNs16F2/ofrXNJCdfTmx/VEE0EKRT+2+L0G3GAC
mI7Uj9iBochmG2/SShIDUuncwIhtKwmXb9/YzZdwixqBr9VkjbIcdoKPIUVorQOj
uRL/OADpNbkmd80MGDMsRIFXx0Vl2j3mt+Prb+tp3olaM5qRI1WlLd5epxAhtsPb
ETmwii9M1+MqEMfl2yV/URK+edjYNlMXm6rCa+IyQ5UW77kDvQl82BOuyydrg2ZY
5Kickv2BYYhR/SshqnqHUw1Vg9V1rSBOZ3GEwVCsJ6EDXUQ1hi2UU3L7iNnT594e
/EKzN78D3LZxnujLkgBGhYvbssaeh+UBE0y/AD65jFBbjwjPXRQbSx8EClcBlTSo
tTMlJQOD1du4t4DLZdTYI+QMs0nUIsS7G0s9lWs8IfBe/md3HRtfBeDc/Dq/bZmb
DUoLBr4fv3O8Uu+GwQjy4nM1yMNfgywuTZmShV/RJOzE8PWUs1GGdMdC9JpcdiQX
p6IdHrTLagdPAVC7fptUDBRBjlTHo5lFs0HiTSbwCznoSDNIfaOsgxJPOV2NObmo
yaPDVz3JLu2d4NRO9XYGPZAvVJSmrHE+MZUp5cglrA31hr1DaNF5/wg36HM/CfWq
FLlsgHhC8BvnnQbk8T4PNYiOQkso+uHK9OChI4WAbPH1fjzsTwejpV4hM/nEarWO
Y6lSqvtGCk5QKNbdpgR4Nd3VsgKeipS2qsfuKwrBmC6gVlqtg7WNY/f9PmD6hC9r
MpESWcxgkImwJ9jcV6XQH03brCqz+hUUgXLtG/H3WTW2XQBaWBgKU43s5kJja75I
VbGCLpsrv/nLki3RJ6vkmws/yUonEeey0wEuF+3SS2mC11BOO6TNyBMpg5joK5wu
SstKKgBluy4lp3JtlFfDuRNeOzB59TVF1Dh1R1GWHzH5OECP8/FHMuFYOHjH7l/h
d1rR6ZglcWadmfwrziSOnApnnGmuydDfA1CEmYeoiF7Zozi997LsgP3q2q+9OXqJ
Hl36ZEY+An4BGCBW72gSRU8IbfoJfLrJmbFNuAbFqnEpYXwsNaZEuEH+pyvhFMIa
vcp+ITSZKOaDLbimwuHFw32YnJpYuFdSNKXVdx0glzl5UIwiSD4b6M63Syz1dXQC
8dTjk22S+PSa10529yuWhrFaaCiJ8FAVfXA9PXXRhgzIQUE3ZXUChNGYUTFFAiGp
3O5ghIvMC4OznUiDx2zIihWrA21vQfsWTtjVAuYDmLrI52ENOsxQZ4KWSMGHexcK
06jf+jlOqSyD6r93mQhJ+0wGYmdzdBnwDOblmgJVrMIcSizYEsyNhssp5zKSYs32
W7S7rMG+DjZbfn4PBG+iwaNJj2YxUjZ6iNo73BSr84/eabYzNCH83SGQVmpdnvst
sMbGwjGSPMG9bhll7F3IYuL9dMU8nsHdbg36C97uaqwd0VSZ+8q2YbRHiZH/h2/+
mIMRoE1sS7DRkK/wDvEObEaYuhToAj32hDK7iVySI8Yvfivc5L23MkaaicYQZP8M
WZ7xfCpEPDyD1yaVj1ylpcp3mB+WS7w8OLT649icYmTWoYnisGvR9fa7Gk7QNewJ
XDZH9OSnrnWZNJBbJyTsBAqACzLsdfZyi1uFQJJP3TVb3VzIsdHW7XlCHug5xsRx
gcKm/IzKtVlUDkA8tYkH0vY6p3TEOJgTX+jnprPwlnlW6NZit55Fqd3zPFH5MsNU
yrJ9spkpLVfB0xHIqFhc7mnkvIqPkerrtar1kiY6rCyuKJDjTLn7ISIJ4E5hL+eY
0XRLxSPMkiF+GTD8bpT4hmNW401PRqFsuuWcT1JHWiynFOG/9G9DjtftTdLLRE0n
nWHy7P6EX6SjJEcfIcWaefV+Vux1oYhsPaYMUEAvRRgLeAJh5zL3mVIho8J0BXjX
rMGuxL665lz28MY8fYlz554oqV9V8kPZxAZO/xklWXNT38H1R6W/NwC0CXpJxHVv
HeV0P+TLKi9mcx2mrRnGy5peFiHEsfCp5UBdl6Fe09HQjqvgzHtc1sJqON1loj/y
yW/B/DMw7+LQl8AIeB0XTqXWPfWqbyJIreCjxjU45eWb4wTpaIdRw6KaHTJxJ6bO
OVz8CJJ6bJJsrV2Uqv4tTEPTzO+W/jv1Ufg8sQOET0fM3UxFP8wbFet3KZN74Qz+
LgxjUHHhgLiZrpQwjl5VQajmuQUdYPOjZXDE4i86PX+Rf8fHYk7NDxuVpxNSxsca
m4vV7M82MQTAUacaFglnzr00p79bVulJWenq3NaptMdAfpjxkLla5s+/U9MZSeVk
ru88ASfDZv3DuetlIpcQrH821w4JV9ll4Izdjq6EW+9f/+4waMzU7u+hdglzB0dO
om99NXsgTEs5WQ0cM+fVF7vBspJhxIAiYLieoLDOWA/RDZ+xJL2eSUJi0uW5h9Oy
kjgLeOvu3fWo+j9lzLtkNlCrbqvyZW6vQ0FY9I5sIX/MOoDIQNT0gxiez3glzVJZ
FiNkLqXwqxZqQmLBhBae3vll4r6Y4vKDG4EOvxjixuNCjRfFDrWpbZumuO8jsZNw
Ttn7ZvF+LA8UwFgIzrmuVfTMEzQgmmbsI0TzCta7rJP/HKsV/6lFMxDtOHqhTAW4
w5Sz5BptWDXP1+oVdTT02crVhXPO03yrM9igapucO6HeUA++DQDDSfQbPinR5+D/
gRPxN4kAqUCxKbBVYDYe4ovEaUtni2Gwbh57vMYEeTjWC2N+OhuFyNVLxPlx5RuE
2FPWGtfjjEUCfzJjRz4PcdTW0tP8xhelxKuvIlEwjFIRg0+aSutktwzc1e5JpXgP
sBrIpt4IJWaijvWWK12X1pBLrLuYQl5OgLpL1LoyoNWie312S6sxZ/5qSrZRgFgq
6NC+NKEo0anIwj7208BPzKLanLlQHa5gy5FMbWw9WO1bsW6h27T3oEkfdIrsRDts
qfYjpEApN7CUsbFVufuCC8/vX7/1Jet/VT8jvYrsM7mPuXOBbKVXhqulXqGAN+Ll
bB90aNVb9WAeya66C9UCG0W7CgQkKOfnHrzHMvjlljy03eyxV2DVYFkjTmDEpuyA
kcmIKesw845s0TFoUHiH5o7ZZBx8TyR31foJaZEpBLevzOKWt1H593sETZLfGSfU
t7lXB9QLzxjBHxrS+lBKdAWR+rqdAncenJwkaKCl3TOA14+VMLiQ4CrtnYHPzr53
s5mOq4VrrZaqbG4GFGA1/yEWBh7hNuljalBMtAZkaAR/7paBQEkwHm5/l6hbHdqN
ZgBh1gMPyGXcBpfCbkJSujY9x+TgRT+Qipun0fcil/rmcMb/tvZBH+8YRpYrrm9v
/uoYM3tUO7VnA0v7+fyqCnGOtmvryAnKQTQUsNX0IFQk/O53nngd1n6RM4EmWWZC
yrCrVr8dKn731L+fDp4wwneNegeFvRDq8QteVCgsBipV5h2+isAeAkOLhiWhDK5f
PM0HezhXCygxG0Hpc7Y8axiAJZJbt50/Ewo9+5cAwL3sTVii2vU/d1vK7raF+Jhr
ENk03+fy+fDnmmXVBsXDy24jAMB12cgZ63IzjzXuA7cP/WoB7BMO83RZgXsaTRDC
ojkPTKhRBrdcx0P2lhDJmM1U5ppmhYpN7pBA4c4bIuK2X+PpeBGdyyD4ryiGvhjg
tgLolQeMeIA34qYBLOADtMlJhD4l/z7USBcyXACqNbkcISAtrjDYWCNPkzyaPqNK
Y/VmOCXU7WL0ePrsfCyPveNc/VyMOMQZaE78uhvX7iuIwKnabL6Vbd5q5O5PGo+E
vg61dmLxyvGn53OK3hmeaKd7WaMTGUaWbGDmXsTt82vheeItnq16QdigmGAzXAtD
Ffb4hxzIhem5sdgb0IG5yk/uzRT23HLPanN8hSRPCDM9HkiqR+rme1K+7q15hYIW
GrbatRkBwje1w8AMia+okuHGSZLhEvY3CHlsmh11zllZEWzkZhUTwrHfnTd1NTch
SsKtH8HBUwe9Pnd0sIXfrZKldzvTRPfX9bc7QPCxEgvaARsvxOkAlvuS86gLaUFQ
7IInypPzN01r1vo8E/xOhtO20ezdZqrWf9B5RlS8OQsqIrKSlX6XfWgINtnsJ5+n
iaQ+zYH6phuy1Y1piICp7eP4wrB4OEnP9Z6AGDcJNY5IC2bBYBswP1vEhEpQZWlI
kqlwxCeA+steOHyMOowec5MDUzRpBpxgSXotH2yEHNQshBgALnEIyU/wI+MWu1ZJ
LmoexYwJJTwiDpZ6O2fM8lLFmrMaYrxdpKaU5DtWXjuR235pKLz1ICkev6C8Nb4l
TVT6XuHm7DyU8PtbiJW1uxswqbawSw00WmptEc8rkG52IWjw5mmdKlZu7nroGaLr
D9e9fsnrTWd6iNibv31vhDLvEKeBHxvANks5LktlmzzdrXvhvQx5cg1mjCI7LV07
wnmk4hn7qvQ17u3I0ly8qRBv7FYOSspZdszAyuSJNdzKSOvj1Ml+JeOhiOOECv/c
AgoL8j4MdnfeuNIdNPhpfMAv58sM6CZZ+qSTA+/NhFaq1Mi1JsO7K9W8tqrvarNq
qFsUngDrcHyGKuK1+juKHq86wU+FAvUWma+yxCI2XSvE54DNsg7nIL0O2Cvz29hQ
5LPNzl/oP0C9hryhq2yvon/0Uft5bWLMbyLS4sniDAJBalA8IsutzdxdIOJ2rAiz
f0pe6gOtcUyCUoPt5NtFL5Qop3/20vJOrU3puLGNInNyZNHbMDkMTxrNF74pf2t5
MeYjgDXX4mYTvKX4Joj281wHf5ho8b9m5eJoldgSOX6XOIEXKnmfYsn9jx30rx/k
DlA66CBNaAOnhKah2WftIHmez5+09GSiL2k/0fLrWlmMJIeaciYer+CHccBp5tos
RNHSy+G50aokKdW2RZBNhRxUldxRswagD/TnG6uyqBRsZ6ilwUrnQ9F9is5KeTxf
6cBO5jBCYjYOlSFaQtwRWU+kP9Y7ujvCimEvVwUO52N0INIrWNh16udk12K/6SDk
LvV1l881rQBVhoGf5kNSfyrK//E/q/hZBy6pn9AEGRKNIZdNbmW7iAejKeUfQNVK
Y1q9cO8X5RWnu+G1wB1Mv9h2Q2DnDPQ4wNli33o5MIgjS11n57HeLSTulp8LL8nO
1Sksv/DuhEyhzjmvbW/e5bdLReDSnuA8c03U6j4mzEklC8Uo7w9CzHxiWBndV4IV
BW6ALrKgdLlpKSIRi8p8coHE/Q0AYA1NIogqSDTJfESdyPNZBzE6qKRS9yPPvkLd
HnfXAn1jYSn+a9ZfcKbymjpUMhCIYlNHNXHDQrKfggca2cY35d5Ds8HOcXm6HlD7
JcPb+9LIOj2WdGmddjVhWTz3RC4fw95/FlwozFiigYdMk+wpht1og0OgRl2U1S5r
1E+WOR/oNDhRtwmtLGrmzxX06oS3itzJST9SElFN5iHnk3sUtyCgUKHQAXuC3Vpx
O3kvcy1NCloYYmLLRIG4wskSJogszp9X4q/xHChAU1pR47uGRF4uz29mU2d+Srmk
MqLbTlsWIhYwY3LAlbDR4OE8VZb/QdMNyRLjrLUP6uJPNcjz0pmLpvrs0tOm3t42
ja/LebDtR+nNNA3ohZ6tg/0E7u+3vw1A6uUWxR3KvPeNOVGgao+6wOSfdyOz3w4X
p83ZCwWtdXSfLNgXbyG+DuI+eIMfJFLM8Hmglrs8wxAWzxQEWvGOixBv8dPllP7u
//8l7QMnEOvlnFy5EgH8bcCETpVpZ5Ak+Cbd+02EDJz3iEh25voFsNmuaIiyix4g
f8h2wX1lVk+ycTwFpcMQJWXCKtJhY2VngUAhU6C8eBN3ev9xTojso6sbHVLIWQOf
q4k51EI6Zimay+aO9VEci130H9IJ+vpzZWLUmluSOTIe+Gv8L5qiMnPDDbq6m7qc
4qaD1AJFRa9e/5D65vRJpNGkmwWMJXDjIadMJsWVhaZmlrCPYRQmUpgiJ+PvEDYW
ueHhby9Z/cxWHvNuB+XN30aS+bsRikyL8Kf3XGNOstq+GVnoPsiV+PCb9Bk1L+4N
VFjq0eT/uczwFcdNTvgzJsfnA7c8NiVpv/HEA8EuJXpGLd6Cag28APVmYS8H9aCx
mdIdapgMtzIGFt5ZiMvwkXNDG/79GX9VXdPGSTy9oEBkralrPi71o4OXr66RqQf4
P77gwEG2g0fwU4QBQte72jlEvg8HjKf4n7AGIcgEdOPjQhwBDLeAS070Ezm/POit
Iy7Z087n0nOCIIv+QauNoMIgAj8YK3YymB8ORjU0/4t2VcVKNLUvFM4LMDvLzBuo
NdpyfGP6NODrv2XnzLnK8e5wZPrjyCesZ9l0M8PEShuiit6HkUUoVbdr41nDaFFr
IMqeVwD091KfkuDrtLXa+XMsvPf80qerkll2kVjvzHaUPhjEiSv4rYMGW6rKMgeE
o8vKp6P+II3g2mxtiScM0UB1l6NTMExB3giFSj/CXU/qGhv8H4ZABIMt1RX5sENn
9QpWwVmGXqWKRrM1e/JLjf3JKTtNcJnuZdQqRkw1k66ey/JGmtWc4Jfic9sCxxwJ
zWw6HeRW1kysBMb3eHOq2JoCEhcNXxLoIXu2IFJhhGrM1wk2FEJFZUTlytZUjeXX
RuCJXjLzMcepUF44krmkq1EaPHRzKsgnkBRXf9x/+cKhghcnt285XjJ2nEAt368m
cP8pIIMxo2xBLLvnU7xax2OfX7uRh9LvpwvWdUDxZK06nSWxP5TW+tjpi4QOYFEC
gb7/gfF0WLC5GtanIzp/GPwGZLybpwUiNLxUkUVDNctfywJp1kqtcMW9myCfazuB
ghpcH+ZnktBdw55B5CRpe5hI2f3ePefwAhvBqRu9Ron6JYVC347osOAK9FxQoZHD
RQ8Ezcojm2B2O2vIhIhSp5fPKi4CnU0CtzofWEjMpBZJ2+Rujs5B/otgYF4ZJwFS
3kDLtC1YZk0ajwXU2Fo7rQlczgNE+xEQ/Qh7cHBTVqrtCCKJvMuVIy0zS0O7Sbma
0BtwA/KGD+wMzkhNdLjZUiyiajHYOGHGVhC+zdUmTH/nIEZCq7Bmxaxn3/U4zz74
gbpo+fLM9UvLq6/lLrdLFbzvI+MmFiikUYSJD7Icvu8pQYGdGWC/CackwY+z/TM9
1lesplwlJPmqqJl1xAi981YF87gc2lN7qQBx7qEcVg/0wbmPo2jp0tHXbkZyAs6z
ajiokLfifaA+ps4livfN6q+Eb+4p7J4LQ6pcz6fi9RjGCyMizMQmJ7/Odt66csUf
TyiFOm0oG/XRpWRUD0xMyBywBk8Wea6bgYH2b5wNZf6HIhfZkE2xqXvLiFlW5up2
etRGtOTyHNezMaN5/yRp79BvljIEXb5mwQ610nY8H6vN/4uAhjYHMqwfM/jj0DoR
FhuZ9kz19j2Ob54MpYPaHjf6wiwv5XDuWPsDOZsoxgNtV8yXFCszSgbcV4hglTg2
dZYXA+r8YZ0ZIOu5RTJWzXAeLQQIut2IOnslvLIFy78dCufhRlGezS9YfQWgTFje
qhlDGILH42rNOhB9oO816K0ECBgj1OiFL/UbobPW+MpU2i4R30e6COMwTLKHCwDK
pVzG+xYPSNVXO+cPh/RN/3dLB0w9zZ4syFsxIe8L9ar2SmFmbaM3RrHQ6/nig+b7
Gh0bPyfOwj7epEMXAwfM5GLPS2ernRXPkmKr+2afrSl51mmQuReyi4Exod12mm6E
kcW/h98nbAuiRimrxW5oSPzVZL5m1+Ogp1QAiDwBwUwWA/fK07D7vH1HsbJ6hPua
kSNMz96iDdVz+UJi3FTD7F+7l8/Ne8a480tIRQJRd5T6JC7eBrMKVNFgADYnLdZ9
VnUFxTts14y0MZnKiOih/Zr4CPG/j6bJBLkm3nFgsfWm73+xRdNMbwIoz2OO/qS1
YlSlKSRXgbGlzYhWFtk59Voyt9xeUPvh/MHesQ7Ke5Jtv05Oynt+LCaGGHPch8Bj
VgSzTWdubQjFgutHIGxqIjnNXwt2V/DI7lOe/eiHdwsqvvtrydg3hmOtnPFbjJVw
n18BekWz3W79sFSDp/4Y8iPVwtpfWbi75a5wtOV5lOwK61LUilqY8DJF9tB0uh85
oIoypjQ6xos6NDS3R/2OYBp/3oyO6gdEXuYbXNzQG9Qb4EdHTwRgze1lUAzEdUuo
7RRx7BETz94CuW/z2rfRAh5m0ERMzzUjTkMZN13yOdbkdgWQnkZ2vA3maciNbntf
E9YbaIgjkzRqJ1HqNJqVTWnYtUo0nQYf34dLKyTlQIVed0VexZFtsunIYGIBrEc6
cO/D6JyuoRBAFGSUOFdamya8jGzovSusCqzTCk/Or/os+AXPqLeZA1wJ9KUAM3nI
5zjAgUc9qUy9/GIq5ekT1Agh488DYW1NP9uXf++bQooccn5nTbjzQGPodkbEUoBi
PKb8n2drfoaKmNEuu8sCdCk7+1MlHTZbVvZfEQEIXdz119K0XHp6EKydmLSAWya0
aAg9aILkdG4UZLiNmx2FzGP4QPIHU8XHt7U0gidaEuOcDyPFU7hgrN2qTqXhy3i0
zJvdqTqGeIyIj9ruIogKHXz+QojPd9iQ8Sdm2vH7P4c5OKmYhYqKtFKO6YJ5Gs51
YOJax2SID6d8y4E8dVx1ru2QwkaEmtH6yWwK6xxp9Q0UTzkoNrl+hr1R7hgvYQj7
DmZ5mpwZhE8P/PGvTMDZz1l2CpfUS6fGtaZRgDfv3laiaO/55pBxAAIxtMIjKl54
2nHv4im5AqVkbPhNV5u63HJdMbXeak6AxeYj9k41/Jyk9lSXLv0KjNrtB4Y4pX11
w60XDlWMQOVcqvIsFYccidn3ipQOHSrr7ZaFVBr/kItShvadf4a3Se34WqoUTywt
sRAM8R/TjESwLM2NJ6b93yPR64ogAK0P0ldFrHhmCT+KskDH2gOlJEKXEgIYDiEa
ziEJ6rtJ/vyUoUMLoak3dgYiwc7dn8yRn26GWWuOZjPaRJchY4cY+WQhhJQLtmoC
uaTRU8oTAeNz8jv2sE5hj7UUmRuY+ph7quuZ5v8h6Pe+nvODttmLVOUsSJqmeloL
ONPGz/J94VzbuWSUCdIaRhqRTTYyXirOQz5wb1R5r6wtW8ID7An7XqegYjK9iILt
iXyuKN8AX6S/uzoPho9hZGAwaUsYSmvVBg3QCDcsj+XGcURfhZmwEAj0+7WatKeR
AneAbLB7o0SNmwQmI4VV6K9gzbmBCMnv9pw3daa/7AfgXSm8InmsZTgdYbuhzdL7
dJvoQPuPu7C91XpZ+Z1Avvv9oWrGUVfTp5sdF6BEdl791guU2c15UJpKBlVYduNY
5ULSFbnHBJ5vN+HuNNYORsa+w8v5ghVQxNNk/dAiVvWIBN+Uz3p9TTB46tn34U82
2tU+0vMGVQhu0Hs2Tz82NLodlz72f/H9fWXpo0nT5ZBsoOiC0DgZ/9JA066AA/uG
shdF4bf0C6rvXb9MFNzPvoJK9/gu/wG1TvN/wkB5A9O9KKOgRjnC9EwUqsXIYfbK
x8l500x5ooMMID6Euu042e9kNTCaUy8dlTZg+ZX3YFUd69H6TIOHXLvz+rH0sMEN
iEh3e1oAEWcf/HXYdulqB5NRfdk2/QR8slcF1qgaYkHEUmOs5htdNrtRfNInHiK5
Haj8NDHhldyUjRyxcGiCbMZMGoIW+5Mu5ptm11uM7zjubeBPbNgT/ipvYg5eDPkg
38i/AXqtivCdblRd47fQgjJ8koKV2AIPFYD0W/YL0q73X4k7+ax3e7sZjGHn4/k2
2jbJ8MAKLKB7ypIZ++HR5G2/NiBJnDzPEIZJYAyFJEjYqR+wojMKLxFPtFcqc4hf
0NzT4XOTFF4X8yDKDHlZ9vH4hBYdZmiHDWJErxuHE5uWwTi6YXnTqgmmnwlBUMrl
WRGnyTpE+bxnXmClCjHPHQHsZskfDoYIy0Ii7S+h2Np9McHRtlD9ANxFZjhWmTNN
zjYWfn5deiqatGo+zJpt+TN5sY2TmUDA5obDOPI8yFDRnPbYMf0kACaiG8cKrctG
y3O2KL+TL35QpjN3d2hrI1dHmis/M6xoSyML+0I7E/cMaSTKoGtspktNC6cajd9/
x/vCxD+6W5cavF5/f+Nj/BVqrQDvpkd6qwBDV+NkAyMS5EkUw3leZ6SqdhzZLVtO
PTpR6bfefuOmUQtpV4fvyapMVJYq3Ht2mcYiqsDETpTDEkmhvzTlPKVQP0Pvj1h7
G+EAS2rrnVuyr0onxH9qsbobOJ72OI8QjyjsyReD0+BQXuuRaqVmKz3W4QT3I16k
XuuWB3w0/CB5H30IHwCKb1vYxkjohwbPXjf49lFhhg3pGon3jRkeo049Nb2jFZ2W
XmUADVaoUR75Qmt/iY65eNlQNsAWeRlfT8yuwe40vmBYDzTt4p3ePc9H/J5xrzyR
d+ajtnDt8Z1MAxOVfAltxNLGI0rxKWxm3ZAztu4OMyUluW/O2YybkqmmkwiqHSsF
PonuASz/yBZv+1ejKB09zj9eMmuNg5SGquxVhu3tz/k7EjJv3xiBnrzC89z+FOTN
MgxjehZ167dObzKHU9Vd4CnCLtrF2cLKPjyMzQySdWGfc7cEXZoVX2IRtnued9LX
FdBKni4Qdy1MnvPviNR1pGNTs36HpFuamCeqaA/ur+d+kRO7TkcuHsCeRp7KrNGi
CNII+38dKMylhWGqYv1ZHFOUo8R2bxOKuVG+IFn8+9IAY1zML5Ct9FzOR1noHg2k
ZbtVMLgooXbT3EoFryoGQ0rBY3vdIoc/zD9kDyP/q5gEeP2WXs+w5+gSJY6dwjE0
x6VzPW5StP2Bs7Ps16sbnEdkWPJpXhX2pate+VQGkSXH7n+TE2k/HZJ8SZW4ng+2
fzhio2GmhF5jrPo8oqr88/ZbAu2nMrfIbCVVmge4rPf0kyZYO/o/sZ25q/3Tmdxa
+yVB53Mq7TaaYjW5m5XXWM0joDOxgeJ5LyaSvFkZUAJOEL5dN+eL/Wmj28UyGaUO
u/1CC8pjU+OjsnGaeUQbaPPvPxV9f5gQT4kMtbHjspcmemeUdsr4AaeyqhXoLndS
eoDpWFnmrIYefMPrKiy6x/Dc6xVu2iZ/vQxwK+6GD+ZzE/SIXXgEc7GXNHVHFsQY
MGAlAqSMu92oqo2uAoULi7Q4Z+bSS8vMSSCWAF71D4TzP4Sge/qbv+8FxN/2aFis
wYhBNYFRRoTfxrWawGnO45Sj7hI/LrLd0fyDQ7QQ/bR69mGZU/222t9V6hQl1vwH
x/uql1zqlKr1P+6/kRp4Pzv+WcJ0pZbZ5COieHLqA2KuM8qPq/RZLFnVuk+4rFlN
8XOygZiuETpV59zrA3gD53K6KEa5sfFgboDCpKyUgIjsc/FmzWcXIxn8+tp7vSok
41iWjY+T1qJClaiS3uRGcZjnwsBKMf2auF9zQsBNfsK/cZ1lCJ1Als4SLmRU21m5
A5jyAlegKaYOHILWoo3zzyIzqNcCLlss5Jx3cIlBoi8U3DdJyWeXx2JTQIHC7UZH
OEE6Xvea+eg6cIVhYT8uIVNtKDaJu4qMq/2I9wLUArwNYFjsBRWXApIhafryhRYF
KVTvIz2Qk+MaZMfNvNPXCZ8PvFM/rO5tAgVss9THp0Gv5ECKrfJ23jeVF9RKACew
Eh8M2Kxs44xHjyl6GSMIuCDuhRM9n0apbIjyyjM4496fpwP78vbHIIvKUDQW1LSl
Szj3gVSLq2xH+wM7E8oCPThX3ZJufT18033UqsYFGGhHZWJjBRsnS34Io2RSWe1C
UP9iTvAoNkKVRR9fwNlM5dfStzO8KPES2HxBvJ7Vk5OyPiKiGwhpfy1ax3QOd7Fc
DqLShYNRosKEx8oWpNj92o8gebyjlC7UYfypsDBHoef/GdF1m7Z1LF0ePDed8wIJ
7WSUIYCl6/8Abkt0e4q8C1fo5Av7VXL5I1SiGs/TX2JanlW7gPr2o1QVjaZGP9+5
lc/Qh81WEPm0hlH3ai19zV1YS9fkDuUh0ZLiMriFclqqy9N/CkJOtPWZa4lpnXVF
NrXyuAje/KNfCIZcjkw5kRnwSi3VaEH/vJLs4WfUHvKYJVx6fry9e776wQPiPokA
qEJttG2EwJR0JnSCSiAWG5W5pxIG2kOVGjEr2lnewl3Uu6K78tC29JvHJYTEONex
dF5tfmQ8IkWK1gGCwqm0cx05gEF78CYd5RRquFTtnZkpvp+RzsRASAUTnRxUn7bb
WFh7Dna6xtbAuVWQELtpfNr0r7Lo36KKJ6U5wTd5TekVR0gIrO7WHdH4eEDEZwPA
H0y+oDJIR6vnaX3XXDH6eF5fzzlubUIwF9ahBi+Oc5ST9IuCI/9DpoT09Ce/P5im
YjZY6ms5g2IUxND7wRTedPSVa7HXM5hyC5CY+u/m2dUB7F/4N5Mx+i/SqerHRVII
weHHBraZcgCsP4th7wBTgyN/n8eqaorjs/F3Z5+yKAEVhbGyRJaH3QuIZgYcbSpx
x7yUnRSxMwrbRw5y7zi4+GN2+cmB8/jtXVqpXT8UcwEP98SXgt0hEXT3lL3HOjoj
mN4Dvlgh0XI+lZWq9vrcb5b0V7R0Jin0aT8unjPT11Pcf0w5Bn6DWWWE7MRCA4cW
In4/kxCNtN6RlpFgIVTD+oAlB39q2mFOpzQQK7iTpl9AseXwj0Z+fcV9FASpRO3r
WnCwIEw3NMHiIbF/muqPcM/H4C855UFPODG2mwKffxanWsInzpfghNJweadUjVFt
DB2smPDMyDsqXCG/iKFw9igOUg6jMOXW0LJ3pUS7OH9D13gd6Ff4YjJDf+hurJbE
oypCU2E3i7YYxb0pLo7cue5MRfV2XH3vJZVI5ehTkyUK6FFXTzROKn3I11/VIJZJ
Ayfp50/6qqQ8CPMecLBhjZfun6Q7Wk//2TMZ2Ydh4p3hN7ZxD7BCyYdDRIWB0cxn
go7v48buosHu37SSzDWD6VGxWoPZ8mvzZ9BusmIL5tHVDsfNtu6a+Av9i6IW9Xa1
HCT230SuXKq7zIhPANg+W2mmTtZQovH1Pa4/1hevqzs3/2o+t42HHmCWNDXfdFfr
YgVCcFGAhVbxxcc29ZhwxTXgDS5ZPz22dgo0ZZTqKR1mfdfTVMc997abg+ob+CVR
zM6YmSekiPJYOQC6mBGenLqMSzy237zDnwh/nanBW62zYa54vG5idzy1czxtkE1K
kUtBMCboYGhCsyHJkAp7ZZhK9qXIvS5P55VpGERdY3QUA+LhK3uwssB7mBO2G4RF
9KubYq03DwCwJG62aDcDiDqGjJ2EPkR8L/b9Wu6w0FuNre7joCeQ3CuIngNN2yMK
+cXCS52lfqRc43CQGO6YQwkRiW5SY93cL/rYhHLMui05RIw+2fkTAyT52D77kIXm
QK3w4K8mXUMwQnTJ/HCsr4oHtTgh22riAbX2fBAHImsQyI3fXG1oiB3S0RqYzFdM
IysRk3E/gt1ARKoWV274fvXeAfkHKAPwLQsEtakSI3hPM+B0m+LmHfCZSAuWEuh8
GQE2hRRvgWfgV5e51o81d+3OWHBnOixZQcC22L9ohGjQfrEzMTC+r8ssMjpYBW30
NOimvJ4gkqzU/SOeTMh9gXJLixY7l5b365eTQzdfFv2Ozuk64wFeVwVaCvu+0DQQ
oX1+e2Cxh6RvyNsRLiodLkTB8o2lEbaorhdka4M72+nQQyqgreuF51ct3miXi/NW
nNSeHtX1LyCLwiLKqwkNyhL3sOhpwMyg5A8nAc0kR83Z4cGCNQNgpQ5a7Nq+yOYN
t5tGSscrE64aFTFHZm0i+Gl4mu+zHqtOeKVYzUSQhzO2Gnd/TLn79Xp2NLpJUuGV
5cgUkWC3lA09G+g0CyPg8iWdF+nzQpeqr5cvI3cPQVjvHG7ihjh0hCbGKIEbRW9T
15emNdQqoAzCO5IR/sHnJOllKjMFvMVGc4PcLQKwgCBL0zvNs6/4tcy+99m99WlJ
7fBnsJtTXv+Um6MJQE6hb5k4PS07oCE1nWOkxVCEuQzsbITD9ssc+lWMBZyMXzDS
Cu/iB+pzAgOwOWruLO0w2JOMP6FWIXh1CUWnt2MYgCPxYmunGk00zU2VfACAV82U
jVe8bGHlD5OIvkXdALJsyFSkaM0gkpfCOORM4nkq8WMxeaakWqp0RakUqJRC1V5W
hYiUC6jLf0Zk9KLvylrjMn8wBZEtlppMwIP1Z8eM41he90Czs/xU0p4Cc/e420sl
YDBonnT0MpXWyUP1RbSxYEkh0Awz/oFbhNw8twXkALM7vVtEbBarPKGtGr8Mo89S
wwe2JvPxwXvbWHnfIPhcF9S2OqlufQMRRt4zDu7hhChlgloI5snfTy2QEAyNYjMu
lJLtGU99HtYNqaojmYT9Wl+roGZgWArqpLM4x6y3nv+shKI8ijnTKZinmOKa+nX4
vL99JL9YWNIWkn/76a/FAOyhGeX4DGF93BUsrOcVBPnHTDaOdwEOSVKtItE1qJaE
NFcf/I0Lq4zeMSwH/2+oLlrfoe+m1VVLeIIzFc/STtjdMV7QEoY/gD6ZAW+Tr3Uk
uRJXzoPim/sbfKOAU1cXlsg/eGqx5k0yRjShT8R5rqnUPuh0i+bs5JsjUoZr/cs3
2p1F48AEo7leXcPKa35A/ObdQVsX9D7EnHARvJrOdC9URW2WsgTZpIZPVooMqWTZ
hk0vYeKZi/zwV9w/gOO0lWyyOTiCT1DhQOa/1Ll0RjAzUhT2CdTeytpdnRRqE1Gl
UKiWt9IbPcVxjX0UA5W5dJemQcphbw/5x1r+Orxdl1XV9M15V/C3MNsJ1c7bBfC5
NwJEGUxpvP/6bryeJ+JKjjA3qdd/s9QOfnsSoQtWuqchSNBrzOvET3XUUODFtzRw
5vZnIlgV3/l1cwEpnjwh+vgUQ+E1E9dRpWs/HUTJLMqvsY98Ts/OJsk+sQYs3imA
RzkKs5IhRwPJ21vRLMpQ3CPzFKLQTn+Tmnws8+qZGUjeUW+O1/vWVA1MdWXyap7E
WyVV/otf+8MyrEjOC3V+1sSV9DO8svjxs+VQSLW4xLI8jMH2Aef03cAKTw1VOwAS
77FufR3J6+I/MWsPHf/EVZITj0AJ11JQ1VUFwKEs8/kMvzkNQeirFNGNWGCIHBiW
IgRNafjabybxaNLy4Uq+n/Ze+DIQ+lkvEzaJUfy4X6QkxAm+DdlwlaQIL5m/3Zp4
Nv2RbX+yuFt8hfsKoZ0kZ+HyuVWJnLE97/jlFOT0iXVZtGo0P7apKMhMgdZz15VO
B5BHelqyOAq842F5SNyo+iuUZjWGqFwAZOnaOZgnKJvzpNGgNCiMxpmvZ2Lbyfx6
z8g2+io9tUgYAj6ev45FnKAoVMmdQAiz7C4ecn0wjJz1gQqVqoTQ5haYDHBORk1l
CzIoQre/qAHWKvC/uQPhgZSLCcf9o6MIKw1KlvD5lbKYisDOMeoz03Ad4u+QOxgJ
z58vDaLsy5AcRL+b3Xth9m3bKckw4raQ1o6GsK4RG1N/uuduHElSh1z2hOk/QUJp
xYxAT8vNPMx81vg7TCdggmFONm/w5OyBKTQZi3wZk4S3srN/Y5q8WCAY0pxtIBd7
v/nZmljHx9wwIEkRBTNwC4Yye8kNo0R1gtukJPqIIxj7DntryfcVTiAO1GbsBJyF
rKZTmaRW58E2/cnpYKtfAGh1ehAenOoz3FHdi7+g/FDTfT0h4ulWtpan5LY4PJdB
AXA/LzqvUVBqoULIl9PkzUdu2Uc4D0GsrMxEMDvvwthirrT18gB4qFHRvGKhU4e+
JDTGJhdMqdybw8qV0XKcEhwIYrmGOOPZznyh5MAJshpSu9L5QbcDaXrYPxLDTtQ5
5MT5DTHb2odJn3AFroKYJv+ndB57r/tW3EoI21M20mSj8ADnHa2J+G7WSBMlmCo1
10niuQO4ssNue9Est2VOhPr/grAo7d2WorDlht0mdWr2aiebgcfVTele1JtbhyBa
yZ899C1OT4zTVHhS3UjidqKprSWJFLGFB9WdfxGpdr2KGaCnIGAyGCC1el0fvl5V
KJOLTDunbwaT94rEgs5ltT40n9lpaWfeON/T5i2Ltkm6YX8HVNfZhXHOfCfexjqL
VT17l11Ubdrwa2gGd4N2fmsI4zDZC3G8dQsJyJ0a4fvvnIv8oFpNnS3GkJ4nTRZD
mkdFiSb/IgtTbWbu/WX4KMICBDpOdVP7C/HRhS/8fgujvvGYqKJu89cRkE5t/+Ac
oUUG4nR1BYH0N4zHcI0PavnAI15johY4j1ni0L4vKgZ9dsJBIpRfOSeico6/QFac
IxEL70czhzkvOlpi4CEz/Cm00DSVSVotaWD6Pe81XvScgUcyds2ouasAJM74F5A2
aaG7ayJNvQGxzvqJcaf7jk2tJPKwfwnpUg6N+zqrilfdY9FNhEfhs2MjEUoofK5B
5hzcy4RkbxUg0TKKgJUY5GXrM1B5CzdgqFtQxfYc/MHRjXDZkprjdnCbVw9nQvOu
QPnXZxd2MGPvLJPKRrxPY2j/kaknUy/Mx9ZgUbbqJcjTSjGoNYWYHDkWt7q98HUc
BSBVgzHJWURSqNWTaEdinc/j/JhuJ6FFR/xjgEqV/T5SYDB3MqAb0tTg3/bFmU7a
W2F5ErzJBVFWpQX+nTDi2UcUkms0jrLQ6WtrowSFJSsrNucfrtmrDDCyMGHE/0za
vEvN5Jymb13vXaWldxDj8fZVPR2orE0gEvgJdl+pwS/QA+y2l57iDSh9ciu3JsoB
HtSFmr6p1kbqA08JeCfW6jARzJ2w1LNW+Jnpq1534DDhgyVtbPlZN3L5W4YRzfBc
qEETszb8zOApiE1BN3lmRnHMUqF4mw40CsG40cQKnJ6fNgi1YAVRtiGtmDoXqD/k
rRUsYSOk9RTV+gNF0uzimscRdPLtd+ZRtau2AwrcQVQBoxA3mKK1SYR4XBxpjPTg
muGAvkOojIZBbzAaP2F3CUv4LMyuDiVO6IIakuKswVGjeDjhSIcxJ9+PR5YJcjJh
GEDnoUjrY6WcKvYjEDkhs7yabV0RY2gBz+j+MTCOhn9OythbDS4m7ORGbTQq/9tc
Qf072m5wZ15y2Cavo0zbZVtyiNYWq2YNBECVm/MVMzEMYCb5a2xXXNg1dcxXeho0
XATcz9uy0wJnRAYSe0KHyNlBZ8FGVVOYC77fvs7iiIglae9baokxrspG5bbIV0KL
rrLrFWxB53OIE+JxRn8+eHXaJfA8WmnJ4LEVzy/odAB2AqQ0PBZiabnCehQ330C7
VMfOY0+dQ5UZZrBIplqtOjK+7L+X8JeimNSxwG/Ysv2gnUuiDe2YgTD6A2ZaKLVC
dp1rT8usjphTB2RymqaqLDwjrzEE8o4uq53FiE7C7TLeLMhs9iiDAz5COXm6Dkfg
cyw6b6eeYufqxengNYS9Dxb6BsltGgmboOmrPpfJkVLFHUMq66INsz/TFiCEYEmi
X9aLtDvejcTl+yHmWuCLXco5oSOubl0szk2J0L+OKq8zuM1gqEShLqDqCVqOTyfQ
lPB4EZ1bh6830SRDRGSkZCoNWDZ7YyJkUAqo7B96OcMS5ipoOGpeuyM2bbY9fNnT
tKtfDekngoUR8kGGOWeBuiJF73E1fXB5Qb6fUeqcd1mifDEDY/5wLz8FkGOCGyhT
k0+1RzW6j5uj6AYVicWu/VxKIqTHArUlwfCr5MLXfCeawcgxa673WveJLshdxYky
4yC4UdZOVg92rPDb7pbn4k2LYd5Xdrn1AhE7t7G/L5w7b4nwGNIx1HNsP0sbV1DR
cDQJItGdIm9Lgen9yd5mpwkRzKnzr0jXdi3kmMh7w7q73CgRq811i20oN5Qn7hkj
o+DnnC2yBbQ2Y4CgYz8cjWHQbCa0gIaTouK4Bd/r3iskZfaRgEE2EsTWlw+ayJWa
VvlWlMVWLI37+nKUrp1iqtraiRKxH4g4SEiBLL0SGWv8k8FK6A1Z4PNA5v6QIUKD
t4PFyrx54mmhVexjOlZepkXVhLMc5SoeYnZtsumTSqTMAPg+9TBRlfAGihfrzhmR
/cBw4w4nzcQJOndO5uCuZmi1GGwb4bbHjXivS9jTdh1DhZpzMCKVhc23wl+hSRJZ
LnOAxqGcIKAru09cfydGWPa2xjrmzDDf+WvYxjVyruEaV9xy3p5h2HvOG8KCCkeN
/korOYz1vDQWdDn4aNu7S49VtMFdgWSqrolroeCND3bKYULa+kAAEQL3GCZVyCVI
wjO66qHDWRIOy3w5stevi1KImd26LzmR5jrjdxJJoGk46wR+RfouQT9ELMW24lgO
LW+62AFa1WZzeFm1AAfXB7FZgUKMnjwkH/djqXrXeXOf0S3S/qgJVXwmdtZyogwy
K4ictx7ZFi06Cd2hGVGj/A/FGN3Ou5C+Tb482TxgqEEkvFH36VGs5+Ws3b+cFyLC
CZGUMzZHYML5qQtTHmsIIxBY/RH1rd9G7Grl1ASu4yJy1pUNbvVpkzSBzQ2DBgXN
pHuvOvcucHnE7GX0FkTAZvFZGDKy8JozJdNRxiyWJQViaMjxzaYvuQLBo4/T6Goo
+q6Jc+pNVPUEgiTcdal5Af1y8B7B3sR1q01QA+uPkSom6Jvs7EnEn3G8GEWV38+T
8U+gu/Lw3hgv9QHciL0fv0A9aM9+oeIE7eYKU+3Cx/NYjmJUkJahJEdVxbSJwKlA
YWDMU1rUmPVfjYoGd8Xr+g7F/HiMuveFLAD7/DklqaXNqkTfrsb5zvA4rcufZyAL
W7no+vWvjjHn8qYDhWxK+xdai2n98D/h0DbRjha373fEoP0mv6rmMMbwOZn/K+RO
rMy0gY2HAH9KNQ7L1XK5L44npmc/hnT7R7HcL4ZDx1iptFB8BuCNtGdUnJHaxAt1
70Axdhr6cnDU6cW/orQZfec2b+bWyN2VgyZ8QNgW0zufdoB/AvIBu3I2XrOmj+wp
ntdd0svba3hWBHWhQQcoFcOpycW9xK559J17/0zLwJwdnPGTm2J5DwQLR6h8mRqU
+BJZYGMsOOu9+QluzPYj2VUGjrLV9Kjrd7MGf2Qe3suLJp9H8FV72TUcO4FxqgQa
i3oIf05byZiDZAWMsalzeTEuRlSAs2b/KKWlYOm23qeRv3WBLjkjgkJKYtmdT/ZY
nohxSPukjh51cESGTSlgFiEqZQNO0XUooBsiu6HDQyCRApv/7VOjxoB9WYqo4mWH
IIEmChhGuaGnVrB46AyDmAKeyBvK6/aVE2+IBCy71VxwE9hd5lGP3h5834siWAb/
AjVil2K6otf7eEwaAauNFMp1PulLoY/B2fjEnlHL2l3YYFXz7m192MfVchoO1DdV
DCHICk8gJK86CXloCnC+8TMJrAJjuP1o1cU7E6uE7X+B8qOB7bJeJILDlC5IQoTd
hNhDlOZyAlEYOzrdvmx8ipCSXNZstAKQBtndbqhFUG5veRpAQC9PU55YHoaohkFl
oglwQz4dGbgE1a/7htz8HhekP8vKHdM67n6MST28xGX32Jj/PeL98aL2k4h2+wuI
O9Y/7bWs679EQeK8grYWntU7wOh6oRfbJjwUaVKwcZ/on/d09NOdlKMKohgyv9c8
z9G5vT5ek8zeWSS/cPAc7bG4kEmqgUAwGPLFpzpZESDAM1n78XLi3ZO3A1MqzDYe
cgWfGZ5UJaA+d5xPqZx5QPH3brFQEMIL/4TZ1DJS5HhzR4q8qP3keYsAu7vzyStl
MOE4zd42nnaE3VQ3tapsPbt/PMbKpbMw+rH18iGt7Nhb6dLJtlroxsJTomDuH+0O
zcn+5fbYXtTwXWmnhi/e3hIoKLV5WLPGZR34NffNFzw6CrkUawknfc7OnQqHDOQY
UdJT4FiuKDzEfg/AnZZ8BlEL1dyIY6eCNy83jdfuqi/XHBbiupgbGCDW1KsrGh3n
JVwTrjrsenvvFKE6k5eouqhDltuzV4bbcH3ALk6ydBolsamQmdWgolJIn+m902Ut
20/RdlnnY1qPY7BvQupis0DanVve+rq7o1gQrirmKGKQaL3HyYOEuvJqiJseb+FY
/jqWadPuCvoKQJn1gwoSSrZRkE948/W09HB7uGG1pRdO/aPMLRYnmv5keUJA3cHX
iSUfjFYwgTcfaLF+pOUjz8kmmgmJdyOqYjHKbI9ErUPktnRda6uXSi7VABMza/mi
lfyyzcGG6wA5ADufgumO/UdkeWRajvDzHtJIPT8Yj0UPYFhxzFCkZRQH+yvP1ebK
vE9Il4H5ZWFuhyvnwMwc5jSygyfUUmuhp2bmtvUphFEiwoRO365vdOFCayodjaQI
LA7k3qgiJXcUrbrJ3G/+oJky61ztEwUDR4t2pfya7C8tswuoh5+OMgAWSqnDc3DI
ml9C0TP9TVobeWhEDh1T0RSbhaMJ9CY073LIduz6mOvb+8zfPMoUIM4Dy7h1BxQo
209ReCCySBREvvCHH6qZfXMLY29T4U/CaMVfcy9Y7NTdLpvWnAXJJzRZxv0v1gSU
EBjE0femeBG1XvglcYPSPSjDWJ9uBd95Qs8fz9xdY8PXX13SAluvAmR66X6TgbJ0
8j+GAhMBkORsznc+t7EB+Te0eGrqDrd0sh2tGPLQBYNfOUfujNKS1s6M0JVocTw4
T5YYGi4CHxA777pKnSRejz8zKVzOt7ifvHzA2VY4BJf1yF9A18Vq/C2QvNcHewti
FIDGL39veBkLkdxhtetG18YOKNTf1ZAscavWZ4OrRwVXvEDl/xV3pNnt0rIHzqmF
eLKzWdCBnr5Vu4VZuoxRg8ooYjKUXN7WEqb+1in9qqtBjcxB2A3j7AW5uMeCsf/6
4G2c0Th/d8ijU6TgAO6/zlIHl7ywCY+YXhFVb0GAMYst95j4EY0IllLCxN50xHLS
6QLVqk2pu3REUvePrVNQQI4EA2OnRBixPOpvRkgCemGIdeLnfH6k1XLZ3LaqmSq8
prdzgtXvJoeGcHDxBSH5pG33sWAqULvqawn8jVBZon9oM7YpCwUeYg5j/gEyYaNt
VEgE1ohDZloZce23KXTOJoUhq7mLeUnLQ7yumNgZj5pMsWbgO73xiX1lv9ZYLYqa
PsxU31ujFELxxMrAeWaSwAGVw6aEVoano5w9l6O5hzMYNetRCIOMMtohGFOVniMJ
oEjW9N/zxWZmTAEU0IteQL5BcJvgGAi2eT+YyU1WdyLRABCnBvRXTD7H8GlGd/pX
aAvazvPeAHGZnOgrlBrgLJm3X5NVpxvQvKvmMn09sePplLm811nsBadYDPo1rylS
AkHUEpPZkLVTFefbSfSbyF7hybmqpV7yNB1lgWhOf0SUMm3zk5Xstj9arS8dhzbC
IKEU/ahZlb+EPKul7hllgOkl7Ck19tocXDJAtYKyBnVfMCCPQHcvrE5hIwJbDK+k
OQh68SB7cQoYzlMo9ZoRInc7S5cyLaH04d8VUikzO/DPkq9RsOV/wViNyF1yDGcK
JzYZN9yvOT9V/rOuvf6mrGrpwbo87ufEG0F8i3MzlwXY4jumdYnuDC1HL2V4YDJz
Vor528NDErN2FL9FM3fbf3Te6RMwv4WnZC2hi+tws6Y61BQi585S8DuyT09JC3sw
W94QNPhDvk6uxGgXSvZu5FpvNlpbT98+KxDuZME4gzSib/xIW7L7TFh7Wna0Lqep
7wEUwB94M8/9daBWT1wk9zKY1b+G0H5hh5nSa/nBn80amHuj32nW6C1KGxSbpYsa
LtcxNQPgQfc0TPiqCZbxX6SZAtLid8Iilv5uzPhjeIeAIqKsGFAMBoQpcxxXLczr
xIHyKN4jpJMq2NKNm+XI3BcdXzTqwEeCpgGJGnyxr6K6FS0z3AUTewWbyIvjPE8v
z6FFPCnC9OEniWjmaTuYJqXnHUXeLC8uhOKT2tjMsi06v7xjkSFDGyWxoUmbSXEu
237qReNauuQUzmvFra9z7n8hpynvL23PLAOZN1Ekk43Pbb7MKQhcqZ9vA1bxy0Jz
724ZpYjui+4lpzrQXmCRc3+NAcZse2ydSlEhZdK9Jr4iZpDbj35bU3Z4Yqa1N8X7
DYT3dzhKkz6+EUt/BDKA3xEHAbjYBVoSIusqYIi052wPh8DdiejxaFjjCiw9x2O9
2A6fAz1M3mKOSfixtvCNlXDumnVlNT3yOSWVX9/QuTakyLht5g20nHIEaxkgMOBs
GKUB+kc4z6Nl57SdDBuys5iYvjFqVNLrK8pRnaSS2zGDN1F+w5pPNgfVQ1V5u4V9
TNz+ebIW9mfsN1hh/5FMh9uZZcfDNBCNwBEBgoqgwzIRm6cm07aypKHmLLn4L4iv
Q66B9DqoDcda8cqG/gSJMF/DeihCO9BCi1WYWeNv9Mq3eiyCsR5nFS7drG1x2TPx
w67FFVi9brEBrAZ3i90MEyEApz+DAwdNF3lazB83vwnk+aS6XAzjkWgkInYfIpO0
0AipLnuFuNSazNHrNN9EHYQtfo0pC5GLtFfTne8UBX9yQCzybbg1PHKhdlSQZutp
WHeD7fEVzaV2qaIINPyGu93IKZ1IWfn/F6R0g5POGfzVj3ePqAU0on+K9qBBEfKP
13u88KW+l+vgs660m7FsD/LvrypEEkXk9AYke2q0De/473CLnJ3iHksMS3LA8Qy+
GptSssTD4HVwnMbj30l4j7uK+NK6Q+jggd+2Z+BMfPVCpvr7hjACmOEDJEiRMbgn
lsSmG3bJM6diJMAaIj3Fs+Z7lwol+odJ75YGohP5oure63s0Rg7q8vMEV1QwtpqZ
qiZ6rfnn4JwOamD8fR8s0wWslCLNVTWJ1eauNb01r29jkXx//HcXoaui8tHhRhl0
pF+3TpEmIeeP3TDhn5G+jR5esPe5ukND+RJZOQ/nipHWnoAmUsI1mVUQdJ/CatO9
qi4MuP4qKYWRoc97j108hK9cMWqNrKBvI7/xUfkDDfQyFfJSFGcrNL+8VGRS02X6
2As9bqkGddYkhzV6UN1caJvm9s8zQep4mNxqFr8l/9QZPt3yAK7C+2blvWY26oZx
ICMpqWTfdqVt/efGhJoDUxt64UCltDbtqJ3aXaO0vicl6pFVEHrHomW1LJMpCLOo
IyuUv2yLTryo0/ScX7kX04HBHQlVj5sUYMUAYGuDe8v+t+DOZ4YLitZ2M2i9eyx/
EFGlvd8oUQAdD/vrAoEvZKCGw+r6SNK55Z44By7Yx3XXmR1pfrb47fO3SWOn15MP
HqL3gVo9agRcBSvRJgjINysxqKiKImXJITI8dZB+oBO3zzkJQBUvY1K9U/oRyeNd
nHcu/BM7ggHD7Onc7oh8f0yWDOxXqpNnPrC6DZk7cW4v/w542FyoHbeEsNXzfp5E
6WBTAEFKmeLhmiGlX7elXCP4IxQ9FqZyB2gRkyojGCeDduejc4C4z/lUPFfg3QWB
u83ii/I6NGlZQjF1uCWXefnNwA5/hHoXHMviCUwPZaei5+lLp51bPWMCVhRv566n
yVA4SXKVrX7+K518nY3ayM+1/oiLQTqqOOx47/V9cEXBqjGTL6O10+bxN1yV8iOs
ybi6/dkCrMLUIjLcXxQw/247ut6vxoMlequaD+sio7WkHams5DW01zYHKiH2OefI
YjYXRajSUX7T7zbyn4MK4LALXGmJccbYBfYRrGfFI3OzZUO7sY8kR3qFUlp8nKjA
JUi31qyvI+IsdIgZ9zOH/Lhzl+uMu3YZtykYA5KAwu2xiIv1cMYIylLkUjboDogN
ZjwNhGwrhmUKlJeOI/9qU7/Y7Jl9Im5yoofTvYFpt7n6S/fX3ISnA9PvJE8O6gsL
cJIFFs/T6wut67QgCNjuLfbVdTcE9K4LJ4z1TeNRin9eQK/AGDlZeq1ttFSbw/lj
Pvi7Ks6WuDdXSqGbdPG4cDuHGtI2jMNBLqy715Por3u7wUYzFh+q9R04YViM7+w5
YfAz7VN5/vOPXsARW08qTwiSehXvV6dDrtydhbaK3Jpk4cSgP9TTq9prCB6sNNJG
QUIvgQPWcqATSMUf8hGKYEGgc//j5MAqSHGx6v7GY+rXy8VwhVGgXCbogSyY6F0t
FcFrAsQ5L3WSj/LVzVYciXqIft7qrfCwqrCA8QdBSNkXHSKXYdOpi5rt3KnEZcWV
JSHDXwADHVBdvQ09rfFHWdHds7nDz2IVAT8cIcY+i++pX8Ibdt1FhtOtlbcAuStQ
qJCsHtT0GEnP3ss9t8n5IZmyMWwvWomebN5zR8iuv+pEbYOeR9Yw03k0tBs2MZOG
C7y7qxJFNC+UONn8BB3ywHMjNHVGLZhCCS8dX/u2TbEYPKBfHjaNnK5OxOO2gVyh
QQYHzwAs5WepK8PuwcmSuMcTISx1vpoF6JOWTLyDnz7yWA7ALZTdKuVZUAm+2tSz
OGl7eD9BbMZsbZMC2yt2bavMEOiIdwfxkWjrpN91x6wbqci4N6AY3o5rR2Fs6T6J
cCu7zYBxDaA4fQXyS+8A0TC/+PDZZhPn2T5G6kQ6ZPqwFnKogi8y+Zm3Q/BX5yud
lrQ8x7/4xbh2zD3CToz6DEedPjSnRl9jU4ujlPNSwT65VijX1pZ3RpwerjxDf1hC
Ifd2/qACI0MZgp5ZYBEq+cdf/pqMBcSVKnqbfixX+nTDptq2uSaMpyVXxF8AlXCp
hsXZQLJ02ieRVd9mOIYq3q2QnFaa666sMuBM27b+++xPgOrIsTYqRTsH+oFk/Wsw
sRDpt/Dmf87KKy0+Od9drzUv0qu4mX39ZBdgg0By0znIYO4JduqX6IdsMWEqIWtG
eF4g49f8kpWNTzcRs4nzxzUNi93pCCjLGasZ2lACL8F5r2JL6EG8hJ3boGg+tY+c
36q/CudzkybtyoODN7mIEUj39/LD3SF4aB9/Dk9EgL2Vy259HWkMwHCjVE5TYdNn
p5tP0dDHtIzp4wy8/QJdtaJMf7R6zIIKAYnGZtjFUR18WpxAXnfh9XTb165ECmu/
X7XiT0aDLweqyhwtUsIfo1bh3QbR+8a05jqBHYCW0YcL7RjyKIeZ+wZAGkzbZH1b
zalreWuk1cgl7Q7aSAYrxNV2YWihVnyYWwFCbm2mkHEdOl905/zadAwlZ5+u3l8J
a79/V04euv5x8jtJ0TIFlxiHK4mpLB87brHyEkX6U2icqiZhTYlXivE0PQxxONf8
zr4mlMhT8X/DvDeWozgxk3l+KyXgPeu2SMU7LdggAhQIXDRfwsJ5TKMe3KoJ8n/Z
nnEUJaSOg0M7Q2rnSQYxaH9/0+nlXMWxPDUhXOD3VhFLahSQ6HCw3maSNICMhu7u
PPA1QIs46qOIRExWJwdve4W03GRDORTmetK7utCUcXdIFSnkpsDWypNUbFNMLOTA
GqIOVovtF0uGva52TuyW+W0QJqmOq5fa5NcQh/PauRNOt6O1OkBHakMrPx4KlD0D
YatTR7gSDFonym71j9vdrD/EkmePO/QeP0rAyZAfBRhPgM00SnGwMrjyqzP06XbU
JnoyesIrhrC594NBsOT7gGtx4piGFHf9c+EaaSoKitDMmgDSSf/QNMHgrryV6sji
CXBzeUg2E1OVN5i50+BcndZpd/WDsKKdHvrkc0VccqFShfOrP/qZM9c9RJtQAFiK
cs2w3iwlGsJ+xQ3HY1+CwKSU7cWTfYwDGlla+D9f9yGPRt7Mqfz2lURuiC3mm9Ty
tb20CuWDjcO0gUD64JeMDfVgJ6+EQ8FgO1TNYoJ1fa5PK2n75nhUHi1vacZUwT20
h5p0tgomn/pNs6UWUyUf5VGXH18wXGSMQ+Ne+PMP2Wj+iFlAdjyzaThr2sUw79gn
wdVtCg4vG9CeqARVoB5wboi6Ju0sRiiR53yZcTLPAK+CZGr5y2I00bXy+Rlr8hz3
fVUze1l1jUVHJf0dVTDxP32NKoyjP7T9T/TQIaqKH4wzaLKX3vXFcsLgQbq+VoqU
VyUFwwApn0W042kfzYlQVTmZrjmg1tEUIjB37Pr258cX9y/2kMLlZwQcS91/a8Zi
re68AObWfiylKPZn/0Rp6/RpTH4knpTgzxyp/CFWYyBrlQlcChKe9I6yXn8GO9y8
MEcZQVs0B1YkBnrCNDRR2XI9HatmbVlFXiHGd6cWhNWj1bhCP9oHglqRpgt0K7jJ
iYYzfgiTDNc4bwEiXrPJObvcDQOOHFLuwA1zbzDm4wJB2BIB6XYDq9xBg3DOs6WR
dJYHdToafumh/dSoxt4LWcTUe7ScJzNopKgjCHWr0S20ylfOpfS1jGhi5hVym5lZ
R43tRNweJIg8JSCCLYDmYT+xw23hAmsa5ZoZSzTwxuc1+/ILzyT867deWUa0is6m
sJ1QPH131Ak2ILa1CDQ3j7G6uNSxVY65+9qi4eFyySGnPzp445gI/sUeQKOQTM5o
JX60AyCmhSCLMkAhi+yumw5LbNxEqt4AHLmIh61F7gplIjUPIuvcJXReZZXNCmTQ
lZ9CFqgjlhLgUIgKUdY0QSr5Z8cYART2wAMMK6eUY+ue6ncOqw0Zpn9TUdadseHB
4fMtEemcZ3rBwyZBINGhXY8kIXOemtQAO7jyNceLV/hCcgGix8zAeWcJbe43gOXM
lsTkfo7ag7BVwJzxiVABW6jgUYuM3YHyQzLUz/ctQesGMRlmV8cIda8JNHYQPPSs
tGXXAi2ZwmHYRzFN9ze7z8N/cTWbOBs56ASESFW/6BUFoF8v2sQEubY392kMq0Sl
WSkuKx4kQmQHeaPA+K0bCBILexjDhOYgY69YuneyMpKCHg0Oaw6DOFC35v45N9P0
kNkcI4lcvXe6mijJXfxKpHPE5mPpIzSJUNc+/KOkmyxsDr+DTWJTIZQhj8DIxAOi
75Rm7dN5kk1Zl0mtEoeXNaUYovtHe9zSUTX7PkJjPWcd7e+C+HFrerE6HdxeeWd/
5fIV4j+wbVJhOIKG05H0GfLvZ8wuwjACBiqW4pGt18qpKB8s6pACD87vEzL6xtwV
oGRH8IVJhbU/sbtITgAODtoQLGlt+4mC8ibN5WVp02J5Zp0SnOKRNufAtCHrp/AY
UEJ7a7X8AQgH0tfsPz8ie9N1Ob+vCz35/Ecpoiu3leDVxY1GH1VFg8NOKDClhBn5
4oE9WRZLjEdCzzPZq0PO29Ut1htajRqpiySOiMjFJGFgN1epznwTTDzryjU6IAz1
S5sEfzsxDvyFNgQtPan4rqbm1zrHqwAA8P4r1KZ5Bt3ZvkCick3OD9pprkO/UKX2
W0b48osX0HKB7IBILP4nENzcvtDfcCOAP/uiFm2YcX10au96IC4SM4KUX2kEZFSp
SeNSX/YiF90Ye/TwKMG1Kwpb4FtKwATQ/oTeA09Ur1g61V7MMxCTOqNQITtivKS/
CrS/hLvT3o51NxsvrbyQzdDKd9V6w8vAvu689fJQMiAhQBi1uSzmejusov7ix8EX
WKdFLRQ06t3KhGp8s/uuB24w7XgKqiYGE9VWjtV+GVqTHsbdSEcDS61sG88nxc+l
Obbmq7tRsLkPqLiztGzjMpUO/pKwkqyXTkxhzYphSuPtKNcETWVCofONXI+bgN30
VcfMfiDKNsIMrmVAp+vxqM7/wixMzeWWErTd328AmLhp95sZBf0omxhAaCmbjxvS
PH8aXDAJNnswrwMZZKh/RD8hKLlvbtkPXVNjgQSqCwt33s3xdFvrtMO1XtoP9cQ3
k13KgcSAifqWWdt+VhUFBgkHWKK0wS/d0ljdlF2sxS0YtxIR3pqQA4G6px1PFr9n
nTJgZY8U6RE3RyYDLJzZDzxPg+tdHpDVg3lEdPDOHsbogFv0wZWm5gIbIpIlgMkM
dW+7mbZErjryvWKRkJFGjdw41SbTcYP5swhseROu8/qpIecyh+DRznVbf70jNfnU
b6EWWRY1CQehOWumGTKXEvpy9cDfJ9XlfANg9nXOQ5wSiDyoNdfx8WjpujgqqSzG
BqxDqOY2/nVT2KK8eJu+lw5Jlq79UipKeRWPmOKYR67ezsNjLU8RtxDUTNIHZuto
2igLSiSkVm/UIeU1tORg3qZKVXxZUKqwwH37exswmL3RraGLkZIls0fOQbpvg6Ku
guX4WbMiLhrWZECxhVM8ev+YeTbD2kIr+4rr2hJ8mtp64Z0OdJsjoZQRPovg9K/7
TU+2M4hCbOYky4/waWqkCCtycLd3PPHCUdir3wIzJVbUFlUGjlOHTbU0ohlvYp9r
36HsGzUbS2Vj5fJrMoVUeJmEt+rExmzKpLmH3OnG/cYyuFXe6N+tE0CNAXPmV+QY
J18imQeuNENFuUHUIW324ByHoRcbN+LsszveB/pCvW8SfTFIKO8j4BOWXEKPHuJH
FPIlsiNNspKOYv5VH/DhBMUyhK6Ryq8JS3TE3dTrzYLgXMhg7XDDUfGTMdtP2jj/
Gwzsmbgdz7Ag7rLJSHt94Qzvb72A/rBJ80K5Q1TduXSrFsU55w65NIj5hyGKAJqN
wqxiH1H5R4eOg0Ay/MHmozoIKnDXgircxKdroAEL4jwJuHUdnonuszekbv89NF9n
gSSM8901wp76UFIOEsCEIvzKQzYjNiGArkxuHEU8hZY7z80w7Loy92Vh9BManNWd
34jEd5ubGb8boFMSbku/uaA8MJmQQkLy1LddV6f9Y67cohwUxI1LSmy1g/Ej7XPE
eskRCC4Mc8z3twW3IZmdIFYtSYEIr8+sac2UjfBFjj6DrxzFHYNHt7sAcUPGKr+E
C+ZFtYKygmZo752alSLs+eZn/uUwGWlvacijbonDxYymsm2iTYhuFN5gCg/UtBvF
8sMRWOCHJjFwGs8mw64ffqICbRyVg5PjgQuSEL0h/W4GGimY4K9Ajxb7CWJNv5Jf
n+16T2ZLuoQDTjkqdC+LCNVw2jeJOsACWw+zJ0IBOBip7oX6+9Vxa5zEMXXaqSNr
QzckKvWh0UShuNSKsxqHjmKsZG6ACKcyrNx5lT3cFziMv/uV8U+qKGrkA01thStA
BIljJfPsSVXN8HGCFVgYnMnXdKwa+xJvhePoUkYe2wCY1k6cRX8mrsHUq1F2rCj3
MWUBuD0euBSdpGfmeY7uSUto4HR7nVN6ZcXXPQ9MUaPp3HJNYdZtPjvzt8VHMRix
QpCqrqnRyGHNOzdDug+jX9+IWleFNE7QH+D1W13bTQiYGlaJfcDKySmVKiZYZz2B
UnrD5Bo1+76Nk6opruUmLWiOHRZj9h2uoYOP+hPnzrWBRLSXBLvgX97g1uKgAoNN
JDNOeyg2rhFCW8sRZ6cDBk9Ys32sS3XWpFh6fzZJfynbINHoOplMH2wTjSMGJyGa
3fn9gMyBZphOnnlGTrLTI1CVkM1VnI5FkqoiAByq7f+nEI+9DvNgVCMcX8GYtgTi
0NEdR+T/I3Aic+z1+ZjWzhd3O96AFnZBwFwCuZexnB8zOt0TPaMTwkLkW4fgRsr0
VyxK/NNmsuB4y/hbnuok0vm9Y+v6ZBp8mk9JJMn50m1LC/Nrewq9m5995Ngp5DJe
Q9h5P2safi6Uw9jj9C9Sfp9YF84iHJ+uTKCw6MAF0ZSg+7eb35saZALvk3a7pVYO
LcnAADNTH9IvAtqcpQ7+Q8A1S91kHbgr7Yhh0S9A9ikOdnOFJLg0Q0l/FrD9JPNB
dXKjd6dLYzl9AkVsjox2fwDTQMgeh3MIXoYYxiKWEGPOTFCdxqxjW7M1TqrIADOk
DjMzJnExK0X/hqGFN6n0kSgLQVdBbagEfGkUqAeYMYskGg0zHXDbD+UWZllVnKFh
uxnI9FUFyXhxzCTbyTU5wDwrgMiONBq+/9RP821vgwm8f9vim8XOFufJMFq5Dt8a
Wo1hjJHPqAh9vPgB7rvDiAG9RQmYEhRMPLVatkhyZe2JTAfPzarSK8MD1/SMjnwx
LEZN2K9SaeDYlsXBGtou9smPXhb6y2ZcWlvnR8ehdp8KV7XD9me+P5NN40gEPVPt
js0PiVbuw5BTNpac+dhwhXdKUJ0Ay41Esfy3hNMWuC97Y2T16XPsZGW9prWO7lpr
QpEtilD7GDJDwdM9tREIvgSOOF4/HvIAof3j3qZg9agDcGN2Y1V5u1k6set30ter
UYKv0zwT1nZOfnuLbUWGyJ7P/iW056mDH8jSqoM5tvLAWZXPpcpdAwzMZlyG3nTQ
7Pl4wef+KvbeVZ/c+EpmxbBCMJvv577lEZd8ngLNY71sHdBX2TWfzRXo8vYa60co
spz7IRcj7JXhpCwaXl/m9YOu+J+vRO1KC5SiOktbkAOQdWwlV9w5ErLujDzvNxIV
sQfWXXrSVXFiDKIWsutn8xgyyQy/eUiq5vaIiDALM6i+QjL8EVdW9gVnxlgtlQk7
vapKjh8fbcJY2wnZ75JevKigKygrQZU+VgWkpLjc3czqjoaXn19lEPKwKDYcxpvA
nNH8xEfvT4Ki8vpvNGx6FfEq8F9U5JYvGgMqjzzuxXl1xpLdDoU2LjkMGyQL6kTS
CJ/m32GwX4HwGs5ipavgspB240naWc2ayUVfljBau1WDAjcFoyrenaqPYogUo1Eg
ha1m8ewX8kIV/2quqluZ50nHO9Q9SVkKedHQs4etXXV34PsFRe668InagWW2FKOR
jFmpd4gStIqV+jlSxduiUQmtQOhX2LPaNp+Cr4dBjvqBcbdj6lhcn6pcaSLrMSe/
W29oQpn2WVw/ziwwSVUwL0+k1i4sP8ZuwktHlqTO0rLtye5BDhyuMJSzLM2rwlBh
MRZ7L3swUcBwGl9ptFD9L6ZQ62FVS1tv5JTaayd01Edi74aHvHDKUYpMXxe/yyxn
5nKdBpLH/ihCo4M+ujC/3rPxJHFthjxkGF/hkd/CVA2JXbPUc8TUmEJqXc59WjE7
Fmd4qXEnxrqU625cRhRszzz+S4pHdjTkKdnNK2R0QcU7cj6PJqlS5fdGim0t08pa
Xfe/w/B853OWiAECIciBejzP7zlt0jGcU8h+ZopoBBvrZSQ+Hp3ACLl0XOD9SEnJ
FVQ+YITkCInIDaM8wpaYX+nsnBms2321BC+i/Dw8G5je3LkAMtBSezLG6/Ay9Ghw
CWffSoq8VwJQWxvahSxryd6GlKuDTAgJRoFENiaJ9DXbLdJzty6WPpNidOxG/Vve
wbY1FmKvHC9Ti1AQYAGNpJCjuN0AkfTHgwXgdh03zdhnjs1pQM6BEPVi3I2PFTFG
ODsgkiPXzAZNXqYWsXd26igGmKjvevIvodJ9crAu0aBcn32QQuHa/lKX7u/0NKPl
16ekJAZvHi+rbBPa2R4eZCKio41TeJvVaBLFQ8exZylQtkZbTLeEMLvjP3aBl2Cc
xopBsRZ4yimXTVZxVH0qZLE4f1+lNvhKsC6l26hzi2JK7RdZn6bD3Jv1/9WY5KJZ
hTbjnyV5tYaltEmIL6f5ri7GYpXkms4JmqidrAedtUUuByRNe/Qu4OMPqUo6B0XA
OkBUe8KCPpveHr3Si7KobpXhBmrVyCRCqj3D8+7LMK6M0t5tacUJdVMkfgv9Vxdd
+Q951mS2JPN/vUVRgUHQCk6wTzgscRjEVS9XrYz9Xsvow0shET2vQTl7VGDlE7qX
2SDFo/STYho4MYhg+KXySSCZVzpFfeOAAY4fvu/ARkV4fUdGS2OHj8Ot8RgHzn8c
q8PNbAXiT++dT/7mNzbF3TKtFXwsbec6M8lY0wjgE465aw2Oc2sOFdEb4keQa0QF
2UXBoM8aExvK0u22uaUdeiaLfMJwimO+4F3WtU9syhZ6vDYx0GIOElzM03KiZ8V2
ALRZFXuzzvthSTOmolqQFXMjJCGE9FbRjpvTMRU0kCu/uuuEtrND8BpR6Pag9/Wv
nYcNOwNa32lJxb+rzg2R/FGsrpmHZGsCztxwRmjP/z2iF12OgPj3XbBl/uyqoQOl
NlO8NOBa7SJOUJBab64TN93mRe1dohmb1XEHfTS7hbOTnjxEpy2jM2SfYDsoi6Oh
0nNUaWYyOJRDPABrJ6QgimKgCN4dFAC7ibRNP0MXabPbC9BUVakoh9vy3ScIVdcn
tXHTC3mxDnTcRxhuyqWZuoK2KiNCBoaJyOx0oXGWXkqNgLxaS+uDqxaLcA9+OFWq
3g7bX3qGUhtU4jxsv/PzvBgfq/Vc7UwbL9cHPYAWx4TO3jJtCQePO0oyEUsAo5SH
tgPT2br3+HkVp6Tf37GuPtIK8qF14GmKEf8FewWBrfKObzWSRG0gZMFLZWKJK59j
EbA8bEXmW+PSwW4P10AC1pDdLGVFZjFG0v2pknIiSgb7n+77k3LeB1fr7B11ttaL
whi7E3l17RDK8yqtIcQejavbC5KSyMjbteq95zMxG0tgVnI871Qwfb2wHl0Bsqed
dE6uFI/McFaLWZSLqlydSqbopFRiAWrZdiMElsEMLOroAZmSCz3VMZBX9PXQjfop
aWpoDeXShGkuzKGSF8unImdQB0UpRUAljT8kl3nFvBdGC/L5VCAmK5sYW5nxdpus
wEYvTY7tbRuH+AZcLcEP6dmZfz/ouGPZLwLCQS987HeUv3hz0CK4yLPifyNln6hc
xuFYO48JU78Ov7QjrGoBnN1+K5XhxFUMrnAhyl5TABrSKQpsrS6142E2/e4iLJlB
Lm7LOL2jwKROeMlZN9eK8xt2BFDh9FGVn112cCkCjvgaXaIUToadvQZ/ZL2f2nq9
aWbnWsdqWdy0n6b/UT1s3r/asONK52lP0QcYAtr71mf+QRBRJJT/IP3d3612+INV
93hP0FN0q1kekobU165ccP1uPbOnDZCxFS/PACWPw49CNQ75Ve7v5nvmuEYxtFrB
SSGUMfc55mpI7XoFmaCxMJ/IiEa9oXq3VkIUNljyVyPI2ArM2gRuKJ/I9o42VTtc
Wc0qwRAx+l79C5XJnLBKmaysFHNPd24IcS1uZiG/3O6cF6UbIMnrwfo9NxVzURRR
YT11tuVxNWEi5H8At2Wv/9lLH+G1G2wMoFhpeGT6tViCyegIqmrNbeJ6Zkvg//7a
QPMWr9YolMSbqdJ7oF3t0MMAQuv09FswzONdgdJuh4LMidSxpFEYGRb0qfSmzh8a
pNiK+n7n51hXb1IZySdybc8Ei5ttPvw/m3mRr1jyBNjtsJxJUUTLV+lrCY4msNDM
bzoD9EkC3+pXV/V5neOx09bD3atuMqIL56KMHcWbmUPIGvzqH0mOxl5onxVTmVIQ
dMSxqCnxsQVPOd9NXh++1q30Pe9ePhyNrC5HqEgh6SH3Ud4S6iIlHOeTLIjexhEY
xm4lCWwNug0cqnO26dDi+/cRjWrYFrf9LImauVCUzgvafqzMIm4L67Lu1x5soUVw
lpMdBLfhaYFRLEAe3f597r0D5PXbIIsvc3LNWGrB2xIgpFzS6jIAPzPuXtG4Xucz
9nZZI/0ObBbp6tVhyHWOA/tZjokmT/bBdjhpxW+Wk4Z8nLiRWK22j9//IwZKlqW+
5M4b2c31T0kcyjatHJfMECTXNL1gMcyTnFEhVx9pFaRiwXJF4LZ6JiG0sgZdYds8
FjWj7OCj3wnqi3cMItS3/F2r2+9LBuFncHH7hQwPKAFgdYtvYV6i5n1ubPNjo2wh
Uzoet7uLyKamWBamV4C4TYHXI5oEccCMLSNt9AUmgg/rK1e5m6rbHgnZ6K8ImGo2
iC4NkIZETvbFajO0WW6sYOFS3WoNOx6nGZ2qfP+qkLUJtmlemALIvGPl/CrJc7RK
4ihYOYpp+Mqw/gik4F7Ye1iYYNWJDbdIh3eZUShedWoCVoA4A/lPBG1pzR4ouS2U
bXGH4EI5AMjwIzuaQZdOBMbSf7PCyETNtaaEtI8zsk91e3I/ggGilMcYRewOKQb/
kNMJS4QvyZN+RGcG4KtDqmLOQlmbLfzcAwFmIku46VrrJ1c0ECn4d3+/zgH8dw6u
vuPzHc47iRBZjaSaLIUqoxeXkKHvfl2tN9n1+rhw+oG47lGcE6ey06pA5AbAWeh0
d89QMDN2D1U3Ia2vEQHhpm8F4Cb5Dxv1Vn7FgpRJ5keNyexGtquRA3uQS9TWMlcN
VAAkn/g1y4RRjXFC/c1i59x/a2kRg/tMgOpdJmr/gr39eo03OLu1/MNoAEWHQsBa
ilv4VlpZ0W60ZyNF3qMrJW+7E/IVklLE489kNauMsHcBe6X6FraKmtJ8nRnI5Zm3
yNlBQCg2hfuMOWE649VfhmfhrUny5+TFYaa4sd79Y+4s2Zk0kwXhYarY5zDrsw68
q7b68jCXx8Ngynp72fJa5VDPiOuY7CWadTnJtbcGNjifldDbdMk63+J2ooYCHiKp
Cm4DNVkstjejnujfiq/dBAFtAnQZMFGFywRDCDQnis9XngpfNEjPmVuaEXBOGC/3
y4E3t//jb8ImQIyAwFrtOsU5daM87pbRGyIqr1TJyPQIu21LY0Uc+h+J9DUxd9iK
M9f5Dhv4TikJ1wboE6Ec5NQqMaVK1be6jKbgykzJ2jhlZ1hx5VZYt9/z5J9dxGfx
2x7iUF2gg0z/vu5myIpKGEZbwKT2kBndyGMQvmKcibqtb4W9FgrZe5ahN//RVjEX
LmqhTxj8Qf3KrTC1UHOpiTp9Adg/CKjUVDyPmXiJWXaO2wEbtyB4MNTC8jKsl5pf
Leseyu+dOP0EJkKywpOYvlxMC+iB402VfMPKqt8+xJxFnQC4MM57mwVblRb6aEQi
OnchHOBGZIAOPbLMitQCPiCzuS3+q9TzVZlJe9K03mwrLtgRnLOi+OGd/5Vu4Gaq
itZ9Hq5gBLkI9L6cN7ZC/2ojU7iCwPBAHfplKFJb0TZ6fVDFZr9l4bQDEc91sBH3
nxoV7xHkf4IR2xwuquNLvOYyb9a2nmQNe2PZV4ewq94WuKOzxrZcLIqkL8azAHf5
ZH4UDqqme9+K+RdCVM5C5PTyh1R70+WXnQlFKrQ5pgWUfb9hmSxydJAx4o7kGub5
W4/1Gnp6VZQymMbrxm+nJ0xxJEUt/lelhSlujkCm40eaIBbUPFJ3PKLBp+09r2uI
l+fBHGKnypZ+Yi62qRCfkLKy6W8j0TuDt0pXwg/RbY77mLN+ldXiR7nKTqeliBTr
8ms/tQtIUwZ2GOZt1y6KnaCuFOw/vyIESb6GT45/TpJjTV0SL/4ZJNgcrgGoYjJa
McHPP8z6UnXHDc4FeJXclLZ9ASI4e9b640QmhxmbEgd5BKGuxuBkhhWR3i0a6cEZ
EaR8ULoW8bFU9QYbYMFXOAAKWypjEWglgrkr/RraOUvnc3xM9R0ww5uPzDzfG565
HhtMXEbcbLo1BMmKz71Eso1Mzp5EDrXu96Le3aQsWDe7AKnX9FYqChCs5n72x13i
YILblHyxhLLZ3/LnnaqonhDWzA0Ktg8QTrHqHD02AuViQjx04nk/LJEAvTng/v/a
Igl9zJR5SKbbU9e0VuRqIx5bs2RWvCHu8XWudQskfTOkd8RIg47aNTi9dDSnI//3
pnHTQbC+ShTdgLmvb8tHPLo5ua4O12vcPNTnFER+iLmse8ISVB0kOQhlPOpBZfda
GuqmQ4eu7wPQFH3VyTNC2ALWxdy56AK8RuEndik8BTafVFeSMm+2P/V4T/yWuP6n
bRvos1MybgI+lx4LcSsOEZdbvj7ySwbteQTFTAFuVIFpVKfcVcVKClZd/TlymCc1
4c05w/1Q4jGqeihkHDhoruyEzpybiaMXmcxeNwBQBqV8KxmlVXS//dM1INhnzRwv
NfShmkWY0RVRkAzR5uD9nJf2WHY34l4Ik1LDeiK+FiAfpLc1GUEp9LL9OG2M7x1N
UGaLhIsoWkPlq3MCzCozMe53jCnfrNh9oyrIDLSfegVcotwnLQDusEmdlrM9iA65
dIBiZs3jBeVnM19pr+JA0KY6D1B5V68hVOFjt8uPtBn1pq7CSoLI96yTfeYZRDVC
mYscsOyuqwWXWk3UbZ6+yYAmTJd/54wePJmq4CsNrlJ4DRs4JmAAQ6ih4LaMQm+o
ioNhq+qyDJPOV5g6MIeAtf7RiJyO0L3/tqIsAGThFCKd0dYFB9TakfjGvuh7MIcs
CPDoxPdLch5Lzxh1gkh9VnGT6pIFq0n9cOKUUdfa3mIE2+hF2b0K0tAOpyT1mu+c
vzXGXmGcTRf597Ji9pRCUbjGzSzG4PI+NUkAVjz//0VmrRH8vf54DGal02+9rwVZ
LGv/nBX17+qVnv1e2jbY/XAjtS1m1O2jhDl0eF/hkSu44jKctgwx5kJexyQSh/po
0C+dcmjxrxI+tASbGEpFvXI7Wklue9/YUI26fiVkBufiQ3akrDV7VM8fqaOVppmD
kqTPphkHRifwgdDgcewtno72Sla/cXrCPIPMpGVWcLeJLRypbH3IWAQFvw4fPA/o
z5WGxD3QBfuH+zRU25vJdWsSV5TRDJCT5nB+3q4HLBEf2pOMEtQDLL8t+sLKy+tE
Yqa9dobADTgTffpiJq3FjaQ4HmEfNgS84TyDxnPPXYezglgOJdfi+Bd93OaVjCJh
aJ9GnEGnbYRmcO9z3Jd1PByiyoh+mpAl+K3B43jY2iCWfhZRWRC6GAHEj0IsRVJ4
VieDpYr97LH6xshjxjcePtwUutcD7W/O3ym/hrw7UsgVZWL+I08OIr6hjJlvByDr
IX3YYov8GK17hSf/kj3w0tVwJn6JNh+mJZaiiamsfpvdwvpjzNMxLwxkZdh4GWwg
Sdd7HOBRC+DeRPkHRS3MlMfT2np35wF/0zZRL9e/+jbwldF3AmOuUvOQOIGn2Kqj
YdxLnz6VqDwwq445cDfAa441nZRbjGP3PvURenOvXZMynedfmIrTJRz+CJbsM+r+
d0qnQ2v0MfauMz5pg4yKlxXXzj9EDZ0dLkZ49eMySY2hB6aBt0sNkG20cD/sdoLC
h0Gagrz9VPZQtAxFE2sa4b89vRXgCRc2ht8CMkX2BAWEFt2KZvl9kFor3qDRqk3D
037LX0bxxuXdXQavF6f81tUl0HhZ0+ndXyTO0yfOxDsTM1YlLdPaIEzRuvv7assM
UBqQI1LQ4S3U976alf2n/rrjWFX3Pv2iEhvxiquSIbGXhsWGZymhq/SktHgAFrFm
Pb9TpZDifUSEnmWlNT51NBEjtVpp+49OaEr1ti+YFVYs4nYkF7AdTVeIDUFRK8Bi
LmaiA9R7fZPVhswVPqIqRRFWOVEzUfbQhlYUBkyuBNa/e6LpHjtEvJa5BEzUjdGB
+a8/lECKMD2loFRavASfdHlZ27TZPOTsTMs/MNydLx19EAEtZjAgTUwX+6LqmnC2
hKk14BEFBuEb+1INTBlMsc9g/HzNuP9yBsSsbicMXg9zZnNKlpINxvnYfoEIEX1O
6dsO3dnkEJ0LdOP4UFg8NcJRFLi1y/Zn5wDc2mKj928S8XxgCpU/oCy+ATLKlnbz
zHBbVhsalhrFGtvfPHt9jNMhW+7ZDIq1Xlnw7CLD7tx/R3PwA46t7E526Qf3/irW
YHLlh4NI/IGRv9eFtJXpY2ll5rMChLd/KjNT1WD+VuW/SeciNdmAsAj4XIL/JPKU
SEmmhsX+QKjQlXhcdsI5pWkryGPudrXqrSAJR+KC4Zir3tu+n33QihTgB8qdsgFP
czD+vQnNlnmMfy/y0WYyIYYakMOvj3HiwIa3bbtg0x2DhM3da/FwoSf1ydV3WtwH
B3uaZe2daAq4gZb7HGyd2+eREQsgPr+e9hDhYSoiLY44ttoc6eU5nlfubUfcT3EB
FtGBs8pHGwhXLi58+ZMasScs51bM2SKWjvqW6+LxLhsgN5FmTb0y9Ws2tx0iye2O
EGZwinZnG+ww07C5MnRou61U4S8zMcPjnBgR3P/h6So19NvKkmxeqrLZvQTmKFjX
XsZnhMV59kM/0QqPvF2tIuICcXO+IqKRdYD17KDNMdMcA9J4BZQFCpxEkfVvkgrv
RwXN0f3g544A3cdkfkavOALLB4LpMCHV5va+wBqEGRV/f3TfCbRjCwjvu2PeRZty
xoPr/QjXgIyAYKiuZmm8B/f/r3OXdVOPFiSjfWoZaxM2B/erW97M+zrEnXLr00R2
AEp6N0vb78ZaV/eFaRk7IM5c5oQ4h/Rmy6Rf7TxQ09DE18lDBik8N9wbUiSbT+ak
yBB2o3PAGHr8gyiURUC61+ZxOyoz2jtpe0BAB+qnX7ujbQVLYVsYvL3AzQUvIfrp
uZ+OgX3bmz/IZOkIRfVx3L1ihCQZJl+/kV5yypCTeSBW69e7bAes6SxoIYTjNcJi
ht7X2jzDAOZ708YsWtgTEo3Pr1FzYaeksur3ee1aWMtH3JQII/YJ7bmddQ84SPSc
rP/LblpDJlX7cTxCgeQeaQVBwToyCHeMVNNN1W3ZPtXWYHrWu25q/gRS83OsO17W
WuAQXuvT89fNjG4AC2y1PQZpt7Z71fk1ATolksZM1RNK5PuavQMTKcVozP44KWyD
pXCeW4vOeExaAU4TdqiTf7viGi9/i8b9E9QdrKLT+ngP+0jTVk0cHF+9EuyLr9qb
5e8ySV0K7nRRVTeppzuvUDQMj28s94m0nXezar3U2cG9id0rw9VLQat14kfqpxSc
vW046ofohCbVogOMxy2NnO/L6M2YUO/81thgtwi4xb7h4sbBwyHOJxcy/WrnFsFW
uwTaeTsAHcyzX1ScWLe0UsV7mU2rCXCwcyWz9/B8NIlqn88+t75KV652XrtH013Z
YzyvT2hFjOK9rBYfLruYNw5fac6tDSsvO00tjU+lid3D5sDxUzhVVJQegoLgp6XS
ivM6ftb0Hc9WAhvOTzyBJyk4YZCt+B/3I++eT9qNAPgNE/TF9vgviJdhR0eUHIle
nL7HIKuv88yzCjZ2hxbM702UY5QbOy+M61hZnl4S+ymR1BMU4Zy62RTqiSOAjMOz
k9+z9Nj7jAwlRiDrTOkxE4LRiRUFWLOVN1fXm7PKbnzgNLzJ2YZTFnmzDfoUefGe
dnAck3YbhVlrhrBnWE8LYWsPVEG1lxySR8pkjvrPqvYqW/75guZ/Rh+PTyz/iZ5I
SrsQ3PGxidC/0z8y0bNH7SAsZFlSvoEvAbU5OCTFuk7q0+CtR+3e1YsJinwjMyNF
k6274t8krRJxuMyvRFAeaLuDmApusjR12RB9EDPIrEnc26orRVDkkCPO3rzx6que
P91AZkYXEbJc21g/KaIS4P2oCiRPoLsMwLYEQRWt382a9z7IvBcx/vcrzuWBkMxw
jdtwKZqon6oTO8i0R1ZofHKs5Td34qvdauOSw8ZGNuCUn1gE/mteATXZZB8AJ5AC
jYreAqL0YAf2GMMhcIbTmjoisnfMR2cChYbdVQQ4AVc7VpvSB9fpH+RA74NhLOFS
weufxrTOQnEWVPoeOuFLLV8eWlOjRafDkI164ZV9oZBCElHpiL/1Yh7Vm4lb58h6
1P344ZdyiRc8IghT5CzEwZhlgrRkNsYo9QRe6J8BudL7ZxT94xQNZU3oIGfRR46l
rhPgsCtNxB33HkUTZ7naHJlkiQIHnH2PghehGSU+06Smvkt50V+HpDKY+cfCi20Q
xtZI3LouVjCY4Gf3Y3Hr3mZCuki9JzOU1b2B+OEfMlW6rtMN5KjcPuqu9r7QwjpQ
eMR2tXKE72DGWwRazc3kM5smlKzLxmoNTm886kYf2IgpK1ThuQwDy8RswMbLcgiJ
cETRsqLrRgAZsYEYF9LSV9ORxFhHG5EG7qORH4ShHv0xbNh1AEseqFY/IASqKf1a
LZj+qUUyIan2amw0y9cO2CVle14BbrgVa95BHuIGlBVi2nELEHPcOY/CV4c2HOLk
CADlayn6FY628M6BBxB6KN1D4dtZsO/mWRxOxe4JqYtmzvyr4iNkha0Vl6rCvaMO
y+Sh68wnOrWkT7UFz8+nX/BBSmpujRorQwElVkIafQ0Lfl+516n3H/Kv1RV5WM62
++Z5Vvc6JLKyaWk6ftIEepzN2UWvkhAO47lc6nQG7A652LiKSd028clnzEF6kbOB
ud0/6e0yAGIwC3VShX++OdxobKj3jLSOwpVYvLtAzNIVXIp0ttujOHGPkHZesSfs
gp+JR0NJXrQ8MMhsBcw+imI9S11EqwxfYrdniG1/HM92Ud2FoaIS58AJN/CdKm0w
2zCARKFaghGHV0pghWZc+ayGJxJf1vXE7RnJUyHbUlaF0ojKwtzcms5AV+SFjPqy
WdLivVrdCfDQD+fAHENk7O9NhHmTXmlMAzPeLBMrEFI5JwVAPGU/QJKRh+GcYT5S
OLri3ULM8JWDDMGTnZvSTsQFjrtOW+Dx3p8MMxWxUv1p1bTlJ/p0M9QRUjCABdKq
HzIGZIj6Q7Xt7Mg8vWTlWW5sCO9XWL6SXeczfeThPQw7PNgyLWReUpKeNtddzft3
mvx6RgH0h4JL/oCb4ppqRu/AbCle7i2MNUam9rf8JZyCQme/EkFHVt5IowtchlAc
MgS67gnstB8mW5H05wG7U9iiyFyN/UTTTaw+g3YeDH7eUhaDVfSYnRrzTjx1mY2F
yQCzmIWYu5AXwkmRaYyIvs678UdkFHc5mlv8l/cKJGN5bVkxmSdBlaGUkklPJnP1
uGd2uSDCW1FGUeBP4TjaySMtrUkh6GmbpDAi0cruX2ZG4RiJllBIfdMVJruvQd9s
OKc8ShB7frX8QNwioq1Zx8iNQYfkTudPNaUjCDbRfvBVDXYaQUMAeb85AuX/Q5CG
VA7n8JVZ42VoPmLsJLtnjV3Xgg5T7kmebosr5H6jpnrA8IoCNzTdTqW4RKnSsQ57
X1lENPpept5cSUO+EBpeftpc34JlWfKhPux2GrE2FtiALEsWKL1RL43AtZzf9rJ2
GbiYoP62yGK7wyEd0vkAvKpn4KqqiSLMikVzZSVCCgQz6EhGeGfMHTny558IFgiw
okO+74r18WUxh39xmQw7aEzgl2t1MwviROaeLNLW5I2GMq2gG8uAo81NGPope8rq
ZdfgYc3gMMh5ooZAL/K6WcnygOCa6YsbPDOSKihbn6UtUjhZRYooCxasb3vfbKio
eq7fS4Egze9NQQllnBeO6oMD8tz6TtCf3vAVR7ZXBAoi0gsSmvebRDLOBb6YKGb7
VS3tdHse62aUQoS82WIagTw4qt5loT4+FKh7TrKa5Ii9K1Znk8c4VNydaiqFOtIm
yvPD7oIXzr3yQGgUyAaTo90tTQKyejjpPMUheaFBlzarsNCB7ATPvGQJbQfCciIA
oMD2oAWXoPtfzWSR+nzCNGTcGZFa7oNCBebrPtceI4DIWQKPVHjrUK/Aoj4/3Sz8
fLbFlhzg6zPLPBqxorbZMxwkjLMPVkwFu4oWxPo1IRpb/lqJfO1rayZmG3WgLo49
1w90hJErlJhqArBPmkwD4uWlJ4y67nLnb9rg1ZbTR6JsotzQjCWt2OZ6Yn6J7jiW
NTuLxj9fi6lnk8WI5rzWcyziuvUy73N3P09Fz0O5RMoGypyruoRJXIb9lPDJ8/pO
V9CZzNB/fnI1CAPYqaJYT0etO4NNmlNqCD8HGpvZHlxlbADba38CfbuB83zLpsOW
7dM6AkClFraPNJgWc0hMlPjtiBVipHgpcC5JSfoAzdjdJH4oWzAQdLdvmc1JwiOg
voCyXZXmbzVEHzHSGQnh4dQpDPaCZLLs+IcKWgrQvDNmfqgtT76dVjg5boZ9xnkw
6txbpXtQmm6QCmaNn0UcnumvSUL60g6dqouML2rXSj9KQXFhBct74u+Czermceob
cnu6A+nC08sWlUON6A0aWmz9/OWmkSO2VhZoA4JNhjgUMdXKBwsdh5HZ20orlYJ/
r945Yhh7QW4tO8zDqVKQorrkdJr7E1SqKLQXnfDQ8evPmrB0r8scUM052oq3i/j+
QyF2FiPWgp3Gto+0FXg4kGNL5p0OFJqsCBkWnXg+RaYaCkJvSQhTkbaJwAYfF1AC
j+SkLt2q4jrKDuu1s1X5z0M4HEei7+48wWECwoYstCQBpcJPD9HuZxQD89ECurN7
rKS1dGw8wKtWFWhz1eRiOtIFhPmDmuQrlvXVJnHZuY+F77Qqh18wrF8m+AdB1OhT
IoTt3yInu5CgP+8f6IfRRYeTVq23DkJnwKwGN0UaUmJ6eUxo9nqX2hJQ5U979TIx
YTPcnLigp4pWixugJSL9IppqMivnN3XvvdktRnKypd/fmQ3vOYsCJPMl6e3BbY1f
UG5UsIu6Yel/6zV31rnDJXIdbAgyBYlzF2085QayaphNsXAikvN5P00qMWmzMfYM
ShQIoXvulhJlGFXyIfEgH50apHzyUeItgUe3y2k9mqvdcvcJqe59n7sG8t2SQwWS
3BGPv18LB6UC3GgzAekPiLlJ5BIARv8Jr9RAjoomVf7CGHOB3caP4ct6lCOJLSVm
gvRU4HTDhixmSEZigBhUkDouiFLXiEBu2hKaWN62xkA0hArAT91qZXBDoAMDMEwz
mXVIAJDWWnt3nIwbNZQJDtqYNJXJjHGzSQ3SQ7IbpMK35j9qJHfRl4klr/6r/eXz
co7GDUXGL9MPi7r3bFBluROwaK7Y/vqpD+UUA6JkFjv5Ec+5ukEZxOBO1IYy7UfH
+KBfvf2jUo2Kb0/CHVfeFk/mEgITN8/uo6GLNKWK4q2nvh86TJfO6XVhxQrCLtRC
MycxABt2xLsr24iDR/SkC7jB+9axbBbi/8PLiy3ykWAf5Bx68PR1B8CXIwzsSgiO
ODEGR+18WxLyqsgeheOqZ82/wReJrgKXmLhO+C1tF+spdhNQk/5I7FnPUlDsEsUp
dRq/jYAB55un0YsBkej7FIKprcksKWUpdijUeJAfvPHJlLxtLj6+Lmy8cRQ/iUuw
NzfoMd6xOysARzzln5s6vQNFi9rAj2z1q6LxPhSsXTfkx+1F9z36NVuWk7sN5cJ0
RyctzJmbksUPnKL+/Q7cfYrwXhb/y0zYzNeYy3SrfYqZvGFoWg0HHMPIzlPw3y3s
8gmT+OoZGBaBWEg7AVxp7u2rEv+EyW7lULTOzywI4dobXLKYYwxGpJHjJzzhxKRU
WlGlxYZ5sBqGEDT7s/13H7qsCFdfHOsZrSEDlnSGDbUKKkNx9XH2sUqotcu7m2eb
nf7ov6sU5T+7qFJRULImhOcyjPkzqbtkq4DbHC3DFTOGINIiBTgdx/gs6Gm3sasz
/JscUpIWNjSyX2oYit8xXeLlABRp12gKe0+mh9wH2T0jhn7LwtOuHX0kKOXNCE+f
gfziO4CxujFVt9lEyZWjOAFVaLRSuTZTjJSRIl4rHzH8eqbyvRmN1ODdOyi1lkP1
VSkaFw6HxUmSoqVWFKjlbw0n8Yecl7wKuMotuatThQjkrYWApR+sKWI5jtZ0wuf1
we1qhYYhmdnWPc1ddW0pCi7vQtqlhyY0SLLu7OgdUj9st6nduLQzr+AQkXMn0woD
xX4UJnlAPSNMnK/4dQbhONIG2Dt/Ji2NBNGzEY5AhFZd14Hew+466Ce1jurYn56r
nqdjK20KbbTnQKeU52kQthQwiAM18OrOYEo2hd+Vkre4Co1OZ0e4geFZkvvi41J1
Gzj64J7o5+3SO4Pf8xnSb4W/pRtAvbnOgvIzgRqQSM/DNOyiJ3NsprdDDS9WblZp
GQdrSw+oOJ5ailxAZu9LU6T5i4LCJ3hwjpfwYrJ7irYniuK1wPlKzC268ZmaJSaB
hg4ol1XZQ9e8ifnN2tl4lwMCGp7IRy4VQdeDjn/I7+hIsTaeDA8FRlaGJbVwo8KW
gIT9/NvClGsnZNBSa61JuQSx1GzRk5enRz4aPad00q59OyLLL2r6wfKgoFm4Q893
iJqniDF+yMNqob5A9NkVvNzhXUN4yJ3oqvv0KSXVPE3nq3qL6HmYG1EKECatPep9
dAf6IRZZXZdrt3/RKW38xc15H2+arIRTfySc5ZSydBLHe7MzRcgqgv2mz/aH1ymk
TbIM8J31xa3RfylsPfctmIvmTQfTHJ20U1uFgn0Ocpn4hfJLh5e+KkU4or1XeXK6
uvpOAld6FpEj8N5UC+mIYozM7EnVRg7VIWx8Ezr4cjzo1KAneYEhvFrfyKH/napq
dpx49UwBan9IBYaK+BFKqPGPq7kjEd22URaRaAaZpUgeYolbJXMyeG1fBpyBI6P+
hgkM7niVlaC80UQotdqUb1be1h5tl+95Hk+TGUUt7IVkX1WBFSQNiVkBrNoaouxB
BmT2985ZslCugt0CG7TEPrI0kFSpgLnNv8Ay9D81UosKpYc19Gq3IjrTHxiXX7gV
JUGdgv5Qlqm88zJqy/F6bS4aNrMrPnNyJfOK+tLu4uUOCeBJyuGwizzBBZC7PWyx
41zFmaq0sB5eZ+4eBfjy4CE/KyevIpnNIMDUC6mD3a2fmpsi8YkevI1QoHjphj79
LQybTysI6nu0ZncPOSauKSSYiUCb1CA2ZTGMfGN/JiqyT6Fy21vLPRt+EHP2eh96
sgkICn8eujGw6w4H8R7ZWRY2qzNi2wdyHT+V/QpqpOafTE8YD7fGJggtN09FpgjA
Nt4bDPSKEG4YDwmZFN9e4Aw+RzC4TsKZZBTlA/cl1A/SN5LJKhEqlmOJsR9gbqcT
zZCVzhZsY8QSofK63/SVX4xodiTLcZr1z6AfApn8HB8exvhYOnfgGoY34LDbqxQ1
5rDyjPxQ3BUWswNZ6CgAGP6382zkCtrloSjPss/mqmnlbTkas9rXtV1hjFHdkUt5
oWoqAi3Llm2wxtQ8tOK/xYiTOjJRSR0UzMsv+/IJRPxj3N/EBpvnFMMJtzBT6ksk
dRckLN6TTr6fl67LMVpxxoIcuVQ1SJx3rNbU0jgl1kx6brcabnVwA1nONpaO5h1Y
/KT+lq8u3C+88psnbXUKEMzeFWMtyfq4GH25JYGpKRAYAe+VxuE6NnczeVntCCmw
ZUa2AdaFoOrpj4VCYKMnuG/u0jMKedV8oEHcr9ZWPTNhAehnutSLGCk8zxtxu84Y
BNB+w5PlyhNDpddDnhEpfRERJdqhHNbEqiSld2cMcopxEfCu5YxY3bpW3WrNhLdV
2VNj60S+cvXwEGKHFnpvnva6Sg9Sv6OCyDpHIPA4dQavYBNHe0GMXRhwep1leiZJ
s6hHTri3/jAIYYvpiJlgvaW7IEhmp9z5BlcYDXglVdxm42Tl7L691OXOHBmEoPCw
JE2pdf6OjKXIRBh5VzQffFAm3kBU8S/i6JDGhBn6ZHSxFxroCXGu1AFByLDKqRfJ
Bwd5kMcdyikbZyG+xGRrgnDfZpBbb400yMDBYerK6+69FtwGUR05f78CRBL9CQEM
O5wWvIaFXVXT7z5HuCkuwPpn/w4JH1rxQ/RpPrUn8YcTwmn5HuL5iCUkg1FB2SRt
Pv9rdvnNljant8BSlZ+HK7znlDd+hzOQ7Qg/8GzIpWneaWDWUqmuLMH3NAcS2QnN
FkQXVpDuCWc4vFXpScPGYFPQKpS9FWzYnzoUOSlnOwGzHaWUgnk0rfc7b7en9Qze
Myw/NONXT/TphpDGisgGUNMzIPKrMR6gPt06Y+tMG3I3H9a+NnlrLs4DYavnbcnH
aw+86UGYDQrVY2lX0PvWAg15NcgKfHHRg1nQ83tT19yGbl8KxEaeKquDmZzLzhVc
oKjQQRlZWyWjy/TNYzCbG7Mk+Bj+MCGVzWPCTAHs5CCfxNv373F6QSYDh89OTTob
IymYheatp6fAMtqdoZu/tRfLY6oVrA2CWjNWj/sL9yii6w+XMp2pf8D9Ox0aCwQX
KuEb+stlMxAMY5KzSMsUAnU8134rO597W9leTU/MjJY5/zzt1b2sC3AwVp9GLZ1r
TW1jUlJvgEppM2vTX122e5hYoCZAzp4pKOoD2NrrjPZ6XBS1BpGHwB3Y85hcgjQe
NK834zpH3mKHe4j/m9Gtrx9xPLHqTGS3CPmZ9vAmlXEc2Y2sDlWMil2Yutm9L3CN
Ib1VIHNjMuOjMal90j2uRvcb1YDZiRhEpUff1pVw5M3PxPJrGoD6YSKwHHU2ugq5
ke4m2ihJ7yqLuOFGJBm1NR57za/LZYmnv0Xto7qxcGVMeAMzAb9sbrqPpD5ldkwJ
5AjVVUbSho3CJmo+ga3/1Hi9bdJje5TwhvNutAdT2c3OQef7+bsMOp5ywBqwW6iL
uAVUajKqYsApzLjSonvn0qUyflXbaWh8Jz2BLlE15JYUzGoQWwkhGrLIxx6uITxu
gsHgA128Z3L0sa8WisZn/dC+lVFEo2yr+Ybrqg5W9hwOzQqGJ3TmxvGTClRlW2e1
R2xo3uv6cl7PIY1/E4wCeFdkSW+zYsekKCBsRJdMKvGJWGEHP4yynqBb6U4deswv
l0CmOJsiwSOhoKcRY6xcpskfLUhCwTnqsU6gUsnoBCPQiupYThD9veKR+Nxpyxlq
7zPqv6avkW5ZIPzCfROvvCKZyxzUNX4cLXKLMumwr2F/69fwKRYOGv28/KDMBAgb
lYjtmJwc4wF5gKODX6U5hSmi3qSxfll3u1LoApA36yUSgjbhy+rdAeiTuCcMXZUV
HBYBKTi0tTkcbGtZ2By0ItH9GV7/cYlJVGAXBNQ0FFmH4lBQ41SQwLfMZhp2+RCU
wNup0pt6KWWt32t133+J5tWgsVRj8TTgDgZpduRnhy6yub1QnO04BEB4FxT9DEwr
/dLMqIchJRxXnkHnXTbL2cSU4JnU07dJTAPZO8dQTsf4k6FRawUh7x72TKxLxd6x
vKpo/YEegQ2ItRRqsiAKyGkRFhgPUuE/RBo9m+b10oraKb+W05JFf0gzcVNUQkhq
UWHxn2eNnq0gdycNmYRbXQyY0QGiGEUPcVFsXNH3PfqyvXk84eA20wUphdBNB/Bk
n4Lj05VCovdMjPUDwfE1zw9qrI1lKPJdEyQ5ABY7NOl1oVTlEri0W/74pVnTvPvY
pjE3YxfGAR+ugem3T6UcPhgvPx/caxPJU+5bsBu9Ggbm/CvM4CrIy2AqLiQrTCU4
fsQj9GQi8uV6MlCUtvasMUmwnQ4PKtLQaZO5nAc7BniDLVf++5IxccEW4Mhj9OrH
UtMQa1CrjGGMYJdYbSXek/Hf9NhCOIYfDaBDUn/KqgDyHUiTLrv+oKanLyefqbQX
FnzCKn0kaYR2Mcglely95tsxAIRK1ABmn56O2jrayntsLN+bMQREQq0Q5qIT2cfK
RiWUjDj1lB1XYtTPS+8SbUR6HO7ZpxsT+Zj7M+NIn9cYNB6lMXXQbDURiuWJqLyj
78JlY8ogY42Gkkj6ESVdubwu2DVACzNBXaDeNUrWw6WrJ2uRAjxF4yzOAE0kI3Ll
ovhH+GkPZJ8W9fYnnCoVfOM8AYIyzxyBxq8QzQ2clzuqrf2hYi5odUeJKw348xwE
846erDZUGKDMcqICIXBu1gx79Rp5NRwNv4gZeC5KJskOYShgkJMizijjA98bL7sV
mksfj97se0i1BqhSBe/G3NdvJ8xT2NSGtrTBEaWHYQtkBwWW2K8d4mhoiyEhcPKa
FDV/pcYG+9G18OYjRLKUggthNJ8hZdb9iCe2cr8WJI44SVRaUKIheqLrQ4styDhO
3ru0SsI/IB+IuFt2k6w2b2bvw6q3kPjkyKkG9jH+42Qnc2hn8Pyy72ga/9b95+9z
bC3h5xsancKg0EYGkV4YyEEZ1gu6VyTJuyW3CHcEZEadYJnPk5kpHUOkWPF2dEWD
0XgyCC5noC3XGTyyHWhGtltEctn4eSXpY1wlJj5zk0+lzI3mFWwnbCEZGBoVKYVz
FmKraxYc7emWsXLijEW1TYfmOzb+jpro6vEt9Q3N0wk5a10pvd9H/Z8Jl7DU0qEx
5tcZTD9ohmEvkfFoz7nb/yXIufRa4maNCOGTJ/xgRtF8Zhuf9dmtASkd9UNqJvzM
GRn2NRE61NWn1dwTtAysMAYKX/DUY2l7hyz37Dr5XHJv0voana9JZV6vKUljsVRc
HisLMyjYvJeayUU/XEzexGSJRsIL09j8lwC6PUUnC4mkxCVHhscF5cFdKKggmiBU
Un/iXFtYrF678egbprRrqkNqKGKzIoeIVCnw0mnCyLBKHDu19XmpuIPiWdWHaBPf
U20CnOADbJHmzcZrUXNWWHKvcf4WVQ7nd8Qme9MrrgLAXpk8490oWTckTwemiCNk
2hUwzqCoVLXkTUig52SQXRAkfQGVsGHYXmBdmqWQR/zweBVbn7aS240VgEoUQ4pj
0IJ+gNRyDwhNKclf3aVrBujITNBIjrtRdEG1Hux/wYrny5AKxPvvA4XsKFBynQuS
9Vtd417hV2S9D0tbyunQ8eY+PJzzchSx7wEKUOm9SBA5CbZI0k+cd5GDLdaVt6P7
gmhNQ6T1yKCJDRCUBMvMMitUPUau8WvgJAWwEvIoADFgqjU2nVe76bmeWtt4/IBC
onja+flaZSGs9T2zUNstx/fDqKzoa0Otl1hC9gqESQu7rKg+2+vbnsNy4dP743CL
oHND/mrZcwnsP/3RGHEdTlvlqvJy3YvcDboVRodVEwGdWS4H3FoUYsq6I4OuLRM8
QG+CLkaIWHsylvqEe8rHEyur+z0MHLKpbQSReuLSatNcOOY7jAyjKRyKSYJrJ2vT
GPlXh9QkBI7WkYUbyV+wvjc/RZKbRqTw5dSB7pNh++kxEXlJxiNpLzjAkiZX7qda
WjklooZls1cHoZHjPBHtzWyOZuS0O2dtW4LZhxcOYcrmgIk/bFZc+j+4NpBhPSA5
nG74z3cvaS8qzUvcSuxSrnr1DjexuznpIVNzGhGxPhIGP6/HlhQoyxEQwQKEbpo1
RBNu/+YS7TiL4iszgpKDoY2uSwVl0ggjfhGwLoAoRfSKtc7zNaXZD95xPhtH/KxF
BJhZ6CRz8ga9K7eZLaZbkn/alp08UqUnAUQq1EPwCYq9keUOEF/OkhSx+FVrXoP8
UlQOf4EZtTXX9FMscPMrmMbj4j6VFyvqwsHg0dfbFjvhS0S3GFd0UEJwOt9zR/4s
JU6nUyYaZU6EIbOd0Lgtd7Ck9XXK6Azv77AI3NeqpF74z+uQv33ExI/tBheLgeGR
2pK2cNab3W7vqwt3Bc0YLzpkS3cGXxBp/PrWHgLKaLzgPsEKrBG52hMYR9IWIC4q
jt5fd+Z0jvnVd93unJgWJOyuLSLIYOiM/baaJwruwGfbO4y60308HloRnz2tYZ/6
xsSWCiSjmsApudOX2Z4Y4TiIT/VgaH48LIoCrdvHf9vK8BOCoF/6dzeegusNC21N
xczXeRmsCa02Zj7q7TB/SoBV0gqwvuLHR8Ll8VZ4gvkzMdKuP8HzV6nkPGFbGVY6
fvd78cBYiFlgjVQw3UfTLzohqVOS41ObIxiJYs6hew/Jki+5Dsiw10hXXaz7/yBK
jhPBkKIA6utyEj8ImWb4cJWnspcQkmmhAd7FIdsLDrfty4b2n6zKcco8U5gokXPB
xw2BKVCRy7UKxJCsvlyzYnGcePvJFJSnbd7ypdQJHMHroEqoOPdyu89mZZTHcT13
6CBozL/SAAfFfN0+lvMZ1eMKeY8rSXXYwBVVC5sje4Fk7TPwxpfkdP19ZQh0dBxh
4b7W6WC2mPDW+L1ipUrYPKtI1vOSqSz6RhSEQhuQrDGRkwdfj2gHOXmht5VcrlRD
Ui6IqWNuoLvg4LV95YOJY6nsqeD+BsOgWmTz1iZO1dKrAAwRKZKyViENlZU6exnu
u632KzePvTjCwu2oRc4Emai4dGXDjsqNk0oGmvBvcWkrIiYqTKfdj4QOCQs38+3l
xD9llQ00fhxV/9XOzfQpMHvmk5DV3m/E77OeaHN+8b7ZIZOnIc0+3OYV5S9cgybl
CJ6a51N0PjmXA88jhTRtxI/sTwK6e6qLC4wcocUdjDtsDp84WpoOHANwt4hWLUGd
mX/sADulG2E6AM+HGZRud+q2Et+TZerTuTc0LCprO4iUycjzqYy14MUSA6KHLjMe
nm14NYXiY4Xu1F8wvZ3zW8nuCcWUlw+mBiQrGndrOU1y83QOOkGVKMWL7NmelhtU
hAh/wQ5MyE0+W0rQuQg2jze/nHsAAnHjIK/KUL27MvYsKp7mGwlcz6esGMZaduyC
x4biS9LlCVV5CQn/QOmuL/vfsec7CGpRdzjzLuf0oRqwL60Iag8MtaeeztgJanQf
A2srGsv+KSneVs37XoJMjF0RgH7uW+PehucpOgeu+/HGcZIJFyImROiBDMvDMHgf
iEQyCxcWAYbX9ZSsy1Dqoq8LAoK5vmWB74DekyggN5EUdR7CoeDhSNAXGoZxpatK
A5f/w7BhNOR6nWTsoGqJUS+W8WIrJP7JXFCQhpvbiVimoLXzCzic1SQjiUuz6TAQ
65vrBeRUNzQXWzXcQKmkfzVQ0uHhPrbwuu6ji0uXLqiCKaEmHF93ovB2uhT+QV5T
8H6TTr7TKoSFt4j0sjAktSIwT385NSuXCoH0DkLElI08hHPPPRVigy8cfefTxJ8p
ND5wEtNw3T6iJkrXEuPqCFIm53ElZoKM6tdt2DQG8LkZqCiWOAFs8V4WQFepC0mx
LT7ZZVOSLQjMhud5ODWge9plyfboVzBfczLCskv9Yohy4SHmUKviApZcBO/9kjM6
49MBPo6ZJWnS5+D5HI+damMlx+PclNsPBWlIKiAWQzoo7ICkr7RjA/Hr1zpCpjgL
my13NVn+1MJF7RsC7Q1zHKDkOXb/SPwtnkFQaZ4C4AVj96+3k+KsJjfaBLp3kzhd
oXqOnEImmyrtTZgWByyOkY4T1CUKE7qj3qtGWryDN4rfjAHMoN+S27TigyXoy5eu
LTzd2YhLAWYimkWd2+dYSX8ksQQaBkb+oeMq925LALcbFDmqnn4sJ8DWAWjJoWV2
0a5/kttzPyge0lZO1js4psjTMhMVvRAzrz83DOC4nOy0d4cXSK/BY4xbeVkan9kN
pkkWJmd+WrSe+FSOgXVEeZTPnfQs9zlTpSrDF2SylLQDJSd5ENVV8ve1x7pujCiW
bqM0Gp4c1QHEYUaIqrt+TeI+OVk+MZipq7KM6Fj0+6Zy+BAc6Lm4L+ceUq9u5n1w
7kNFTpnhFttkK1m+6hasI30udyZsqUl94T4WBg2AUL7yvvTIcsjjDsteBiC5lpQT
NZg4nAGRKN7sIZJkh7+xLqAnpyYnPZIdWm+FdfCQ8pEmp4HfdadZvAmEI7DZtK/6
pTInqV56+K/7NDoVKclDc6vewoFPrIEahWbgLjElrz9A1YAoLiDqJ6FhgbSYUYfA
l8P0o/RRlRpPaMXp7AT7ewr9zH7Y07KIsE/sqFfo4gAHsjjp5/mc7Vu7pjds7F4N
UTNF/mbXUhsKIYQnsg8OsgQ8smyVJB2HweNOyiC9bM78/N2AqeGzQxZsP0KjmlvD
S7Jvz1xUCBdKSKe1nmNhHA6KrYsPDT69EXe/T7HFwbmV5dXBVuUgUQNEgwl2RcE4
si8Gqbgi/RTBhE4cOeCtTxZ3U++JKhs/qk1Dpkh0fYNYJKHvPFK5po7rLFijaAuh
nMX/UGsrWNyEwW4ar6gY+EF8fZsARJpW8bdp1w7eNntIi+DeSovH6QN06yuaedh7
cNq/pUC8BWaEk0z5x1LrrxQkw91/S6XLyrCOkm2DzPe9PQS5NOs27Bq0uCCMJ93Y
C0D/yur/1mxl5a1irFy2NNx8Z74wF5RjV6KQv2ueXZpmqBtMnrTQmDriFzD9td6E
B7R2l6XEUKk2BjNTz5Z9j+0WCcKC7hZFIN/kaDAM1o2yIIJJwdk+AoZTMuEujc7Z
MqWp0oO9pBoKUfGLXNMcTx0SHrsawBCcSyfpRznFtdsGFHNoqE7pbL8NWXLfA3fY
IcSkmYGWSpUmIFbs3/aZ8aFn2io2+AgvVb3aN9uZWwHS++wlguGLUGQea3NInPbR
9srcS2dkmd+ZsQXKNcxXC2K2Uz9sXBN988Wd9/Bn8KXYHoLnbSx6qD7sD43SMUTb
6D0ZR6YBXRPWraUGr8vSBQDh2sk0KEXuYVL01D+JA/6qLOdilnnaN7dfkD8YaIHR
0N/pdg1ZOWjH5b4n9xarSkaL9If+URTl5UhYPQCtmB5YmleeRtCU0VTDv/3R6CpV
3I8ff1BHT4wFhCDSR+Hfvo5QHLtnhCh46kbQUhtklIE7rUn6p6ln2ojUc/X83kM0
rqGJn5xOm1go+AQBd3ijW5mmxWm421uJEcQ/V9Jrsgm8T537azrDwvbycEPGiVYS
bUAB+DK7jL7j+Cs5IdWxIlwpvZQbtss5cu1qzccNMyAtClkl4k1Kpc2mIhGGM3Ti
kdjkpTXEie1SNGXcOOkzc7znScf5EkgSiT/6m86bHL+YtzZo5yS3Xt4X9ytncllp
932DeZ1NBRHAXvPh6i5pG0q/ASr1b/ZXodKj2xLy/CgDgQ/bCHbeJ10XM2up/UFT
uulmPjPqmBmXZ2ii5pQd6XTWK3FLF4WaeSuzvAe/xd0RduJG4mv8Nmsalm5rgqtf
33IyILHYFqzCZdMr4QP4rWWr/15Dm05EZCdaqLwNwXsD2cv5Q6+4dsREgEWBmKjK
geiok77mQ1GjU9/ubHQb9tl44nDEkWJjTO2jaoxtMb0MbESWZCO9AQzCyQ68Uv8v
GvBuLKpRHWz98rJnHTdwvE2g2nxa08JYnOluvGTPqgmwWQnibINn6tuH62JLEmC7
rnvIRoCjIaNMs3fcb3CZu+OEPAg/2nmHCIJtDiAu4wv7Gdy/5cHVaX/3MyHRlz2M
u9PRXRyyeDstVm5dP6ChFTowZrSDGM9RspawHnUGFBzPLtw9kyXCFRqSRoLD5UqC
Rp1KQNxx0TeZq0E5nUdUn9HyGnYJWgTwCA3he4jvR7RcSKIbg/JOsjHcQeqU7718
1noiLBI9E+SN0JonRb/BBs+kox2f/YX1mrAkgmVPEh+9iCP+5Ybkr/FUkoxoAzEW
XWYUpNdCymDmv0OkNUhXQPL6evgdPcoeGyukc4FKgXqivX9CbFVMCiAe+Lopss4z
JtjlZ9h/lZD3yY6ChjhyGBWmzMxvznKm4W3v9ssuTjnOuDF2g7F0/2hE5L6dtizS
US9LXHvXNRb3trKIaFSzLeHDRKadcGv0fZteL/a5BgfDGHydJKmktazBQeaBM4uc
o1HsKIQv7/EhjtQXiV771yFUl/6MPUGK2wi9mdhwxVKGai98XkfGLpe5h6IyrPAL
FyApSXbLfhFPJZoxkHUj5W/+QR7y9ApF0vdmi9eTMLYIB58P0JAfDg2CShZsFggd
2au/k+jxRaF2/GkpMxTXYVHNP7F0XOPt5g7BNSds5QELvAxM5wv0nkLb64HuZB00
GefXwPpD/rZDUscmkqtu6k4+hZiwH49QXB5D7p9wed/ro8QpZPlAyYZrYXP7J0Y9
+eZzrlWM9QUDhXLqqeID/8U6M4h1wPBHmbJ4Z4Uwt5sLvXrBZU/Ab+79Ln2tKTTd
H87vnHswmeNXW4dyazg0VCt+7tj//NV+s38pTpATNgSalj3047OhxM9ETDUmdioM
0U8ho6bx4XNgaKQ2B6T+Uozu/ZfQj129mL0fVqrajsGD5fDY9yuZl43fy3gy/FWj
1OC+bl8WH/iyFUYGEJYLrpooCF0Bbn5OzR14V7tSMpLwzIJLmWmPDLqJWj7IqEF5
8Iy8YaRtc14XfirGptHtn66y5idTlz2ihWwhodn5dQ7gFSHErcz0s9DSJNjwcaJX
dDw6Ch3XhyI9Vx/OdGmin5griocc+erhbQ8kIklKucvoCAY5XrVQzbYMuIQWvA/3
8VFHT2sHYsM+dOV3zK7dWBwwLsbLLYjdvO80e26a3GJsnd6IcYj9f9AUcyfJxTsT
tEyK0W6cNYgKMnVnNwhJaAmJgvHT0hM1I9tmm4ZxFn6r6NTZQlLYS8QMYmR+gewg
CeUIf1d9WiVxqvvyaiNxchab5/g8Vmt9dt5rShI6X53P2cXmCSCviX6uSUeAby43
LbvCmHsk59h/6hw3DrJVZs+gNqXQFHZNb01HghSjLlUa10yFHYM7DYjg6VFNYbZ3
chhASEfsGtLlVq5H9mZ3ORDK61LtIWwmE/e04INTUosJGmLjdLTWYSbOFYhHftJh
NjGOe8GmAoaKQj0tbaybdnJ64xTpdGHRl2k3a2GORR/kMWZ/7zEjIBAeWEhWYzkC
q7bJMQeTyEC2Yc/x/YN5uAm8X/4lW/8NJrRnJfx/kwmbdn4rByBbyS2Q0gv/vYYc
AgnYAUJjOp47b4lucwqRZR3jWtEph5bq9MAoebrXZhAYo2noWM1LEkLr+ps/u5aX
8BuYFQvqfu37CpuE2bS2eLz1QqJisxss+u1AEbeGl40gzgYtHz96UvlZhqRhg156
jMSebspgSBSoPIv9flWH2wE7lInr984q4w1Gu9rJbW7eCjWIimaaNcu0QCccdPH2
UmXs+R7L8NXLePxwkKKJ0O+41Ly4XAEJHoT8YTs4l/hvsSUOBStzOS5ZcYmVrXWc
ERGythrAvg50vb2Zui5eF2y1UXLaAlepHZYfaz9AHLslvyXOpQo66PAvtljys5Ra
9a15bEK86wYbe/Dwya7mYtSTVEaRTm0CS0hTL/Xon/rIO9BoNC482NNtFhaHNnhk
ULXyB4HQt6bT5+WUoD6p8zKCtSHpU4964bbck381POv05nl/x9AUBWTFZZfuSOJO
68e3xZ6lVXC60uGtp5IsQMBkkPRTVeGgCVELUTYN0gkGHsRT91Mkm+/sfAVlKuKa
4ODVCUHgvI8Zf3F+sfGIEqkgSh+9bH2ggYO2h5LF8yjJJb+gSaybL5FwdCC3N0oM
WchOwvzt5A8BDtb/jIyVEn26YvBYHyoQikhWQ+vfKQF5ufspka15SxRAQOOheEEO
jahWA65c1UFqKimKBdgF+dr/Ckkfydcfn3gGQPQg6FhTzTJSjh4inLIo1gEJtQkU
Rwk0GoveZqZ03gY17G5I09h7nXQHMEJDdaWtmf1VhbPxHVRnBbeBmVgYbHTFT/ma
c300CeFnf9zL3Xo43U4kpewFaccJbeMIqQ85LvL0cNjuKkEbJ4vlIY1L5bLy+nby
OcnK2UvcxCS8AtxmdnO8n+avCRO3IoIJi5e3bhXXe1lG/2CPiut78ZGIgRNIncdL
+SdvZDJi3ao0qeN2DAY+GjDBcd4qn8Vwy7W7keSM0Bu3R8bm68u17SABRPVe223x
Oxy/Se6Eod37LRmswMxYN6SS0r2fgsvto2bg5LvLdnUktY2Png8nkEIrn+9azGft
DeJ4pSYUxfd+xKrra2ER7uD8u9yUt/TIsQo87SUl942cTyzn9rNCepbULGlrxXL7
VOPC+uJUQxoPhohj0RlxTcU9pvfy1XTq0dTr007K26Ya6Wzf4snqWRxWS491iIkK
YQ73Uxp2hGeNsF3AkXwGPcBFzXYvi6Ya1zXVDtFX90akEAnDLtwHYdCRMJwf7Jd1
+fFvR3DnIp5Duent3QrVj6q50QHGoztAu//wUnnhMJ0GkpYXGXZMdOQWn+Itx27O
hTUIMSUqjVic+tUALXwvDUyJDUITHeeNWl2Gt1kqMTMhRSxh3PkkcuIBKU+fWt8k
s4yEAM0YkWOWsJkSPadPVovwwr+qFHLjNegQKL6V3k+5AOT3NZJcBMIO2dWClw/L
QwEEUT64rQmYy/rnc1l3fgAS6UMVJfnpCTqM+SkblrPzGxeSxni0iKfunOebRm+S
PR3N8hEAoHZf28Nd7KSL8zDYQTOom4QAcEwsd8poNEkb9iuPgbZ04oBGvJxTGvn9
7e5ygE/tEkDiwizzvpKwF1NQk2quYBGk1CegWhCCBCvF5QG6iRVXku9F5578wzd9
DORGFjfSiR+a7TCY6BLbCd99zgMjcmuhRogGCOnKMRCzikQj7joNhhN8/+KZdE4V
gnTql6Lxkvll9b+J/YbTJO+X/GDEmH7yGbQzGfOkTgRpeWnADiQVcx7J/ZRSHpP1
tfedT38Ifz8Qm/IgaAN+DQGgGrt5WSAAMLRIg9bZinVpZBn01pktXg/6Q6Km5NgB
QDNLT9+uraLsZBLVg4TqpVkFSr4TU1EDGOuIZrlj36DbqYAKMhMu3jVzT/Ec8aWx
erIQ+oMT3Euf+7Flf3XnG0r0cdUWM4vfqFFwyAicsM0ReNyJawt1gGtmjmxw8wP6
z3W5UOui+6SLsaFEDRGRpLKCpKBP2RiD6K+zRHiCfgDIHGXAcp9FSinA/d3jFrHR
89UP5lc/O1qeyDmk4dyzCqlFdVQz+kULqegSAITFvnU5QbpriK2qg6dD1PQvdJy5
Jze9m3rdFU8xnRs5cAfAXTgunDI4GD7og2yTUclqmK1nbzxbAgoDzibFymZ7/4Wz
lvci4FXLWHNpyz+6snkQHvblEeiK5EeNTFMTruFkzYio6MDIn1zJn+pqVc7Xtjmx
85FodieKMQVor/CPToSC8qUkOag3Adcr0ZUAZLxdVNGthHgVgFaDUe4DlKD8Aq1X
K+UkVmtd1R5ocIVaKHgs1wATGhsgNi81vy171QUtjpbXb/brVcLuOtzAkQlVgHAJ
YSLO0kvNv1qQIQA/j8uel/eNUfaC8ZgQ+LFynIMrlkfTp99cB6yHgHmPl+MNbP7A
N5itr4MJfr8jEjX43ptOMhF7yXPbNoODTsrxaG3BNJre0ewcHMLG0WoLnmiIc5HX
ueMK5OtuoLvDCJpi+EuNZCJqk+gCk9Hk1qFbFXaconwhVo8271nOZ5Jioz0rxczg
QXgA8/RZyHxdELcEd77H2TFV++Th7mX03IBbolKwdASFp/hs4MgVFemFElJAY5M6
T7sb5tIqeQjtrX4jxcq0BixJhxNdeXhahXAG2kbaPHnntYgfPyrcryWqe7cFtOtu
Ad6zBRCYdxFY+TInw0wK76CkLXDx0QxrIDAws8N4kwE2SINvAaY4D3Iof7c4oMtA
WO4XSqRJs92zcHr80Ph+Ow77wfGBXnT1CXB/JObzoRqdyO/HzVh7KXH++/hibWXE
3w5DeiR3JWOm9Gu5JBBzt2kwUsekwmpKmgmZVYqh4zKnz/FXjfdpPjQzUPmKkWI6
Gs+G8M9Q8gWC30vcdT+I3U7llsmWuHO21HM3UO0dVS60uyk6npxqYZtrh7eMAVPe
9LBT+CFGJhjjUWmMRfxqH04HqRqJDDRJmZE7pT1vryEDBLn4Y5FxQM9O2G4M1IAz
XIBYZB9KaahbhzNxUOBKKpQofSFqozlmgCk85XzO0qcMueAAhreo7fMPAJCJiyOf
1W1QQCPWzCA7k6qJigzvg/UbO+SzMrsmBOrKH6RlG38rHIuI1BwR2praAbItSWLf
OI2dCpqpqsU0K5jxeLxXCDmhw9hT6nIUQH5NpA1eAZu2hD5xq1a8wX5OXFHAmuGR
oPSp0t3ysOLPa450J8rJg2LOXc2/7ztHrLaRy63seX1imEMaPeonhCYBepeXyR52
pengPwLZ+gtUX3bu8Gowoir33mLWKgL/cuNaCFlqFVjpoElSceih6MrgM1/+Vzo6
F1M8ecWMs308q0KrY2HSjFxRjL7D1eC0n5TfEpS//NGECYGf5CXBHYnyTk+4AMQD
LZRdm9JmRLoog+i0o2m4bWblbdP63kkaqpIhpvjFNZ2i2T4zzbmvZYbsy291pWSH
vrnsMyeLGazr1ZuYF39KaKgg9GDq4ET/LE1t4gEPtqSU3w16nDrDu/rrFY2pdK3o
tLeAu1EbnVrs1VNI6MvQPA5IvbX4lm7hx0BUzz+FqeaPGQrdiPcpysan0iAEnivJ
6TwoX+15JfC8M+lOFi338ETiKzD3FhNfCZ15EDD9JaggNNBL6dSe12lJwo1KF7hG
mE+DHoyrfAwmHklQ/ly1iwoZm0dvJKiWTKv2zQi+lJBgmM8srwlsCXhsP1pCYczj
0AXA0kviI462qIxSwA7cIJ4cWfhaBodySvBeD21ehsYjlBSUnAwgHqgGkdA+cd5Z
WCdy4RpPZKRFv0SyHRBlMtOIbZaT5qUCvwoUcfVQP0YQ2Ek2AhviJ81hFlOCtgSZ
zunpkZUv/Ve/STNwEk1Z/dgCk80a79LBNO+pFIpNZt7PmZEINonR4uK7r3jKSi9Y
1a4Uo8xE391GcvtKr55trJqMYXBoaev0LyshhbwQE95DuO2Z6gHE/PWMOcXgl75L
amVGMdm00AHIMnrTEgA4yIcJ3m3qjjqFGYRbGTZbHmYgwkyEs93/3wPH6KqZCmLg
NLyU2+943nrFC9n7ZhVSerVva9Js3jl8KvgqckIvjhR7iELxHEYpy9o6XPFI2dWO
xHeQRyZ1lBsuVHeGZAjHqVXNjyubnFNxk5oumJJj7yAhMiEbc/9HaWmUfaZgP5aF
LvShK+ahEtckdOGqASNqJ1CxCfh2y1apW3lTMfAfxYmtKQlX0qDeaEyXveUaPHZI
+4FsS8ByIrI9TAVoQqEG8AwXaHRJxIAklxTnb+8TGXAVpGLp5VfZ/tFmYZIBgG6x
x6l4t+LcdVBmfDHCajSN9O3PLf9cgbrSFgMC34P+RzlqQw2KTK8EldJHVWNtaSeO
VK50wXLXoIWcETSUg/xlE3r/trw2tPfUzKHXI+w8QhmE4Fk670oOf5AZVMyQQm+j
MEJpS9SUuuBHz35h7iGng1vOEaP2nuZXe1Zqs7ylUBy/HWCxAvTom6wGhJOcKAr8
3Y+kStFjsOYHS4SV4kohYowz2uh+rhOBjB1tVA9fAWf0P4NpUfqwAa5IkUB9uMD8
gJoymLfdjCNdPTSz3qFKRBktddhOznds9rAPV+icRwjavCeCVUidAj1D80q49+/7
ozfZkgmsxAPQqALy2wvF9QrwkU0tqiFlANhgF/dqBph2Vg6CUVHVg61OXowzluNx
n802GGqOhK9lLgkujo8+HPkIMDukofkp33DSwLfQpq7r576CFsxACrkPmtV0TTy6
/y6Gbw8GyVuUcQMRQtfJDT20zDcwmXmB4aQpC8NwTgNl9GybvaX77UrXFX5OGmkL
LTfWO9KaQdLZ1fzWXoau+TgD4xlO6SUFhwDaeGL043Kts0f6MXnoJtSREV3z6Du8
pJbzl4teLmCQgZQgIM7sLmsxlYHO3h+hZJNTLPOqIFZ3zeM2u/mxpYi7kC43e+xr
hkyU6x3+3AcjtE7nRHwAQZ2BCSj6fFarn2HUoC+5Aq7UbniaQ97NS6Npz7Tc7FKX
89367bG8gaCvTrx85tJBHtEAvTiZ6uiDFw9Uk01pV7YvNYqpiFiz3fWnydfiO6B9
qVdpZ8CZXmv9+4Kk5F3Qp3S/Z9MW/hWBoAyvZ1SOycT7+O8ka9TnB/ZhvXzdx/2X
2PNcvilAYnBVpYbOERrJA5pnWJlqrxnB0xkrLTcTWJ9wdT7Qfi+smp1MKv4KQvwG
PGyVHFyGZ1YfEKoeEF2tQl5qT6VU9EjM2rOvBIMEDBa44R+zid+FyWhhNG6i7YyW
nooCUdNWn0ffOFp/qGBtw+Q3wfagZGJN32akhmUHPYw+gHZQm+oyXaxJj27/dLev
mYAhoUwBp1QghBAFCaGUhJqi72OfoKbKpiHKiIYKqjM0b2Nuz7ceOxaqTHuSzqS0
ero014y7141KJ7oYQ4n0VDmJuZ9yuxuvfKFJ0hrqkNpP3FvxA1cVFydf97g6+ZMQ
EcG3IQ8lbNG93jgDPU2V82XZMmQ1rGJSDqtotmBo/2/5P04y6qgjPubPkdj9JXN4
sevpxs7wgPr9A+AKWafypAAEROvL3nZ5IFkEGK0D6VJJIKqZXEe81gXa2KnyjXup
K/l33ol67qrblaYrEVXYQPK+7ugHWeLzVBe6Cbk6Rqsh31X1BLtZEPMu1tWqDuI4
4J2Wj/Z/qwSuG6FCzljtWFqnGlyLDpbnBVmquv3AWuEkOwjRFtyJRGkwMivFCLMC
Fpueh3JUfwk9tOVLk6ZUfaBKBYe6acEuEOG1KTPmSLjAIdvVMaZ5uoJ4Z8iGIYH/
+ZeAUgo5Kgti6HP6LIMqwftjxv2I6StRewTgHqfbt7xivQtMRErTk+i5R+gXx6dd
VOnhXxExx8N0RCL4nM3mbPyG0O9GbZhMJd7orFRI2LJvYQvCWBwnx+62T4/dOMbO
TEmN7sHZuGOjYpkPWBMnGheqHY+Gr8zlOkKYdNS3Bat5Sp8Irqhn6p9/CDdYTF8p
rIIEmSRKNOox7apZMJ9y4KuiJ8J1QhyTsAyXSQ3dnUch4JosU/J8E2XK2R1iJfKP
MXftEPn+kwDZEcDjYjedNiOCV9nU9AZ3Gf4hcYxrR7SSRWUyr02JUEWZXt/QU1EU
9eULevjuLFI/u5ROhC6w3SfJ2zhx9xzXMLcUDZn4s7oMch5P+iahqft3zvT6ZHre
XcA6CVmirs+4MIVhc3ZgKnP+zCIB/20szGRA6Gr9qSjGrEqY6UAbQkJF7OAMXbKK
Q+pQ+2x4UBheR9qdu+rPHPx/eojUoiTsIQQz/6rPGqMZD19eni4/SL7CgdP4Xxqf
KzThFd2s5aH3EWSw7zPypPTFZ4R2zUlnoQT2g/R3pk4hbcV9XjJiOvKyaE12S/n+
M4+ZhU9A5XiT5xqCEJkTZT+VdOPsJQNsSXM+eSnBIlQTSkzBaL1QoM6XPtz5A8yT
ZzxhDWgaknE4aPJqniGfbOD5gCdlvaB4EEKka5XO2a6OK1zdtJRxANz3kprIdEQt
YTiUHuKmZ5pyGX67jOZQhu4PabdSMyHK1bSEj7Pse/haRWc9oM5b7JhtTAY5/QqY
UzlYUgfZ/YKQIrsA1edzBOu4FzblJ0sD70QjXb6mn0+cIXxPLCJqSc90cz9uhese
WteEZQNT/SsuyG0dFyPOF5sG3ThcgdhVlaoDgTkuhK5zOOKRDGXTbOGXw34cwwp/
kn3ybehE10/+TWTHN9gDeWqHegQ9IyQuebxiauB7E92/1Z/WgYHE061xo0vrStL/
mI6U8fLJhyKEj3f73PzkDJUxv3LxuHTduB6vfLhL1Ylo0UGQB8y4l6RHgDa66S2q
LCzQV/2LQWkz7Qs4JxHvc66LbaLnQXBi8ePucPwK9P+Zv5lkzV3iHQninHXt2Ivk
VvMJMDvv2N82ypzn3jLhmlUo5zy/38LI3uceyMWEvzsy6kBprZZCsN4IdmFNswNG
A3zACwxgNj4IvAe09GN86PCTa2nYk6VsU7w3O5iXGAnR76/j5cpMf0TFIfm2j/uO
6FyRkVn/1Thc3QIG80coaU1d6IpPM00Vg7svtEA0XKdVnvQK27DeG1iNIt+8GifL
nCBlaVNZYqJ24UajQhPWeLpxsRgGMErms/W4MYVKy5RfNwCLe30rxUiofw9E2Wpr
G3UCLMWY1zuv4fjh4NCf7lh0EFp/sF0tvWwUCKqB9ggBbCwlz0lYW4A9W0io2+Kl
9xzv+I/tKZZHqPSRvZnYgneju0nLJkEIuMlp+kN288HL6FlbaMpKP08qcE9XWdeO
kbrlOzaPUZkv9TTxGJtfaNkmvHEbWX3enfreRwlEzQ1BHTaUxwxUBRZ5y25Umfua
u/mvsIqHqri7f/y1JL8XbUzI7ISIcM0qZSKF3qagdFgmFXvIMqvXSra7ZspW6G6D
12H5Fk7Jxv1mSXVvmwtsbC5HBZmFGON23VJQJQcC5eZayLWRYuPPvsIdtcoFq59j
5ZyuOS8ELeuSaxk4b0drJZD0JQorc1bgJBDp1smPx/2zG7rzUyZlW99GhLwhxpCd
4lQB8yW3GEoOo+yURdALSJmTcRvpi6PV8GwBn58NPoRu9G0f6Ygno5QCgYEt+maB
9xMg6cV9VJkiBHXexdGY5XEZsiLTJOyKTV0KJwBSP6jeXrMBo8mc2pLjUXjyFlmA
yNcsQGmgQ53OU/YBOdK1Vv3+caYpjUYDvcnPEODHb421/iCFzTRlWoVpFM8s8kkl
FsPCLuLFnJpgRU7wmYWX/KMjT/HCUoAIJ0xdKVs3d6ZsbLrhs9xwKrqXI9BHITWC
8yAp7puM5bTW8BjnabDpFBHv4T+56Jv0VxN3AymSFwr7qm599L9BLmmwjtd/aRF+
GTLZS4XIYhQuA7+6rENto5kGwZIeZ5RU1PFaDerd8ygWv9/fNf35L1dqG4dEKNf3
33nSemWKd2gCaeVtlbxukytVJgW1PN9RC0QEjoWHUVn/NSj68WnDolQ/2R5JWwOv
H/BKd2p/klbVO/Fnt+OXK+5qJs4wbpoLBUmcLuYmdjg3Jq8ew2uIgVGC+1oaNpGq
3XHR/HexZrcl0w0CABmJ8SYSM/4Gr7iWxB7ihfhfi48yw0ITvDtErIb+5E+K8W1I
JLbg0Heg9uvpi8TbdRVvDJgkQfAebYpkXnyC5c6nG5F9Hqs8RzeMZb5Qb1Rz0Zyc
Im0p3dEq8622/iMwglWUzawL7Ztp0YpTxlYChNMXf2qV/V+Jgxl0RRNga8RCaqC2
OC7ESbyaeOGuosCoQ8m7u6MJarLQRGeh1oI95qr4B8U/I3cM9XW+KVV5o2vxweYU
/XSFkGK+qFmZfbLNZ8WBJoPmekQEzaP4OmGBlnv8+BNn9tT9oJ6xmI/umY1yXeQu
Rqw+2vJ2KFkatxbWINn3ORG/liEf8AFN8WZ+5C8ZvdmfE/fDfNMTG9Ia3RyyVbCz
Va8E7WVENgIcqvdyhpPS3Qqs+6nQyO64ebthlixaiPs7Wo4CZLuHLQg8L4adngOl
rn/pI2dK9P5iAigsXOzDfOTAlUywSEJCuY8gkhCXSgV4zy1hyqzyTlG3Z0Hl33BU
mHs7pFY3mIECVguf31rDGxrF9/z0lGFuIApEEMuIMR6B2cN/43NpJ96kB2XYncJY
AIHBeXfIfSN0mgcQ1vhAxwpdT59OHR0S/rLsxbS2FjgUBf4jZC4NS3E9w1XM682D
xU2nfDyzof5YlByIc0onwZA6ePHvYEclKgMDkYyrWmLA9hsQnAQ4AV15suPLDBoT
n43w/8lDRhzWilA12xHKVHcgMGcS6lp9/Em+wg5MH65+5VpsS2h1pkcOEVgxEi38
qroBNYfq4mbQ1bx7tagA5ISFfRiFeNV7SEbx9so5H4Djldvl1i7ajHjVsRruwqZn
trEoC9nxiCtfArJkpR7l9m4pCcQQSD+hrfs1G3qFzex8B1BgklZUrzIoNCuzKTMY
PpIWPohcMyhlw17eEFvnIuotuEWUN0iglm/Tycz6Ef+heD0JgdTarc1De/9EZgOS
DFhTbLcYEEw0hEjQZdXuUd+CNfIe3aPBFuD8rYlD58djdEo/tELh7yqJYS50tabU
ncS3BMAFOVRm6mg5zvYNMJLGrIMy3pNZgWPdsGEd/zxzgxQUX9DWgd+l0jcQbBPv
fSAUMQO+CxyNbCopyNNE59CqMcsPuFbVmqfEI2PYQ678FxzLHTp/4nZeti2YWGHA
w02ziFJPDp726oDEw7YgvAW258VBHG6xQUVES41PYKBEM0AVVgi3dCf1AWxUa3Jd
1LuPKoop0yh0qpDKSF3uGJ8WOAyGXiIbZF6Y4qv+im2F7TowrFIB+7cYz4V5sqwd
bniHOBd047fbVf+alvSIusp511CjDnpGJz98y66NSWdwlMmZTu6puqKaz7YUO582
MuMt/86NmfeTvZ/zvUc6HlfSgpn4qkS0u2T+7ZwJRMGCAV2zWneVOS3zSQYsmaiO
ycU+OZ5C2FD+ro2COBCC7UadE2UcrzfRPLuwssl4wCJEv9S3hd3Ysr7ipvoKehQC
X3IcqWma5sLyxkrLk7ehuY0qJd522r/+94YPXfmc6nwKJavTYBbr/ROAipW0DplY
s9jlt7B0IAfXQXxTK1A4ZtGi8SxO4lSUqIW/h6JfFD1EPc3TNyLgOVyC6++rxFJz
IOyHouvi2Gdyj0sL60U1poVue3969PtyCRbYNIJJyiIZa8zWbj33Pu2y0zY4sWiw
yzlkGVPWKyakSuqP1BJhhUiyS2VxfCiNq5va14YEr6TplPPIGR07laDkwbsTe7t3
eu/c3PMQcSI7j5gJc31CKMbCvwf2pJG23f5clzawL82XQvEnQ9rLt05fU+3qxVT0
TIQdfmXNMhcMWv1WUXE0JJsiCojvZKoJ0jh4wATG6ky4oR5VO7AWIi7/SHyd2TYl
IUaR/CP4k3cX/sPOxCxG7dXPvWJHZ+O5K/WO9M6Zr8kPnjxYnK6A8y43fHRP/B4D
ElN9Wtnkos5c67cdcZ+zUUAI2iJwEcgtwB790l0Kn7KZCRvjKBjzghQdA7BNKl4B
mhMu/jmhBRsffkBQ2stNn3y1OT2ZcCBOpYRSw73Jgdb3+0M7U0TMQNJYP1ZsDVDi
pvFoyljh1sqv4ONSQK4TNiKjLIftZM5xFYzdmodHxxbGgLptO0Ap+rn1cgRtPht1
Riom8/hq6DBS/PnvdEkGy5nSsgyRWyeI3SbwJI4nHC7nQmknuEHRMq7QvFo6Qzwx
YOdfuDkAgHxXM0QpEtMJgb8UZO/XwGveyJgsBfy0jHsCmtO9MtCsnUU0jjYxaL14
SlQbTTANXldkWQOVu3J5fbHtDkTIU8hjrtG8CF44ZIyae7hWQErVtJqgiZ/MWcxF
x0yDTP89OAfIyK9jSCl8IrD835Rgmr94SIbDmNUrSN5bN/Juo6t4bi7VqBM0yhUF
ir3LvXj1vPmKO6kYfFcmSGjT0CnhumlSBglk39xFUuyEjmf/oxtGSF+kf/BRDGZ2
+8atV6RtXm8NA8xUPM0A4HfzAeXHlYXzL0I6SrCPR3S3fFVPDewguewEbGypfO+r
MhZsybjSgqMmnFWlo9lTpOi/KCuxRmaX1A5dB+4cV+lihUw42jzC6GQrxuM8/kBk
A8EETV5CwYoHcSMH7/Y71uocmDYa9qv33sTod1Iu8EknnOgguKFTlZSMj7D2vfpW
8iSMMSkBjH3TijPPtY1uPpitr5r9/64yTo/zH/hEOdxV4AhwYgDmHwKdBUPmbDhd
Zxu+EOClu0e5vj5sTvD+77cKmxgZiUQeVgfC68J5bHfeMY6SQVCkUFKz1auTLgRu
qKyiLj6mYWvNz3m2aZm/OWSlUFtxz2hy0jpuqiOIHSQYU2BlB759Pa1EDilphBS3
rCVnGHQODNNUkr7gNYMz4HR7bmZucOfjS1sURE3E6LyFEgUQCk+tKOv3J14Dp5+L
w0rCzjpbMB2hLOEuQwY2q3qGDRLLTNPNdmAOM1W+5OipTLJ4YlAtZRF/VD+O1pMI
d0hhQn3pLTV03v8dissQN3/vf8A69IzvZYPRs2GOrIV7I+LpZzb1lDAtGJxCIADi
AYHowpfmmMGQ5yROGLXfK97Q8R0YK5sqALmAN7cvq6bPZpBDysYZ1Wauu/qA1LZN
kHECmvCxkHQR+apbmjTNzO2ftQfP8iTlr5NBnyO/kw8lPRrXBrLKX2jopmYBjr2n
xBYilvvVKnCtugSia/u599NLJET9KFbJPRuDYPphJl5dqW+1UzWH1lklXSWbVMD5
oimBkCLSZ18LGNWJ+7nLWHR2/iaupNGbuAzJ2R6tYJmd0Y/+PHMLj4+meZpOQz5r
rafmp6KkjTjXQ2u7691VqxL5JNvpewubC5UxS88aijPgZ+Zavk13yju+VQ33Bui6
6oDcvMuPMKgsFeCqHeQ6QKCKJnboBKcl1rQgLJEi9DQDY81wflFcYO+pm/6zLphI
pVSeaENas+EMwO703egAZMS80Lez0cub8eyNtd6TtEjt72KrDclOhIUUkPn3/eoD
DkkfwxQZcvtkEmpmDRoSnwEzzkaQjfCPvcJj6jl0lN4gy/6xOVXTvhuQy3RmMx2+
ZJQCIRtsV/HmyA0k5KT5rXKaK4bcAnljnCqeI2QHw3/yTHN4vUmDGuvcI9+IbVsS
1GDnry/jWTQpwZOsXFXkuOn4j+Igu4zp612rFzuhxHjy0CzdPHyYK8/UMCWMjZ8W
sJWDfY6csf0NG8Pv7+JE07ev6nGOYqHHwGow2+r0EIwPaf2oCZDDGBGqWLk9JGfJ
pZTSdI9fQu2LkvVY8ipEkDSCn8AdTaGWHmtLHlz3TgkGiyEiVS1LTO46FejQazLE
QWAEDlA5vJm6ROM/6KxOjtk6YXMjMAKAxYoRxk1pZeFrv91YVxvRiFLmu3cSAJei
v9PIQRUy9awfVyN33m9imTlH6Qng2HFh9mAiQMswr+H2HHMA/gI/bd6/9sgaKsOl
rc036BFH4MsBK41ukUmWK6iik4/MZZFDZpJEDxa9MW9fYABYdPRcyrn/nkGy/W0j
FxNHz6GN9UwSsLReQhmWiXktYXpCO0Q26e2YQF5mmme4YCGhmcY2lQrhAi+Oczmx
OjLIwIGgpsH45N1Ht0pGGvIwyu8Cu0dTXPgw+/8wR5D9+38sSpo9ZcsOTidOE+lw
6YC1eqSeIhnY6DucI8a/Hw3/dqDbbvhZ1jlbIc5ahHBtxmV7n4fdulv2Hzy+FToM
0uHEwLle/WFmjkpN6zjduxw3mgbv+AH96jH5go7hyxc4HC6T9lRi1GQ7YMWU643X
Qdkhz7azrDStJeOkEG4M4dfi4DE+4ytRO8YtW2pMoQ1YhyWcOyeUrgMW1YcpYucc
TjZFvtu06LybSpxs7iSqcQ3+nAynDXxQKymQeoFUAp4krWSckU/0IYhOW4H3xpUx
TJzej02SIrrYXHhJ80teQfeEiIuQ0+C/KdPvfKdlFzg12vFt/nfYoO5QZHNGIffO
1HVjr89q9l4jv+HLktKUg10gFMkBV3u4y6hRavb0O99py5mbtzjrkQQm5TfZUcx0
FaV9jw/1R2fpBqHnpMrwnmwm74cCWJnuJgv4r7p5Ug57uri7rQy9iCWEdisGn5RL
hUbZxneB3HVgYGhkm/izVGemN9ifzeSrN/nFJsE45AwgmCe6cQRYETKc0+mZHkJB
x4q8KDu+0I7ZgI6wNsqgbjIAotT9VXhjO0+R7PDi03RX2RKb2QW0hDLuQa/IhwJe
I1T3QIaPeFTDY4XOnpntyEnLA0b1eb68i57oCQAwMlZgfFK2Y5kpPMmDimDFti2f
YDUlGpcy5bBWPr2+zrQ4FDocFJznZ7pav5+j5TEAFOEm/yXGltY234C1sh9FlnIr
1BnYhXFshyWpBZIVI53Es58N7ZuSyHcYPywzL8llAjQECByHekILqIZu/o0KK4hO
6O5vHq7cJEom3sED61BSGDh/Hts4lfn1RsS82tbH3iRRIyvtMfQOpUxWjnHaYw4T
JgHkBYVoJr1C8x4rfTi+a9zP14bGVE7ovy1a1Cn0DZpuyfy0CFqYYF7jJb99NNQW
qWX1Ctj8dtz8zzvV/3h+pnOwreF9LAjVI1iIpcZ8VvYXcCX9jy9ylJugLdzahYOM
Rs0V0qDtlv1zz0BbJ79QZx/27GRqJp+oGDSj4/Pb+fpBk61m/hRJGZabGrOngZAO
tqUQw/WcTr368SlkzluDagHh31FTfBNF/MX8sv8JUMofmBxotoFNSPERK3bDvaVh
qUILkztp1gngSipgUaX5/8BsT+gFjaXPrIwh7ECsUr33Z9KnGUbXx3rYhxJWO6C3
6Kj81obqKhNAosiAgMIr4zQCiOJvd4EaJnyTHHqbzk0/qi8NKHYVczxrtDDJQk1R
ehI/deNsluLa9UW5MMseSRRRRq8Q4kPMFWV3AK36xFL14kxe6fujNVdE4kE+69NU
dg5Z+9m07Bk9Rqx/TEAa/5rUK3FxCLdQL8um7jPUdGVGJknTFlyOiaM/fsvdzyQw
q8dCLXrRcmhQY80qqfbyRvljysyhBXcVxKldaJ/FaGIeprGPtMsOdMVC8jCNA2Kb
j5KGdgnsr4yRYRAqGHp20LGqSY7AvSxHKg9Af7V1+wIShkEn1mbhRs2Ht2SmOxeA
avsaUibZeSG55lgVW95t3fa2xCa2X6zID/j9zK7dyOKpAWrlIHXty4OHIFwMSn3o
eIIXoaHEnAOWdmpSI/9RZAAxxsrKd8s8lnQy0DIgymHMJjrrZKfa0b1L99oHVRMb
LFAv+Pxl4QlsVjas3SvJhiuTIWzBKYcCPNOE3rNcduPDyV+bWzNdqr/sEdHtXcHj
o+UcXGVq0ONbBt69Yeuz+xDhTTsCg5G2TpbHPYdnc9CIl2IXxNFaJuO5JNiu++w2
ExgcMMLmgyoIQqL12bumlxdNyfAz1QRJPceK2xLZ34WWM8VWsRDClsQniy8HZlxV
JGVUh+NqAyOpSyXqB/SbhsZCG/tYNH+GUi4rEunlV/RrmRhC9x/3dCzknieaxACU
YcnYim4E556k5jm8eRs35fBRXl4GTs3EgpBcCk+3Iq4MBzsf1rniqvCjCStIJ5HQ
8WcdtE8zQvWqyV2bU5LbvHJd/jqD1NpO4VoQcVUZBoM3gQE7kWjP/sDrXW1L7/gF
8bu73adL6WtGp4Wpp0klXGbqY1VpSWwxyYOKPwNVzKs223M605pqyNS0/CzKIn06
aCIzOdzuAunVY5H0LUfqvehX0ww5l3BTggr7SZffWsB1u3xc3BJA+lMkXUfaYywb
MgeeTTYqdP54AvIb2Jo2OrfrdXHOc1sM4q0PCSMWCs1+toDSVtuulPi3fqpZMVYv
ErnnQBa2xeMC5IlLn1axCXw/f16P4mQ8SlNUIc/gMLAlJRJgJ3OaA9C3QMl5i+X8
c4vnIFDXy5pExtKhVQqziPQZ6FZ85s+wm+8RE89x51lcMQKL7dB9gCnBgZmjZa2j
PfGW9q+rk+FXFoIyy4jyUGcoZm1YtNkJIpxBUZSGWU3rQlCd1puOyFXKSCYXWE7j
WdARSO3LIdnwyhCnnVbQBcxgRFBv3RK6oVq7w/0oA2ntgxnfArY1xUgil3LtxYHj
N+Dsx3YXR+Mse+g9HGD3HF9pX8aQe2IScCie8WzqZDNhMiLsxmcM0JKHrkoiQQcb
p+4mXN+cQq6e5zChXwyyqsmo1Zwmm+z5JMm+1vNnY/g7vKxX3jbNEozEEKJHUAiF
vUPcvYX+MA+NKUxWjflPPFszpRF2qbsvKp4mA+NI0TNZkOyARRojbo5vpZJ7dJd4
Jfbeg0m1muCPS+hCC76kBBJm6wVgwOI47h7O4lGYSBxM8baGH8K/ew8dcVunrbKw
5ZBCCn5bvNN2i/RPePNpT9Nksthdz4NklBbSfH3nvPurRcMS9P8X0J4s96Aaax3G
tcEplE6AgF64FPqbtbnnpWXxJETqOIMcAbtcTlAxA1WRgvKuJfqHbD5tzjWiidG3
X9W8trBf5FnH0nwW8cnyeRYMv7FtH63ZoGy/T4ikGp8FCaLG0Whhc6Cn+busP4Tq
idbIiEBiQCprzH3aFOARv/4EfiyPAer0ctITxQeNuB0tMTiU+8v8u+wetBhaJlo+
a9OSpFOIoku6DcrjwSxX0yqze9jsjiCBEufOAc6b3lrftqjh3QFyttvfAqdA+lmS
keuRG00NjJN2solfch6QbNJ5gzgS2iA0iwSziTnZOehgOssOY9sEHttGEjL4g7vx
C0XyBNmMvyDww24Qeb5JibznDBu9skjN942HSPNdNlUsnE5UZ7VFrCjCqfR0PF1M
wTQOpUVS4zhdXNJfnA5fI6SciYv0t62WIdXFIuhWY3Dw5R4VSME3GUxDgRC+UPvE
aLTRBSMWZ12D/xCidBOQKQR0VtxX7SKO7u3qJYvnbHy/YhGYIzRBYRsMN2tVFtCp
l3+/e8IARck8TAO/Fl+nCoibRVZqbjQ2dXgiq7rDbS2N6xMJwsTrf2NDA316dxwB
wywmv1tF0/DFUWrXKm3pkTw8vnBsPPJsjSrv5tFTSiiHbW7DQzbJot8On0RSMfiN
ovf9QCJm6555S0QwcgSovaIBzTLjJEcEZE5jbK7vLo3N4SAsGajObPPwC1SwTnrC
nxG0xXDJn2Bk6QNPLXkV56Y29aVeQCcVLmEsJVcJeRuLG80ccYTwirsWGgUiz7o8
uT2gVe1it+8CNYNd305kOxKBAEuM1KPFbJBxIyABVT1XhQFkNLVv74tR2h80SaP3
obDSLryszkAjIeV0pkBxML3nII1pXFlHbO/vCMe35frnaG+bXridBWXoESwRCWsa
uoTzj/FL3w/up91abshkb8WQaroMW0vkxaUVhLsMLKZr9v/kh0RhCYPzg5J3FNU4
DbJJDFqvAVd9VLg1OxCZhXBSgE79BGRI38yyxL4gbSWdEOY/yNEQ3P9AcdO0zQks
GrFg775w1j1Ntg62yKDueQfY1RFk3UnIakjPywEdrdcy8ryqxFZLXrDM8ZxeDHMz
YzuOFQNzceQN/znMC4UoiboQ9Nz2N/F+PXGiZzmaJ0psSddRX4h0bt9tJHvorqb/
/l36zNbyFw8t2Hh+t7Rb20hyNfQInUr1vM26agRHWDIpFkiRhnj9iZ2fzu+ydDa9
isHx6iEkCrKxpWu+go13xhxCbZQicwcEGXyAHaS7gsNXSi4tn687j6JwHAbdAlzl
1HFug62QDDzyfU4T1pmBIhxkAA68MxRB2UCSN93Bg6jepSFWCQK3N+Agx4AGR3cw
+dDeQq2hyOmTYVjHwIAE0QhPEKh13pHjGa34RwJL+7A4oeYCEfm48OcRH4wJIZfr
w9JirSd6kNzBEsZz5nyiYMpE2YhqChGr/cNGG+TUUJKiIwD1y+tbj6ChEjRrODMl
mXni8eean2kXdtR8RcHhVIjatgt4ENZi0C1y4u5OgFAm/lqJfOCSjYlTNqWRU73B
0TmMzCLtwoawxMstwAKFR498U/8q/g/ERJdOGUlIM5POBl0nvmmKIJPGlX1NYOU1
LzXelbBUSHTTHnnqR5Sy2rbPOEwnXlmSlo7FkYqdO4x+b8B+BxBBrn3sXAeBNaDa
s/Wgw1BILFuQ0+QenKpoULBfdaneFP/bS/Gby0BLsor/8Ab++XJVQZ+Q1m85bpF4
OVN/pwNHESvptjfNSr+xm0/srTBPyUhItDzaSJtycuHH/1aBJ622wZlGGaSKC0QJ
49MHHYfbFTlAWWJ0LqpZh/2IvtXAsLApfNSC/Fnl2AN7lpUrjEL80EGRbUNzCvL5
L+9J/B0so0O6cKdG0BNlpn4pG2JgXMjZpKhPsbKSEdaqKUZg3Bllt/vssZ6eXcFz
eC0ELlB7eLtsOFFDqY4c57AEWXYdF5L2xHAy1XhqePbb16ibBt+vs6APjxckp5xp
OoTZQUXZWpN9b9hJWq0p/ZZHnD5HP7b9SnH1nvtoL3jpb7XYlxLjh7adrvrwtft/
xcvelUhGRyt/qdViSHfqSly6RwPvPfyIjnlVZMbzXcDH8518XSqNguUtvB/uov5L
Jh2neYzuqHJmzS3+Tx0tOSAcOmrdqKTwi5LUG+CTjL57j3hLucwYaHNsk8P9KO18
LJzq2rsY5dUgz29HPTywCqvvQ7by41y+xmWmqUhRT6mPaBr1xHLqE5zJ1jTmMuNH
FWyL54XMMHVyUzn80Cr4ZR01yednRTZg0iupYT8jeeO8L51dMYXuFwrGUwHunHqv
wVcpd+cemTQy8SmH4on79jXitoD84YfpeJh8J44sahnJayhJ1JW8Q/tLORHQWaDM
8RLBnNN64ufo8+SbomZpBJ4Xi8K0OMrOWtVQnwxqKLO5WwSPjmhj9O2YlyBg2TyT
pYmCxB3PnvbmROzxpPAa5lBJpwzmxCtKKeLpWOEMpwnQ2ZOQV/m30ZEjsVU5gn7V
uW9/0jeGNcc04oNXFWv4EElFdAGVIUvbS2k9HiPdXHuNX9IY8HUCySMEvULVsTch
ih3RPvEQeRTGEMduRPB+JYmXGUJSd+SC2BlhsHVEdQ/C2C2RpOgecjwuXjQcxVp9
y0UyqmBVT9iAiUbM6VseQfbW5zDFvhszp8PjZip276sPMtsJ7IITrAiHLCcLbx/K
FzI9GACR+eOI0VIYoUQ2AHtYuPhbAafVeP1JCr0O9quuMWgLyZqtGD1j8SuV3WsZ
id31RIhm+LTRd3qZzDvo//1SkkLrhMk0co1HTlvF6V6YstRNrl+Ic/XAdFind0vQ
DcHs1n7PMfh4+bWndcnzpDmWeS/WuxubmQl8KgCbiMjkUsaPQrNjfe/s0sA1DNsw
gL03WLwSph7DUzKq0mDL+MCviDCB0Iy3rr1aoaeKHxmSKYijZSG1YZAt7+yrdDNm
umtX8+53IQYVde6uRHQFulUvlry3eYeZb3MZYqi1kx6OtbwS4uZTvq2w6WPUYxaa
bvNgxcm752tSeYeaNfilRx2eTcYoX3Sb0oJigZaggVC71e/+E6/DypqFv0TUh9TG
JRI3OSJi2CGqFObszp/2zeC3IRoYXkZZt6OrM89U5mh35CFf2drE0ECGto+YgmhQ
4y4p+Av5baLxf2z6oa2iYIk+89Q5PuIDy4M9H6e76e8lQupmixac4btRqYUW3hDW
XILaMVu9dcLFsP0MkojhjoTaP9UKW2fHoh/3BUa6OduXLkPvfFW1pofqkyqq+3SB
c2nOmLH52pnLlZC1Bi+68ciP2g+wM1axZBP3dwINd+QdSAZtNd97OZHdYc69jniN
uDSSf1Gyo/EySBCDjwjwetZoAv5zTHBYbsKKawSoQ2ucnp3758MT5M0XvmiAu49o
1eiyqY+k6jKUZbRbY37nvBL6I9Cvok5u0fd7kuz/f6sa8ChKs3g8IGR1NVKYrxj7
/uhHacTH4nQQs2n0tnrKgAmgopDywDdXIxP3zshiT/tuPySDYZDLozSXMmHYdsmU
2TwHby3lSFfWlGmihQlixbgtMg8Dx7L22/Ia8OEzKUM/KAvlZpF04PzAohtSQsEI
zJ6XaCm8VzieJAF4tZLFdt0FzNe3bUOIlWbuBqIvMzna0I3mJjxI+Q9VLBYURoTh
jvccLFi0eYZyNqypKIAaAE6b7d0P5SBcUyuaxsRt7Bljy1lOf+SsVfZLUIGp/Qox
EVL/kRwhnTlnVL1EF+p0AD4IjrB2zEuXoXgF/Gpi6COskrwnruRRhCFW/RURlZuz
qUFjLuSKbY2UEOpkDOvlLdw2HtngI+ruz5Sth5FTJ8HuCsXZX8EFehUo/YIQ7EEB
Ao6SSA3VHne8U/R+39t2PJlPgtxS75+dFuhB0NhQxmMkGGSeJwqubD3i2Nx+M5/7
CuABGLnuXMNuEp1YHGS+CvWheS+taO0IxJsqMz3Zph2RZ1ZLfv6NGyTG+gZWhms9
6NgnuU4X4D9bDuJ3mPislogTu7Z7uzIvU/ac6Kxil2CxLbJ3ubCss9Rvql4r38+j
HfAOlK5J+2t/XVEQL17cdEEu0SmMy77LNvy5F3wYsmu3ZGhAj4AJiJC2j/CdL7Pu
pYzhXm6bak2K4l0v7KSn2zJtXZloxKsxsfhVjfX+HcEs8qhfvk4+IJQr+FDmx/Ej
ikQ3r364R7x56J1+bO+WlMIWdg82gH0vf1BvYFxhZo8GKOAi9k1kCpbzt4oB5FFV
hbBC99jxa0gfs2VdMI6hocuA0d7HtV06fQbZF+pHYpedfInd9gYwzjIsGWfR6eWe
PKdFwpapSbrkujD0KKd4m5xC1ZCud+0uTUtekzvsb7Y2LeZWsakr7Z2gxzhaIZRX
SjXh8BTdzufXIQd0Ode1CXQjF/CXXv6Lc+bi4n/iS4ek3B5cemJwnj9Q6JQh+3r1
Wpo8aTsDJ629XH0e31oLs2cTF0nvZ+/X6ZiEoAN7lxU8XFelhzlZzly5vEuYpJt1
ZXrIZpna/M3QOG0IVXZe+p5XibMREwnPa06e7Ef5Rpyrp2kVEjz5C7ZCz38RrypN
ThnHODiPd1uFcQNaz0GyeMusbjxcQ+fKlXezYrQTXlQIR/Fg5Ao3UmhlVyo+iFD+
S2tjsfzxYcdDuk/e8Q9SMyKSWN75XTKQgX/k5RxuDM2kVPPwUNratz0y+1RwLjYg
99dDwA728kKV44oAW5pf2dr5te8oNZRMts8S6BqKW1bCcAlM0jLMpPpxNp98r0W9
jDMKMKyHlRN3WyEgRFSaWUkc8Dh/wSPNTlpEXzaOiFt0z13uIW6cxTgP05ganf1K
boF2HTpqtHBXlroD/rr2oYVPlgu/AQP0Bg7r/TIRQmSiM8kdvIUtJr72Z8acVDZ/
f3ZfUCw8vdOBq/NTRYK72JJ3NGl9KBN5GyBreU1JXQ8+hJA1ZzOvCbP6QoPHfzoA
wPCMFQMHhACruVmpHiSyU6oLLrCfLfBLhtIcynscAPo9JdISRVssO1CvGKTks61W
aIX+bF5d/tkINNGBM7HsWo3KHxkxpbuEDlF0hyVDZPYZfykdiqKslyKeJlLA/DT5
389dChh6GSlOw9AaJNBGW7VY1FjsqPHSucJhRmJ7HzDp59yQiynQ0oWiHtiXCXnh
nHMndehUGfN6l3UPrkWYdUfxX8D9ywWGrQiqF0hdS4nt8cgGf7zjj7wztzt9KrjB
S4/1/KzxqAFhD1hzOwKvM7zagW9eI6NmrzwaxxCAplI48fwvdBCO9zSfBar2kSPR
aSmuapr0s2VwNSexQ4Jv3/dAWyPsEawHJMLtYmxf1d6lbncpHREwQaw/daLIe008
guhie0yYiiCY1cJd366RXE0y+MF5wLILBqO8r5jgSRD14SL5G3vXCQdhu9ny8toE
Tv8AgUkNvGY5wAZCZgeU7HixJi0R5kdx9HXSJj4SkgOlXVHXlTbZ04DeTOamVCCB
2imYTwtDGvftoAX1gbafv4BVh/MTfvbhyADnwR1esT4JCr0KNHIvfopKwbzedCeG
Kx2++fZj1DSkNtuVlwJNIRZ82i1XeC74OTWaGZhSxVvVTuUv9OmTLcJZsDN5tu5u
DS+yN8k6mOrOe5DIN8Z0EqjUTUJ2/xdDjvfrBGwY/wxI4f/26YmGf1TXkRnIBYWg
c1rvZn+vxf/qhLYsll39gTW5vgTJ5u8DItE/xYyGUpxKgLfXrVFWlECw5Rd3mnVY
RpxcBe+qZo/DXGj9fak/j103LoXwMlyY4bGUYEh2CKye/QTlOnFiErc4eEw+Rl5B
LaC69xVdBw4FAAPvbC8+CD9qc1RvCKO49Nyr/x6kbAQuf80ZJZ2P9lkbYPrH5WR1
jFJrhQx/xFq4rrYqPuXfeQgJdn7WqqszchH+sqpADdQYVIv26eFz+L9YIA1IrBS4
/UzQgwC4LL4d5SisqiCZex0d11FtYXc9vnjfDnxhiNwO9godfHadQVIupSyHcgEH
wddQuyBLpJl6QAc4OPIyHSw5G5nrlI31K1QAwaJFm5N6FkZ7ckmgfcc9X+7rG3dp
AvXHorsXtb3SAjVCUhZyzyKxCoslaxTlhpbRX0P+0yXGrI8OqKRzd/8n8GnHn8TX
whAAStxcUliqCrQR/2GUtyFOtdMCI5gUNL100Nl66H9qYD45Gbqa7uJW3mlUa9eE
lZiLqMrT+lK/iASKarNv+UZD8E9bsROeFkTwVUvDsGJ9dhKpCn00RbPHN8qfCs78
X2xvdz5x9H2y0KxS/0apW8G7dGX+fvNAXj/kfuP3/Ari2OLCZ3L1LsgVBVb/Wol8
RBKziEilXpdN1gFG2RAcOIn9R/zHJdxW0RBLu5JDnq0NtvaB/oUmrazNFDo2jVCT
JTOwqWKp457WQZlWv5SpFvGfqyA9Td1V6RbK6s4SXfVTth7vzIUm6GE8RFoRS9jc
sTWWfvMyqdJ/U1leztpk8b5j3Wq284EVEibKvAFTfBJXGARmoXGcpRmjlydQ+itx
n+KMEIXOqc2dhU9hYd/fqwgSNXCRCQ8BnZyWV4oOHcDTphvlPmC4hVjd7c0jCDel
Z28za+LCGcX9wuH5AcUQ5Ul7oa9cZ+IUv8bsi8KiQx/DQ4YnCky7ec/DWCSvpqLe
s7XAxgXKCaU9hka1cmwXEypNzTQcWKduQliJj/Ci69R93scCxPSb+Zx+pcPtKo7x
ev92P2ECLaK/wgRjiRJndMihFFjtp1IZ+XFcJvQHy0QOL9MFnbvnmgrNAiJWoJKn
0pu9Cgp8nRSPK1tahpXMib/CeOq9/Mi57PQPTl/0t3dsh53TGDrnu+ikabXCZLwX
35wuWfBAiXfAC6scrui9BqELTiSxzWAkc/HpKnPCEIU5C50GKqXmcZe0gIvw7twC
pBqXV8n54XOzARetyvtkqLYK5r9xr8J+1Yj4dOTwHbahC/dISshSh4cJaI9X1hpJ
36uSPPvgHzMsp3cSTayNhqzhqPBj5OCgNP5bVtYOugHVYGxbA6mLAyuEKNYAM90i
Vg/2sTt3o4AifufQM5c1nLWFs4oAzFipoINf0b5Y+nVuTuAPotGObOxMVTtNw1FT
WKYDQOYJphYAexfZboDBOQfC63ultM2jUrVfx4fTZgU37VYhr03nvbqPWdpBR2ey
3B7NA1gL29+EkB/IVLnqobxKP7MkPnZs4GBYKTD3P2+Jxdvy/EjQ9DERSVTLazZC
kMFefNk2j3teVLKq6cKFyrCxZDtCHnwyHTZz0psHc2WGEbsamgI8/c8oZ2r7RqXS
zxIVlV3htM7dmXPhy8F+VHaqJSwoJb+9f/WGyFA1KHPY5GMHcEkSyNFGwrtgrnXO
VtR48LN7+/KoJ7GtSzY7+aezr041/xM1Ow4JUBrZlcdbEXg/7rK867Ha5G5EE+Wk
v9xZ8xW0yRgEj7j5ME2kB5pZmurgcASZZsnpdraUzKuFGAqTtr1OXdLDeX1Euoz/
l0NJBJLypN8cgqtplxcra5TR0QVGmrVKePLuPB3f8UksXlYS/vGEglRoWWnm//Dl
EHfqe6Ogd0JAPYLYUTtzdfWsfnmKzGrAiJPcGvsLRUGBRtIR44FVOHL7RVhiHLEe
7m62v4OFPlHfCh8FK04OcgAjFoShYrrBgjUxI2SFbPyHnPX5PBi5kf8K6l84fWdk
TG/ywVEEMMeUqK1dEJqBW7ldLlDsI6NcLjZWLrMtqgatKtHlm97OpNOmRlVBo/rC
scO9+Joy8NnRpW/uSu/v/ninqlLZYwkd2/eSA+7tVL28ZfNZvaDEb58NtHO6qej8
nCUnDWvthIW26r1RFwsaLfDw6jZ6sWT/0NzcWB92Y7WMN0xkm7SHa418mlzQqcIl
sX4/OWsJ9UwilOmXVa+rWxAXw7AmOF7BdPmnwEZHjoHqCwDDlgS+PqsRom9LvXLt
upr+9ZbUQJ2hXWhUHzeaXb45fpm4TmWVpGl6vGddMsVbsPT2xpsVU1Vz3nAxoZ4t
ynXNWwIO8zzEAHt5qw/r5MmpsF4Yn2KanQPV35uHC1GhmiIarz5SZJ724kFl9iky
pWaxJyxxkhxI6jk5uAFg4ufAIrBa9vg+bqwaec2C59ZYkn/xr4m9xaS/quW9b7Fr
YqUc+BAa8AwY/5ziVFEtfMgGdRE/VkN4xMF59uy7sDtvVufnHbSZmQRYEtyY10s9
qYEZF0b85f0V/tjxEZbq2Dvcsx+wtVbWW4DSzbrBI5t5HyPgxrxSggtlR3EUad16
eIJmlqQcncJsO0P3tRwiehmdu5IKXTydaL+FDzEdsE18nFjUfA9cgE8ogdJhik7o
Xp3YSUqDIPnCKKNFGXh9qgKlTd9PdIoAuzx78i+F3UDdwm+tI0/H55jCXqMmMNND
8/3WWV6CnqG5SqD2W9LLOM4/APKBWbbMfSceHUj01WBhyzBVshnbkt8n36Y+KX0X
wSnHc6doOrEBMhpLSXpRXP2RLaY13e4hFje2NwqTFArriDa8kr7Ou1tr7LZSLtQy
Hhx7Y61+afhNMfahPx3ueWhiX4kpxZ65U1LyOCiLmNSxCInTjJwSs3HLD7oNizei
9INs6H3sNGwY3qpqaHP9DS7NlZlu7H+Wo+gzmdEDrxg/BUfA8ecAjht8yW4avNPZ
yqqeMEU5geeuJqhatWk7SSWwKVmMxsNg6bvTxZGNtFF/Nn+fejV6zr3sYl51yATO
puxrXqJd4+OFKAXReImTeOXblOyBVevN3s0n6tq/J8SCKyBrTtFf8x1EG3a/z9Q1
4vzskZ31apCykwoVaL3vjXSBlHyaSBrnm4IhAfyD8nOhUGKR4aXo9IQMpNvF0wbQ
B411ABJs5GQuGzyUHE6ztXTCf29aMuTmeEYXFe9obd+85o3fTmFQHwhB6g5WNlfh
h38YrckmdQH3bPU/O0mOHOkfK9qMlClzNvDzvkhANTMUFVjQTF0rw457Rd8eJ7nW
0DEGw4QZ4+g+aHDXKLOdtLiW5SdNCaIHkx57sWfPfc8tj0qWJd013V73GMCPSD9F
zQdCEgmp/t5t6rprC/pn8+6RVRrQFu9WpHbtT+bnPa1g+7luP/YYSHB+ispW563U
py4LGjb2nAfdNAWPRGbhQwBtHITnbjZaJksQndXRQ0P8pGpf1klZcMQsDhCLAQmE
2yk5bkemPxRCHIqn2JPxyndlGOhblzD6Uyo8/I/XWDbcd1tP7IYNOGdXu0spVcy5
KLKZCO8YpZyq6IBiPD5WUNO9byp11hBYS4NXXKDWNVMBQ/zAlghEmFISmZuly1Ky
IXy0aQ4T+nsEheIY7wSjVLdouUptMewFljr1p8h+ONKB8wTCISYerwEohej/ujB6
a/u3pmUmB3tbfG6lB8XSzIqc9sfgnvoAPcZQfZiQEY3M3wLAw+8zsvuNjIsNPsSj
tqiK9AterEac7Iti23r9ZVcfeY22mlRa4V7ZPoJYnFOC4rPxy31w4ZArodXmcKcv
9fsSOtK5YvlQv+UloA8d6mqiuLn3O5Ted+IaqdsZ1vKsx4dAHd3Pn4HPH5aZOyv4
kem4iayy9DAzw4bVIOaYgynxBdAiDNgh+niYCHifC3lQ0H8Ttv1r67+u8ULY2LBI
xkRXT4lGLZcgfWiBlAu1bvnnNj8CRZpB3HE9WXtoWxmlDBz/cJtYE4XUFVyuFw1w
Urv3B4xTB7YV2lTe+zP8cgbIO++/maViAN2xC7uMXNGjCYhiRUZy1P17pRMjki+q
jzuk7ZMnKXX4GPLgEiK79cViTDW3vgoFIzHM4OGBZFIAeOgz0rcgFP8hi/XY9x6Z
CMg1hA7EWxnh4CDZSK4XhN4+i6lEeRGyMSCwxAJ8MkxGi3X09sKNH1brofjdDPEB
no+BbxPENuxGcnHfqTvPlXILaYAYk8/60OmwnwD8HO35lLLuZBzt9SBmXAziLCnm
jI+8ZlUbs3+x22eCG0pTsGxSO0eELWDfW7eMUg8zwMPHh6EhezhW2r6TC+uj9uBk
pkt7R3pvaZRqW26BC0wiIk/gTAnt8/Ee1q1riNjvfKvIkoK2Yb2FcNLbpuogeIfA
8F55IJso4XJPuZoKQ2ak49Z0L2p7H2mpqAiythJaiGsRfbeSTGTiOKSVmnuG0vvh
xBsQ8rWyXeR99GzUU2sB9pLnyZGl+S6r3PhwV7FyyXWVtCRfY56nHhsPrOtKa7rI
gn8s0ii8NUSdw0IZBvAP0iELfK164nNwwiWrM82Z9QVLhDhsOcyc5Zvw09RF8+1R
VBSAPCkW4oVbNnLQLBv7OMs9Nzx9r7A10spoKcmiCI5e96MNU6kU3BNXTbbOXp89
1Ubhlbf1H/0qaCWaLNhVwNyqDQI1+ztuZQJCQvayFjQT9gaFDjua7DaFOp4um87o
7C+Uf2PnlLyakWXJhX6WVDApAZ8JefEQYUhEhiAqNPOTVNSBAybQjNMP6+n0wdwH
TJtnxAi6eB/7dIjdUBY7kunmbQl9My2drmdg4gDNcp1bW1BvcXvAmM1zrhyzwmzo
Km5VTeJH63xnRQhANVtYocMyFneuBbnNu8p5Outdu1WxNQtg+rDRt1yjDhuIt+w4
9yzNdZzWfn0BtXRKMkBUQiTyVzVCCzLuCsaVgWL7bc5kWTDiPmg0JSYUR+BTYR3l
1KeZHR805sSLSN4ZKOlurMXhiN1lDiR2XmTv910b+E0Cpnuh55m4PIWPtfG+PoOC
fD1vsQocaaj3yOTjB5KeUWc7U/TnYwhk4diG1tzC/gQ+huPL8v/osSVe5wxOLLMU
P0fvIIAjRWUn4jH8abYoadzRmEfzSSYuQHS+IyKrke/bSdfYNOdc36IkXTQ4FHnt
kY0397g3/bqmyy15koHwDiE2AkHQ8cVg5IgddQq59Ai7aF7pZfShIK3edAdrLQY6
mVRXPGYSASZC7lqZy1ha+7FW4O2iPkG4WxUcGxlcKofTB1qxTk5WoZWS6bcuivJI
SspRCkYUkqsScH72IigKHxohVLCMJVXXNoaKefTV5IlU5axSSB5IidI8ib5h5MXz
1zey2R+56oenTImRsbbqowYM0LAhkKuZJxPy7B0S0wOg+sXFvfXnsIP02Yb6v1OG
aUQnkz2PCn4+jB54vInARvBHJZyflTW73HOGfFKEWDwzF6WAunkq2SYB11YIvv5O
hjmtpKszQ4u1T+nrK/namALd88JYinSO7uzcPAx1FXgEVKQHAXv76ek8bEjYB7/v
mdIW1ulULWEBdvfH37vL4g99VJj9LY9Y++UaSSWxoUFWomo9PAnZUcVgZo9GecKj
iH17s5fTHNqfjohQcqEG4tRnfV6uFdpU2+CrPH8CiBh4IA8xFrjGQmLelHa8n3Pi
MJ0EqQkXz2xZhlRGBDSRUHO3pitKXMTxTsf6UyszbwDhhKuqj9x706J5j6nzmvKp
z/WMJd/Mn3J4tvSrv8r5nvZOcBvgfZcLj+NKZuUeYWaz2boRh9k5YjRVXrlgpJy6
CNSTNtSklWwFlpLnUM3qnwY51JOR7YUOZrqalWb4CFTat+nYN7tDdhWgd74x2Duu
g+NdGgzJmmF6vwmAzYSzK1PheSSfGvmcwTN8GDn7OH6YCq0EArntiMwdufB1p9SB
77TLHxm9cVnj+SxpH9Q0JgvkVnVZv2P6W6Azq7eLMmOsWO6vbUkTbZNp2bEuaNID
CrT7/6C2HoxnkZMSt0IFN3DD2K5N56Tn3nkcLGuvs3h9PvhbMWX6tqstz1XUavRq
sDwhUdxIxpfoLOKw+8TFJssuGhn8dybJeZkLWAUGwqpmiI+Tfh/E6oNHfE7ID908
b4rAMcYRf+XtPEaKsmHevBrGKq75EElGRsCzRTzSTHyIabK7xysqZLSi9lolmO1M
fpodDQdo075vgt0vT9qLgxm+DYzwAtaJ18QrrdCU+kh7SOXwUlyyVbU107tN4Zw0
O52ksesMKxyzRgHO6maJcpPzwvPWDI7GmRXvvSPs+j/PTPnt7tmdXFdL34c2Rg7N
uAaVQZPVaI7NuUwMUBeNhtyttkJLjFV4ywcspB4lTTgFP8Na3W4+Iqjlwr6z8NQE
VzbD/WTg9rvDFYBCbFMaNUdqDWqMBHlWXw1dtjeO0ycuSShmnLYujmXAEiVeO9WQ
GHvfa6lXDmAxWJqXX602pgjK+Ix4sUFMxXK/PWLKi4McTpATqZMxChFz8rxiccR2
eULyMSNRB7scVnlWafpyG4EznT204pfch4mC1caFjhDG7bOk1QHIZDYCe6/evMrT
DnqeLfwmk7L4CRuvbfH4m6dsuqj8i6ULX+1hFoodn2pj2yWuMtjM8LQDYAUfSM3X
EMxXKnzNUObNjdUm9xjCfIGpJEEAlnld6V1m989MJx+S+v7CfFHnC5FwCv0d2NU8
tbqw/xa6aEhR8RYuqqUNfjwmzUSSHI3PM+i94oH0W0RBGZypDDdBJJ2BzFy0FE9o
cvtQh5yWuU1t3mjm4nRDaBEVX4HEhYN1HG7U+yTLDgrOufoiLTBzzkdkibrkIkIP
l/iJecpSZPatNwdojkqUuPCxqg3+K2ndqUtFVimbQtSX2iMMQ8+ssaiJJCnGc7fa
IH/orsTeF0rZmZ0uu/oXvCnH5SDgOQn79LCHoSVLEWvgMj5lKullponLXApmU8Oo
uG9/RnEMHfWmnGtoMJKG+2Wq/HY9FKE7h6ZAfghBp+EUlqkMR8Zc2mfl7TbHN+D3
DmhJ1OJcK8Z1DnytwMofe3B7Gy4w2HCjYfFh+F034UJ+9oWnCZFN0JPsHKgg1w5M
ojeFnbm3kWdx3BphRRFjT4bVzE3709RyeMtclJChsWx5a1areg8e253Y6rJmGO+p
C3HZyTBPFh49hYRGaMiIKfo2Trb2nO33p/A38XcVV73+LQCidVz45h43usptTnQq
LVHD5ZF4lVVgK0Sdvgdw6NmYgYs8OknoCggd1urYfsbw17CfpZ0iH/a4swKQgA4k
dvtsLGR/77IgCw+SRZxcA8DScS24gChk8JNYKPZCXbF/PfGbFyN6CABlNLfh6igB
RU7ahh0JGXcBaYd3qbD03vIP5M+sPjoDxEQa4vPtfJ3P+Nblj782Yv6VzYA53z51
1G/sV4F/iRHbeN4eXrDH7X1H0O6UfJ+yHmS1p1x3TCgArZWDDs5vO/unm57ZDAP+
fYEqq6qfqrST6/ACOouJjzQQ1ddrPF/XyP/sZaTHAkdTzirKhraVRzlSrb76Dayd
2AULTYuWxQY6X+1VezAQ3WycpSBmVaF9OEsP0CcNg07Q9w5sdOgqQDtKLdkUkptt
f78E9lE5laBpo1TQZ03TAJqVPX45XrIlJkDDugB7vOVqdc2o1E1k5IJNFtY4LCY8
+9zaD2RmstX+87vDr63PZZIeg5jaa3otKtWp5NnwHtbYE1ptyW5WD8uEw/l+1DnO
f2J6UEEVWv3P3cordIPKkMhdRf5LYHX/14w92dNSE1dT82FNTA5WkxX0cSmUBTNV
HHmYtW7ZbFcHHD8jbKYXFN8Eu9TmKtdKFrtgvHXB9O1uCfr3TcHDaQHynXp287FY
usL5uCYz0ID0IbIzR2AIOLXALA0Cgv6v48WGjn5QKT4IBfiK3jjVN3h6KtRzmhsv
roGP/D6KqgXt8B6eUXY9mPIFVtgeOAP8T6+/jFjbsNj6h8KOAQmiyxvjRajCLJtD
xL6/TyxU5rCB/r8QvBj7UO856aD+2ApqD5094ERAnreF4XcxwRC830jwK3SdlNp8
Lj+R9lxykUAEGR9440GXKGsKSAwhC4AJFyLWD5OeDfjuh0kGNg+0RsdiPoX0NK7g
mUaf6839ioaEKDXrYC1nfXEQklsLycH37iJU7i5HUaj5ZYbzghAENTlBB6P1wsPX
xhbi1AsGfwR0OKxZ5KOHCvpTVbrH7HtZuBvWNIaiRabmKNszJ8qTs2X9OqXZJ1Zz
Wws1j/uFO3zsuo2VzUgldW5N+mUSJFPInr1Xk4O9Qt65As9/dX78ij8jep4D7T5A
XHcrhl3or3mCWTFTozBOxbrV5P+BrQJFyRSKfyVFA+9AsyXzaOSoCkQweWLzZoKP
fUqehAIaQ//zpks/mFYzkMUz2twig4Sq+Jy9HbD9PVXQ02IgxdFCMJWuqLZwcudY
R1T9YuKf4+80CB/6pMkwiUq5ipCCyVYU3/seB+BIeNxEHAaObXl57N0bOIpgBcET
knexTVVevQhp2+BNMAkY7Y3SnuXVSUtlZnr17baE8S/ppLVPoKAZKs0id8ebrDMc
aucCT6Ph8qpyIPWnFPYtLfMKkMpxXwZL+gWf4nxEIEiEphFHWndHGzmZhZEXvou0
iZP6pOsC+Yew42IH0ZqdrLJGDpLAsasgHSUkciySNmO8qC0wIizLVB12Tg11Q6Pz
/E9PrrMgxXNFRogC6Rqd7r882ItAtHkSQW8jxe6ouTU97G7cyh2asSotUfzAhx0Q
yfZp/x3OUEya7WZhQ9Vzt8EZ07MC7UBQrbkG7/V6ua1OqttazQJvKkKroPZqJqwV
BAGjn7svwxyXZZwiFdb1LTMGV8FUgIJctEsjDJ3DKzgpCafnWJS5kpozzWa1SNRr
opGalmIZALxTZ1s61aQVhseFpA6Rk3PutGtolFBrnarJuJHZnZdrHRDxjH2SEgiJ
4o0qxwfrWw0LJzgZ4HQB1WBdwDIgXGudqVsso9tpZ1iQuaj7SViJpybl24nJvT1g
Yg8LJQKfqSccfq6/rrcKkPV4OyuGWQwIH+zQi7gtAlCYdhsgypZ2QsxvviUpNi+h
HNkTHWGZIkwesJdhDsyBEcopeN6SfgzYym0h03ENDW2qtNuziaDnJcUcdjUDwr4z
fYahAx4GJaSsRCVa0EmSQebiN8CN0XuWzm8ZtYRnfHe791bJgnDfPeM/E83X+vg9
50KVgwJPWPxaVUzJDAri7wl7MFE8IsNNe1ZbqC01HYsAx2r7spcqHp6pXx0hOFSZ
gUY+wp1CurjW28Wn/7MGIT/Y6WTgmTxlXpShbzgJ71ptK8c62aK2B35f2w/jOHyb
Q6ntiKm+fvHSAB/pFYl+nVWbqXjNU5/yKH62PJRIOhfAEmSo77giaEfJ+U2qg2Dk
eVpgHCQbwpMPOipCYUinXLkTHEesugwvyIETtIOJLS5/byIgy4Gl8otxb4Llzrdm
KV3VWthZxNdmfDYf3+AaYJOGzDK+g90XXbSH6dx7TCpZem4LVyq8dJEinvrrC4lR
Y+v9s4AL1SiSbVEseuRxp/TF3JzE7Xl6Vu3hWMQDdvy5sneGmgW5OEvS2NHlJb9G
e+082yBLaUrwe7QHGfz9nR303enZuLd4CB9RFFpIc6kdLYhHt7Onurhn+yhXpJE+
bub4c6kNS2I68lGMEoJVDCc/dgw4p+B/LA7NfvZBfFcRBUJLCqdjMla1CiBIXJe9
IglRpd+ZaGhTdFLtGN9lCtllLgpwtHAWp/tFXEZUljgvjGrGlmDbp9FgZaWTQbtq
zNG9sOKz+2RhDkfi8DxO9cG+VigR2GnbtXIbTNVLGJ/LydqIwSbNdKNipfBEb9fd
1ukvF9wKNmldxsQCkrXDKXoghjhz94NEwZhtLsFzywMdbhqUqqmfqWGOJUtL52Eg
VcU6//X3sVIZ/si4SWJ29SW60QSMRtKakQax2lIhQa8JHXleQYga189v4J39izYb
vNPcBv4yq8Ho3CNL1GUvONyQyOQyR11x5zc7g2lf02KpiEEx3GVxpSImFrjK10GA
Ry74peBoNIc8mpFlF1PxqFbrZzayMKSijs21uUFznN7Ek3qmhztWBX37CySd054P
V7HjQ75dSxGvsFmkf0wJ4Qo5T1TZR8vKw72NYt+2e2wdFPxeBmz1FUJcnQiRYpET
Z9OGy0rSjuezmCh+ex9CoS1KwzHTEhyyVdEXVR9IE6RcBoSLoxyF6z4oPhc+P93C
PZiIu2blIj+QWCpjudf/GQV3HDwgpbFaQz+iwtowmU5m9M1Y1DABCb0GsC0FWXuJ
nnja186Vn6BRNJguATR1wk3f0pwdgMrWeH9dsq8dk+8rOwQTrBXXh0llNNL9SpyA
AWWb+el9hgb52MggZdtuPOcjQeghe4dgByHTrMwREyR2AdrpbzbBKXSo3R9lEqUj
5TWr2K1S1US88nmC1o8FflS3FsXeoc0a7JkHmdmSp15FLl/u8QiVcFYTSBRcMTe+
28xqNsu8u4w+ucR0qH1wXhZp11wO4ltxFj7DWbLduAkJcHznjUWQQF+NpyLYAbrc
tPLyIezHu1T18kMTWxStJAOwimd2cP90wXtb1fRXeNkSdj3NYjEB/fxAuzDj/map
lPmVNQSl2vGAUYUkFCmCVtVVovDzH0BbCBfSdxez7olqgZYyPF1wavQ4QxquWqCo
FIWe06Y2OMz42KwnB/Vr4CWaaLgEolUQ3SAiy+avKFBgdzrykiIKbhtDGm7IejGJ
OWZ3fTbedan3YdDop6BjovT4SBn7FvAHXIuxYxe0F2JMf7iiQ3gkZjjMRvd2BCiP
hsfViC7N49nahWvsxLOb6Hd3xk8HS50eKKdmr9PQMiGM99r97zg9FLWDmzYRKZni
4q2iQA+X0elBl38sVayYrPumZKKGey8n0sKZMFOKkKOD85vl7nG8kYnUPevtwSzr
HEyPjPkmXErcF2sgaQJ/1DQZvp3W7AxLNJ9Er0LQkwBcbFC6Ku0bNss2MGth9DYN
UMS9p1Q4wfw4zOtG9KWwT5MtlCUsFgrXGej7APYvKqojya5hGr2PLFeDIjihobym
D7CHpJs1ANHow/0ui32cG+2L7be+uVBgHBTLGlSTgd/QEdsfV7hCYm7q2HLq2Bqo
KONPCCHeJsmOCLTrg9CNEF1YgjQPhtpI9WFNh7ZN3UI4xTlQVO5KCZaEqR812Jjd
/0KKAb5LHxzumDFpGPXTfHGOjpcU8bmXrn4qSsR76AJgwlHJT4vl5vYCZ29Ol7SO
dijKaPCjI5Hbc8bPmAOXOOWLMrz3uZEZEq2QtutyK1OLUltMIShxIeN+3Bn/Un3h
c8KZNC66QtEhAuX0qHjVOtF0G5CR6Ry5cCyNtD0dBAE6/s7Eu74aXRXxpXxa87Pg
Vc97exgg0r/mboRhABuWngI1VugLdoVegUYtv6kUSDojkZzfQtagg0/xx/NJSaYJ
sG8DIpF1dQhxKxNOLtTKCTjKd+IoTP3zV17HYVlw9Suw6hh9tGOm8Y0tbVqDW9jk
sK+p5mGP5O9WwYOzJeQMPGYJMIqRveQeEx6e5uQMIKB9DmbKilN1ocTOZq/PhDcv
isoOkJBBP6lQFE2dQsiovnB8eYyw790uZDxC+IOJlsRhoo/idEcTO5BxfcvOqP6y
Tk/lze7kkYtLFOK6iWk0NVlC9DEVi62ggW+4VGHOGJFV8ajgND3szynzQs3gsHTi
QH+qb7QXdLy5X9e2YqRiFv0NAVPV45Lw8vQxYjRiB4aj+ah3gXPeIbarLI38XQEE
NSFQuOODblmQJU2rJyZDJMRNCFt3tDrd+NCBahDuGmoIYBNmnXLBZWk9E7SlpKl/
F8SeVcNz81WI2uM/8DD5U0ZUrTJdBnHY8ELaAFhZZdXFqQQByMV2UuKANwLSzb9N
SoOSb5O8quTyevYY6Gh54rjJ3Pk/lQfPx1ChyeRQNAR7+wX3VYlfOi947ZmgPA6+
/zqkPHXFFSuXu1yh5M9qmEj1B9QZ+zglUC3SAhi63/1Hko4u+EhwAJnwhUG82Gpc
j4bojqgKANlUNqCeWHQFOJDUPzpB1/s52KZWxE30K8OK8RVg9tehZi0nGiXAJbVf
Eeq+WnXhFS0++5OCvPcF+lvZ/TIMlzUHMxXWuwk6anC/8eXDE6TpcsI+fEOns4Jv
tyOhWfCugJQn0NaYA3JY1x3/7DmaOhStWzK9ZK5Lq0J4r0c0856japTHT7Ee6sii
Gi73Y6ppFCmuXepnKe1vNoPhax++BgE4JApBBW9gwzs6w2xiN29z9gUOlYX+z071
ExaDPlti98bhybcEfs1QKC2YmNFx/wxx4B912L/i86sxmB3yd5hCR7UsPl4+bAMI
AquhZ7zdAwUe/ZxedDO+XktsDli8mnwjJEsIqpnllg58bu9gILhfLyw4MXjfdbkN
V5QhjrAgMKx9Io9Al+juHxT4vaIOWdLguhp4T6Q0mBfH4XRF8BLM/p6LjOzeZSgC
NQjM5EHn57BHdEMWvK+kWkgG0ws0O33OWWJoVmX720At89QIMrKLKfIF7SPH7fOA
EbjFYl0JtP2onHpRf9//JDI/6BVrDooGC5XZa2diya7hHugQDLhHx39P+xlNgvLo
Aqs5UmvwKic8pbvh2w5od9JJYfMGcKnjAlsjyFotgCfbqz36C6iDxFCzh4E5+YS0
ws31l1tPn2G0t1FNFLinw1KAcPJNnUAsCDAm9LQwEbv3d9qI1WjZBj0Sz0OF9xcl
XchJEtz204maI2K3AzrB2yC617XQ/X99Sj1TV62I375xwY3hBUwA7wvUx9cfJ1jY
rSmAF/wEuLr5v0HJHKm80FnEjmkPfXKua3IGSXZYCM5Ki0NAKH0ILCIhPxYxv7qB
8Bme7lwKsVde0TZrBz1gUnGKNTDc4cA6aS1BUSBMGuVNTcitw42EzHQTIV+aWw6n
ex+FJ91VDauz3LscbDFWM3mUYwHctyLo1EMZo0YaoXNidFiu/M6H7kEVAJcZorDP
sIZFOXWXNFP2iIZcFawtnbCTcfTQhz9P1APTSRgYL+xh3j+EcQMUFedwxzzIdbjv
7z3eDICu0IarkPWCHWL9hWNp4eS//E2KBI/PbTcB28ABEejdXL7IW8uuu3yeFNjM
cj3Is/agIwpFtFpn8twKwBpEH1IXSiEAPSmnkqjSe4neUxUc5bEojRjPrCsw4Bls
n2znnscdFg1iIuEgoVQoPpCWkFvDWJLPLQKf/JPgMJ64bZFKzbch/DqWAx6Vizq9
5JR6joDduIOvU+Jtmh0e3WwTQkSYwJ5ocKYtK7BbvYyUojmhcN+okdRmgs+s12f6
Iye4eXVVte/10h/UAI/8S78Tz0ei3Yh1SZl1s4l8J5NHaXsotIW1McCjcwVSWJ/V
vvDo4cNef7Z2IhvywjDWsO422APiFy7PVuV6J0i4qzmX73nxqDwRmf4FcnSAv/wx
utvUqMlMiLc7EVWwl5c4znLGRH4v0nrC/kyRxAmBr6ytVyetHClILlpJv6dz/7CN
c2iQj0Z+6YyZeCTKTO1dlRpeAYgI37nYrj4o7101flvoRl3AigRunEilSD7d8RYv
8R6LnVyondayG9ffAL32ISHJfCc1gb8JifvSRZ/SBf2DkB2W8Y5jjUea0vfaxhaw
VqDZOYi1eDP1ifV8fEWzDFzGgonZoCEPoCmY5bX/TvBX2cTIyc8yfmqpU4EgEQwt
Tnly4tf5y2AXPIOsY7K2pww8Rcj6taMBDaG1+SXwQ7OF6dvA4lh/cDSv1hhLFTx4
QM+bqyTSo6O/RAVIeP48sgNDy1j5YWUdb6l8S1HOToKw0bi0Uz0Y1Z48xFH1vQ2o
MYmi6PaZzc5YCIz7QtdXr9W9nQqk9zabDpY68kiSIII4Rtdez4v30LigcMpVAVqv
i3B5KvQe6Kf+Ugll/aCqvmdMtEEFVhMjsTg9MPhWGVEhDinmFJl08OR9xe9Jps2b
F7bd/luv6AKUzPHGySwdKNcxhum07gBpOmVSoYek9cUf2Ge1iYySHaXpKsZ8L7uk
AVA1qvCxZKL1AsMOyRhEpir2UECw8tm30l0LkHmUwD/WRgX1yQlZl4s9Kouo9uaI
d2wWaNQA/IZTFdb5hk0wumlyBEZ7/OTFk8fzp0fKab6ouJgBVwiXXQuFJjmUKx7V
cl0BCOFHZiu4/SgrSIhs9Y/7A1jnbLVsAIf7AuhZdSiN84ZdgCHAFAnFSKY2bGdw
0M3jq7TNJr2BbB8lgqnwmVmh4Go3MdyYSj2KpGahUgVOA0ov/9MXeRMB+MM32T5q
gmDixH3LtPf0cOtSnoWzi2JJ6ZZgXZmSR4sqzotiJKKZVp31Cqd3rm+bFsAlFWQi
tx5nrHk5LyOdYg7VZJj3yQkDV7C0l8SEbV4VSMhMjcxh1Gj6MFs6bahzi5MHZ2Zi
KuU90OZSc88QYpUZlczc+z8wN9ybC6eWPBkCoa/7flxgSzhQAUm3s6ApQXWGPGMt
hngdIioNv8cTG5TCTTLCfSf0K6ntrv4D2t6sm04765eMbFP7ou+++0YtkM8HNF8T
feS3hj/nMKzc4XylIYTpj1yALicKAxhzeQHPoQt23mzUFLyRUsREQk932mf2AstG
zbnrj931+8NxmynDw/QYy0GIDUO+lKLkquw56CW+JhB0EaZwECKVssqgtao4lnCP
te5+FvafvxLECekCgAKG6dJrBL25g06riWJ0R/VwKeJs85kDBxiraNrCZX6HV8q7
t/a+wb0uaM6lN21WGhiVnftSosJ6DcC+/6RZqtYK4J19a9pWLPNWqB5Br0+dBctw
7a0x6RZ/IuQv8vHr3RrWdOuf0CcIRoOlDhYtOhLOCjUBNxMrIrv51kbsQgGm/S88
8XJ4lF0O2xQM6ByQIpgVQ5EAmmdRCklEItkeNgp3Ysj22pVwQCoCp5N3dn4ez7IJ
Wzz/+tI7SJy3AuDuBPYjwXCLl7+pf3/DxEHq/9qoBv1qBJshMaodL56XVJR0f/B0
BmqwTyX39Pv3YuO+czf1XCHxAiNPjoxXniIWVRzlb3AmNhvM0qx14vALzudKi/3C
cWO4hkCvLPpqQE+yUo+M2SNdYxb8tu9zLwtjHjRiRBCb5uGAQ2fLkkfdXW+375yB
060Fx1IMvW0TE3G305GUtka8y8avhau8kvJtHZAveJAGl8g9BZX/+Gg9FoASdZHu
p2aTrYtlByU0HGQbEO3bpWOoGnivFn2onpULfQRzgD6KwFlwmmlhmoqLgjG7Cg7l
FdN/Oqe/KbTODbLAN2MjzT17fbLzAIxtKE0lf/cTUO0GaoyUvhwh1s9DdCQWrIyU
/yeL2JZ/DoRXkStszgiDGg8Yrs9Lckma2Mi/C7NDAmVatEDs2GdcnS0eOk3CSe55
oNiVB9xJf5FJb7CX4x+CBWnB5eWK8VQkTHUnpa6pejgIriRjLtoa/tLXAuNmAZ7e
iuHacZjOl3kiNdfflLSdnr6FHR/ECQIJ/tra0xr04KC7q1y5di6uVdkN00JCDD+7
cDfNgtXaLsR2LZUwV6IKzfgQSTQUo0+/eTdsKUeNNBNDfw+w+g3htBMXP+P8xv/g
RmA/mE5g5a9dmoHtdeEGyjjztY1GVFpuklHs3ecvVBIIyOR4TVHSPvQPnSWVXsr9
sRfo2i2Vq9Ta5Zyru4i+GQ7Y3wKJsmjYwwJGLNcm/+z2mSBvmKFmq45Ed8oGIpj/
n1HzMS0ET5FjT8tANGNbbau08ii9Cq/kAHZdwBYOq/00ag0d7v0OmP6e7jdV2ihp
nMnw7ir8GMRnZ+AI1zxuPzW80gIdKmZWWNqN5AJCShjZuF87pjp9ss6Wrprddo3T
DsNH4B5PgBUUqyQYaOh3YUe1h88HhgYbx/QI2TOBDC32e4N++B88AQzGVN5x4/3B
hvnftP3EtJeINwUhYo2lxP763whz3FuBQM6QQRpiQ4azvU1pfnW64AOz59loLohv
bTY/QST1ieiqjLFaMI2af14bt9IUSKlvMDQ7ack7+/LdgamPxYFpsmUxIbxec5ov
3knTRXaEkSH1B/0+3rRaLwGs9a5kZVwEuiEzN8FuksbrHBUzQqnm0YqI0s89lXWB
F5cKX8EpWQwZaPGJO95vntbrHDNfYwEIe74IG7YZfZJlcUxbNu3vGOAfSDiwKmeV
Yd2trFJBFeHKOiZOxj5RRhAecuwwnOnfQQASM/vt22i2s0oF8bmKAPIXZA1RLaUr
Iz+WibYZqFV4WvHahY/3MKFREM2wpBJSS7ytFHA7R77kCg9L3knwEBT/P6gKjXBn
77FerOSOniOgi4ujuPkv7swvcUbWs3MTOOVrODd5luVdhxU1ze5JGCnrhuT06vvr
si/eZCUQrQEXizcDgKa0kDZVd7mL56CpQl+Qrd185i06t8ZvfVPfdpMURpPoYzSj
Ek6fZtB0sVSDnPl4ZoFP3kmy7abyN2c72Jdyls5htsEsqUo4H8FKt9E5PfdGRF10
tYRTecKhyF4tj3rI5WJBbyoMj4aOUgrcPqqouKzlp0q0MJ5TUnuAp9Vw/IBW8gbA
rHWtVhyvHQop02KrxFHnVRx6WiZPSo0oQMCgokCBX/emYt/KNEU+AvdFDJxzCFB3
Pg5u/718+mX5PfunNRFGZrbAuPBRnDrXD77Klw1Ih2xw0w2lcTevl08NZK6J0jMS
lsgK9OXmXsUQhbqCCjz5PQ5aHu5My3bbMjpVNOTdCzMpj+zSZz62y8Z+DZttaYVa
E0r7O/IdR2cyUK2nlF6BWFYn9fW2bqQchTLu0Ax+bXjyB1Bhgi9ad1WfhVFqEuG7
7g73kG91kYVthKhpI188M9ktTRVilMhcP+Uz5x7jJWliyonouUNaT/3KTjntpTzb
cQkZCn3E6f7shlJu9gmHjn4ONt1rznUsGC20Yzp5qpu56LkvDDw9ZNtK6TsB9dwT
RNnTcufk6TVfrUl2NMPZuHhwEjDFks5wkcQFrVM/DlFSsyRVVU3rgwkg0maKmzI9
4RcZomHfHKluM9e2LDoxxyMMwn8PUmNb/+96iDlkCkvhRHqX7RgvUpSJQK6ualdi
rLmd3MNWvjjkUIdSa4n8Ixh1eNbt9G99jnSekzcMOheD/q31MesEmDTRE6XEGQBl
WkcFvB4dgMX+G58ZG5A06KeFpRqQ7Hpu9m6C7xtKbZE4+ut8kkNdzjn8Iqv7f2Mp
4fRQpS0kFXugxWxdRugjnaVfM/0DBJHOwu+SiOr5+F5RsZ7SQ/cSzZrg0eTkP60g
gwgSg6SuQ5ZUQTdVucK/YvylcujVXHwC/PDuYNbTdcuapZG/xx25hxTkHxorViIi
cC6Hief4bTi3iHRjt3IcAyF6SZwyRhTz8C5rx5nB5Vfb6L2HxIS/rCmuWo7vrmqb
ODNHbhtYW6Sdqa3eDSFNZEZxmYQ1NUT+E/GnOoEjfNEzp1ejZxgBPpVhsLJBPoeM
MZOoUBGhBB0KZm23dJY69Io6lfyZY6CS0JXv8ppHnk6v+sZoVnNcgYiNjj3K2qrW
QP/0g8FWXrziNk+LUjsveFL09DsSUTEcV7tn4ez8T3EUvOAV/Qak8ePkeGCZiSzA
VJHav23ebccVyK5tW8nHUNS9atdjM0WBSzszHktCl6hvAOtZ4N9UPef8T1TdWqGV
HHuu9Es+oz5U7BGO9sB8MKrFud716jNzdmAEhwKCT8Jo7WJ+aYV5XEyO5NZjjUE2
C/FoHh66WhCXfuig2IpvGRQhbOIITl6XUqRHX2Vdv8p8J3OdOOOGEfvTAQosJgkw
zlSLcjKwa4jHn4Z1/Bt5zNw6JnW3OUYh/i5Tt7Mww+DXFfx6QYQmjaNBnsLMESFB
ZNGEEL/655u9pHV5mnOVmP5T0RgFaCsNRjTqSZCgF2WjrrVTxnL96roPJ89Y/HjL
XUtkV1kt31ABoe2i9l3bmf600R5vuZJvBIcaub9Je/sClVBVa3K18sgPbzoeLErU
Srw57NphfvZ2apmL9GFmpl0cyl3rQrgaojmNQCESAxNMNb+b7p7tzqfAC1la+TGQ
XH++5VBHl5ZxG04EQCykRpni/52F69BUFpaDLTvjtTYOwW32Yh6l1pJ2cMMFSMM8
Bd+yyNoAhmZ8Zn+pVDKuraYg6qfA0InxOHAZ6p5jWmui01xbajSBZ79liICDKhZO
p4ESCxVbNMKamMA5W5Gg6xLKkPk+dMAs6uKREdPaPHaCOpfJseNCsMCh7IzHFFe7
ZL5Ax4+hSe8AEh1JOqPAUi9Bwskmggkq7GZpSGBVFb47DzB56/fY3aAQ92x5czoT
zcogufY3ImDQZBW98GhKVtrtMP0buJsT0tK23mQzw5HIHvnQ63vXJ2ZFinf+JEY+
E0RdQjUZLsAyAy0J1enL0JV4noVi5l/pa4wcHMd6RCVS8zNuG9BOrLIjNNEGpcwo
JstShnyhO/2zn/RdDVV0451pCxzbjMTqWrKdZA9iSlQ+S/QQUIcbOlvqajRLqV7x
O8ymZHtt5N933X+M54EccZeXqbksUL3bWUnOg3apy/VkDMoPbwWrXAwjX/hwNIFM
1kYQKMLIJCzOux+QcJtJ/8yJ3BjdYY4mwPb2NjQN6BZwrkv1Sj2wGS+glq36ag20
aRpXMYvGEPdOUC8pSWuRtReMKnHDs3Jwu/MUIk7nI6jgI+KCfVSsUf3MgKFhYZZc
GbxezJJkq/vfZ0CXtn/EbRq28G+0nuL0iN6Lel81Sau7ZpKnZ9DStXXOde4bLAgK
9coOHIq0Db4jDfV8KtmLCltoJWPKyn6Teq9E2Iwmoqslxx/81UAImAyMGSm8fMcF
NuEV614ItLSMCmOwMH6Pbx0O+ldsKKYf0td2lqf8/lX1XOso1tCOFIagfLVwxaIk
t4DYibFmaMImjlyz8uysaorRSTkvN48OOwP2gPRMbjGk/UUHRfh02jR330e1LMmE
N5g8dgNTkKf7xguPaJFZM3mOX8kGp46SCoarSZC2wV/6Dnl2bA37NvoKuIYB8Zgl
D2WYA5B/LcPE4mxht4Gb8x2s9fGqys2lO24i0tEuquvxxOXOwrMnNmAOcEUaCwUR
Bg+QUB1A6o/+ykSveuBdZJmKeBJwPeTsAO01OUC7PgXTM7z7ugKD6lUOSifkgApB
7xXaDp4giO0i8k0ANY/6aC9ndG8r6N9WSmYVRQYaR5GuNbz1gUBZIxU/xGAJVjW6
Ot2RxGQgtdRfaes0s4yFO71GvEQP0PYHJUyQNeOKmQK1nnBCQgrQY4eT2uJ8bgFl
5b7vV1srb7mwDLj0ybDT/uoOMyCHFWMgAOhStplUF8r32r7uZVh486yw2v/e7f8E
jc156+84eyLO7HTXLFgq2ZSjYl6r3oA50AOVgsn8SBS62SJBXsw6WEe2Yrc6jMot
94ZRWSKJK3fh2NDrbYCwcS7vXHQ4zNknJHw7XUUfb82uw0CBo00rF4ji8K36/k7P
FJ4Qx7khf2mhTkkhcgW5cvgX54CqM8gjWbyR+weZUU3myXv4V747eO/YTxcPkw98
+i+Rq0YB5boZu9g5s7CpfChAuKGycAffuuNPj++Q7IO+U4FzcmHInH7FgD6qWhcH
H7owRQvVVo7yrQejOKi8PqDrKvUOmiDpmS43irnnFaRo3acPm/sLG34g0EM/u6A9
qoE8wqkZUTiIXbBZaom85WYNzpdx5wYp+YpT7FD5x5DskYUO5b6RkK2PJJTT99r2
IMNH5fa4fnUIdzK9ZDpqztKBd4J/z8dlqQcPHzg0ExcZR/fRFAkNaLn6gTMjzKv1
HFasPyRYOZwcC6uDeeb2OKWDcT8MG4lGvLO0KF68lPEUfKbXXWdt5GbXcU1D+UH8
snOr0vjy8lOK1MWlF9EnXhTm+QGB9zblChT3O+PIfcX5FH3dUTBa97U2mkFrEluh
sZ6TsOqpPjCTYpNqWoBDzPL2PvzOkKy9jyba8iJUJE7/R5PKFFY9X+dKDOnMSgNt
dBK4y+4wFU0CCw7uQfgqtWAIXfYmv2xL6+fMPqGER6cRcykRKM324HsOvBRMEgVC
sfDsnpRhHcxHAKc2Sfu25urcy0h3/2rmqI/edfeyux+VfrAKBlDh4BnffoYniDxZ
rqwOrZ2+vB3SgowQsYvwGhqlmqzYBWpXmMInsvoqaJHhQdEEiJ/KN0QTUMJPb9H0
N6TkIbqDPHAgXXkEIdyR/iGBefeu90QevNti4eRbEMWPOPnCWilW39HKWGe0eifo
AkzmyIkTiSwAxee0dQiljDl5wpyXePcem3HDlt0PYE8UGdjBWmjXRiMh2lV3nqCS
j4z7fG7F/U1E2P8d87WGFNMFAFAa8Af3DezNqDxExYN2GWkc3ZWzhJX4943Uyo5z
5ew1MuPNAn8FYt9XnQRLPutvoURn3dHKYXA61QMywZGj1kLlndRrZcqFPigySo+u
TwNbUC9/gz0xgrgv/XcZ0mO4hflIoZHCQUXJQ5PAckQUrD4HuLr5cJDI/HqLPZrX
OEsF/m6aM+c0LCv2O7IYrclxFk7n2I8U975OuhsFqK8lKNK7yUU0Bv4/3rZmsa4P
F8ZE3p3dN/ThY4rAyC7fsK6p47Y5In5Euj339PzGXCDACiEECakxWJwPqFPwPzku
OZ7D8VFSD+Ansx2Fq5Arioih3yxtw/+j1ORKDJvSsqjt8KqKylOKcOmBYfS411uv
eN5me0sGMWWKa0Eis0xWV3Dnv00U72NfdybS+FVhlfJz/qK+zWvWM/XK6mQoHj/Z
EMh1tgzBl05rlj4lbE21sEAHtuvbsC8RWu0/QHJmwRCoIBh4SOzgSwMH03WCzwBh
KzrJU8NIWQz3/gg9qRVts1O0287lCYMExWyeVM4xCvVI81JvPY8WjPUEYZIu1qlr
bV1RHbff3krZ1QkRu5MW4UVgLHxRmnTQvnPi28I6DKPwggDct0nNIO33cj4dn2xb
eG0XpJSPb4HSHqaZETYjSiMQg2RN9OSerje0FukyWmqkeb+GGL5RXeauEirQXVRs
+HDGVRFlDJh9qu39xdu61wuxXDRC/wQEMEASC5Ja0aCR65ha5Ny1Oxgrn5OpGcRq
yNXign3JkgptnWYTmue6+5WvgLEAWoA+waeDBYwnrpkUZZNK1wxE2YA4tzPKEkd3
oq24OC8qTpycSiQhwx8SPac4L8W1n7E59GltakaTo4DJ9sH3RpvIu+BctBS6XpVd
D7KfnwAaiBtqBju4/yKM/ywaziZXN+dWE97NSyOKMbkQy9w1Uv9IcPj53fga4K1D
dAsTIYi9M8w2xM7UlhtipYNkmM8Cmjo7FTdjFPKb++mOfNhOg9IfMmRzgWunl93a
45D1VVHoebdoFEbu5QfPaQwvbs/DtrQIsuSQtGiBf4Ans4GjZal/pJxXpSjWX3o9
x1E2A9dvu7rpm1CcgOadxVPWaMd8cBetorez+kkuj/XxrAJMLtZlaqQdWX4YGUAQ
sIXb6KbVV5kf6ZI1e5AYr7H3sDuzbL4+wAqmWwTn7PR0XSZdwU6FZHLtyI/plMM8
aebcuNdx+HVSJVH5OECUJsa/dVlM5Yd/o0RURq53vxooBl9p3+0XsMDCaW62EJWx
/Ygb46bEfBuWrstPl1jiU+51I371VbwAYIBeKl12L2UbCgxbuRLb4ZGlcuVOlpxr
ozQulcyksN1jnilDZ0C33LiA7bVcG3tugAfeMUR/xQeXbFm9igl2sEsyaDVyGbzW
pQet0N811PZ8EIewM/0pJQ28SBl5rAWLdq7bQgck4xk1P1hL/YdZI10Y8gxAIFYl
j5+WhR//tR2i35pC6U0UNxcTzyYYKy1iZucbN/poBJCFBG7P0bDnm2pBasClJwqf
MgyFwvchzS29Mal0ONYQGe922F2vmCz/XJxXggORqT4T6gkFe66E6RnpaOesS7wu
6duv3u7aJ0k0vH9xkqfCMysZKbPvCvBTp/nFClIxcofaHMx93x9ws61ZI+0cdAWA
02i6PMEiw6J7AzMJozjUGTaNsw8+LrfRkwTcE74FF6GERegifX125ipe6uUB8j5c
eDxu/ZAwJNJXYUos2NNktuc50/IEyRQvBL7cYHUI96XbJhpcwfKaKdz6tDK3Y/Ue
PuhtYDt5FREtoz/qG4jpkNFR7+1+MFkrX7Lwz6JzdJsUEeAlpOxrSHdyEtQiRB+p
xpnAGuiG1SM2whXaEqJdpvIfwJilLtCDebbZflB1Uc1vYZ5q+YHW8Pvri92sMZ9y
QDvRmb886HdMIwY7YAWJ3RoYqAzTkTTiBH0ii2W5TK1G63V22hNdXlI2ekEbsk8O
pYlJFnsCwrsgIaZTKPzA6/jU4BF9LDP62mlVqx4yRuIrTHqgiqw6TP2ObfS5yj+F
mzHQlhZgSGChXjx9Wi8xwZc5atG60raYtZplL+2febtPWSH5Oc5qVpQhXHBVJiCk
Q6uYshf34o7FdEido92grDN2n2WHeSJbYqTnFV6nIRrPRs8gkkt9VNERgxcPZHx7
Dh0j18tkLZELuENLjQGoONdsqYxhWxO6+MQd+WPTTCw56ZFYtgYPoEygX0ODRUat
yaneCXkLp4O9/zvqloQquglM2cJswNPvdmRjNlfazt3wzoZVQHGXVNbcV6I9jT+Z
8o7QZ6GLLolNAdCR85omT3OvTMU/erA6//0bm9cAnsJFDC6nPRIqaqVIptWVrPte
vAsOlMKN1FFhD1Ef+0auFHc/Y2nv5wk2S+Ni12SckNbrPSBXtRnpTM/yicNfXTKJ
xm6rufqNZFnleGSU5FOQEx+uS78e36Fks211WEHPh5r+eJmu0tYS7prnS7pXZjcV
SHkJFME7NcDEmp1WUg7oVCbfJYa3CuYeu76X2U9+5GAT+QkIzEqyhOu10U5DQWwO
knCl1D3PDZ6DZq2VTjRi5u5GTPdLbQ4O8+O/D19bV19ZUS6PJMCCr+0i73zy0byM
4Rfcc7ujapW+XHfM4APwMAH1Wr7ocPWi5U5F6VbWAfTaWACYZhRv+XWdO6mlu5ff
rypQ2qvtfvKpMTfjYkYwTNqYSHHYyGETmWdabUxKKZv6FIq/kUU1IL+lU6OgLb/t
05no3FjKgUTiCvqsgGenIY4cUfiN9MuDe6yUhtxRtNqOBaalvBWbsB1mZa9ncxvN
TsjuKY+KThqx81AsZ/c7G373YWjgD+9LE+OiF3swtGSLhRE0uLXCZQG992HG1YC/
Jdfv1LUroho3jBKnUpQT9gLWA90vsYnI85SNsj81QfX6y+R3xNj3g8yHo9rfuYUv
VdP81ylshHIIafvc8KG5e/xa0Hh/SvEqztqy+r5nQHFFcSkvGJDVAUSfoFEoUdXM
WkDSPDrU1QQ9kZfVuLymvmDE6AGrUk/ozmepYsMgXNXshKgOyg2jUHytdWSpD9gO
RgSFWLLsjbYLFCFkKezkcBBHr5RzpcQEvvJhG9mKrArj0QQIaT12o24+/jcVR5S8
/L+S9t2n8sMVPMhtNaoLefB0uNJmNI/Jz0d0z6UQtow3Yx3WLaE4eRpCFYUFSn6X
n2SPXRa6HjjegaGJTCgGEzRLKoELN2eV6k78aT/lftdSI7PmIGKmrUEqLZ8KEp20
MGgjp0WEr7/hXwRixfFlNcpnODNY7Bzm8oxY/KZOsYaOyN1qWjUuok5XKK033gN/
24f0djn6YDOZk8zQG3UWWcFW3RdKZixYZ9yJbklklOSuicByJWQb8UfceUwl48l+
0Tyi4ix1HP+7F7f0druEJ9EVRf44gaUrd9Q6wqCAQMUtKEX+ci7UIaTwYNikqk4f
VTgsoP1v/Gy+VEbUPF0LUwl521ApVdjdNed1i8A+QpoQSiR8B1ZH+kviYmFm+sqU
AiPX1X/RkyBytUKSo3k61qX5Vz0z303gMHjkM/8twUWaLBqNX3lclI5r70sKtM7n
WvNhphNXG9Hdv8m4zk3NuAP7pouLfThPMIV5+uMM91nTnutDDyq7fbhNXRQ3F7Hn
fJ1nXU7Bvq/grteodFmKARgFFU87HBNcCzPE0iI7czEH9sNVLtp+eWCRm/o+Y3LA
XpmSa4mqoV/0y15jECSpatB8ACaS15JRS6rvxUuvM1ZufMegry+azrPM7A9Np3Ja
6AQfeDQUN5xhhoP070qhbjkRsDSPZGq3YeXYAUIOhK5hLNV/HxDeJtuWT4C39KUh
85AUv0smoMttuYFkxDc1dZ1qEVluUlAOzSEow+9IYj3XvZlX5bpxRqvGIHhM0QVt
LXNzNvDiIFw/xIfgE9oy1XcdJxAv4MObUwNZocNoWQEOIMAuPrZYGqWQL1Ay6Bxf
hqEiktvhAKNaP7QqMvzC3/TcKKJhwkNaczUsQAhvJUb5RqDBJrIv+yUP7H6IqcIu
+UIr8pBe51QT0uegqx+WPNv+xWc2oc4UlqjM1diSm9UFvVYHOYNTp1ChMPZwu5xA
wmyEaX4FqV/1uM/9r+7obRNvIsxBLCZ0S75uWnsMyByvwCjzDfbUKFxj6Cgd0gKx
Ylrrld281gbfarZbJt3CSBC1RSutjto3y6hTRSuA++7ZD+4/VgJhLe9ztpTS1Djw
+P1/FwPNvMPfNRSs/PcGFXQNsT0BkNOlP+Q3yGNwR4JzNdXKgfFLIGFGor0KPGXg
mz+xyD/q6EnLZ5gdekaxaDJqWG7B+ZHjdJ5Yf3+0nhR/5iif1GCPA1PNQ/aMB/BN
G8RBjjyAflXdRMfuGS1LxJ1PP7hqAv2ioPrQ7wG43JFFkG6cO6zILjypYtzVR/Rd
InTkXCYYjUW8CMJ7GkVLbLdMI3B88T9l/EtsWcq/WPW+bdyUrVRhLNyHaGAikU3g
YlGKSo4jXczyHECHXTxy4TUn5h24SfsQ48qlye8ISfbOGE91EqcvNYznm5wa4V9M
orJFINFh/fW/669X0NwHBaUf+hc9zihAuYNWU6Fl9r3glJ/87HGprrjRTRY6sy+Q
XUgsYTScCDN2X+4JTxDn14jNnJHoTBHVpmUdZTUMmKwYIBuiqr7tjr7LUW+EH6l5
JE447T+QxKQc/FOvWWw+t3X/MviSFguU2/t+feK1Si2/bTj3PseIPFp/Qxcrm+EY
6vvjAkGeNkA5co8b5DA5E/3jUEYlr5PCPpvkwZZ/RqwOxDEgZxr2jSe7Ryq0ZHSA
yniJfaM6xyR1ACgqbNyaIEjVnJg1vAU96mJrLm/auxlOYOtS0ib2REQ3xxeoG9LQ
MHzkABn2tmv0BwABJ95OgJWHddHsEXjxuFP0qA3e3v4SMuMJfMjLIlul5SXlGZID
8D0xNIOnLMG3aat/Ht46tQ95L8OfTOYf7EwwwtL7O6oVD5PUfh0wkEKRjbF8g/Ee
O271NMEGGjXriUS3V94lzeR3AH/JUFmVExOSQsbCWkRIiTDntFbUsXQf9WqzmdiL
irxslvATWTLoZIQcuL1KLbiwFIpCmHsbMZkOWwRAIQuim4+b0Gc9WctFShtX83/l
/at2i9non7N0zYVW5LN/VJPa3Wof1WXqNx103yYUtucFiD6auMbKoptfFnCLWZvW
otWYYm3e3jNAwoNR5WwE6ZoHXb66MEuHmMQ8RccSS6QYifMd7vKKT3EglAVrG0/B
dIBDjTb++0u7iJwAt2VRuNa+VEAunRMK+fBlG+b7umoaLiJgAUKrp/qpbV8ZbwSf
D+ApRtUBKPwbLfU8o7ALfUjyA+rC0gfbJiciYiwbZixqfvnPLFjSUgr5D1vpKIMN
v/qGl97WWwLkBUqCcWVOPV8UdaGLw6bEseJTKXbWJgt0MaOUJC6M7ugzMPsMEgcG
1UxS0Z/0sS2XoLlhKhan2xMOWOZ/J4ofhxgQO/u9bVWqnSs0xN1Ymn4eCtc0t9Qr
R82TtxmhAmgbm+nwVy6nUR9t7WBSn1SpkDJBhl0wrHLvFLklYUDT+IszTv5OpdMm
sO1SwW6heWVBUbKevqlTq+WCDrtC72NPf7qz8V6Lt+WVl5fFBdg9j6SqMBRkiMP3
HHhcz+lNR42YnROyvkN6Vo+m8mUvlAUI4SD6px7tP0XwyFee8o8y8rUXN2nZJGOv
38l5dMhbETPMmTY/I2YPI1zW8vWM0VQohLU/SXc1/oY9ttUsuap/HXa9DxLYdwAw
hKy/Rox2Es/ScsciH1HY+sjwl50DlrlAX+l816nyWX6uOhEVbtjP7BPZBCdR4NLQ
3J3I05mgQyygkrOaEcY2oBBOUK5GGIwdif0EoaeAt2jqrb4W3JPiI3AFa4hEpC3e
4L5hymPM9dEcW2XZKJcEcyqjxxJsRFxE4RvpFHG9mA2YqNvbN+REYRjwhd08jotY
CnFyNQXQtDLateN3pidauHMfqUL1r7HxTIp3z/Bp96NuWsL8OMRULt7HJW5X3g+6
XDMLjjbqhvnzu9nkELn63kASGke7jeDBP/YTsKJwcLh5BxZ83JOSpBGHGg1tMPyF
wsJa8ejfzE/XFRm2RjvsB9ZJQaJj3M0h2TiDjcOhnMcEacVgUgUI7V5TcNMMErq5
1Hs3SLswZHWhoMovsqcOOPqSLPL4F7mWoHBULD9/UOLPVaV7RbqKRxSM3Ng08G2s
9hjdfQ+IAsCe4bcGWCmBTcdrnPhZ8yZyISdNX3vpp8DDTDN/jJSrvjODuL+SXDxE
RGk7kM700eQGBeWdA1rcn5OkHTCDZDx7dCQ7zE/tSDRBE9AIVJW1i/Y2TfHpAKcJ
BM0XCQA2YJbt9jviD/BfisTu3DWx/Dx3COXHd9M8vEpfy1azB+eTyPDaShk93Rva
sGhV7dXWJrtvK0a1Q5PP/S8YedPqh4UPQNAvXzNAnEokqE+k1CIIRCfd37RoYBIK
PXoVoLsPnc/E5odou7mQ+4ur3/03IM2OcW4UDoYfh8dg3bfxHMvbIHjFFHDaugBN
gLOoOWWPVadHhzU2nnGTwI7ECBEBfFmF+SXdkJ4nRrr67Ts+aDJjPcOXeDGzCGoY
2KtrIOPGg87thOHo8xpJxivkkJOak9orb61zk/rdIrB5d0TRadrYyqCedmlaXm7X
z0qzfEZGQXlHkSNU+j30djKFle4oF33i2I+gOkLj72NYKT2K7QK0l8YAgCVtnb7H
vx+DNUdDjfO/ORd7IWKCFmeOg1Su3uN8CziJ4hOEyTsF8xzpNoQ+aq/pMNoYb8j5
QJsPVBSlZtdumav3wQPeaQ35US7xLIgeDcyhHQc7hb71aAbP+RY2IHG8scqxX6hW
DLz6ithXRnNEYcAi4ucR1M1hOXHeuMcGqs3HumWrcxGovIn+TWhzBeQBEmYtuHoh
4TlfFcS6Cw6/2lddqSXag4jtNbDMvcgg3zpvdvjK9LGMNZ7UiybqazWJpn3sDrG7
mft3qwsRsJ28n+fcRCvjzEuG4h9YjlZVLyDs0bXEe7/0VLe9W2bTs5O7JfD9HKXx
arJIRMiBWN0r8VvNY6yK1qaIn+LS4XE4XoAm6HmaJb/8VydXDDpleWvu6kdXurRM
07Hh4cJbXreKlJX+593gTgCJGG8NxyR1k1cCRA285mBwZr7ydB8VgF7ZH+rM4L8Y
WZU5Cdt4vVZd4njdRS0tiw+rxtV+FzIF2mwMhQfOC6LuE6vaCYI2kuKUVUjg7A/y
HFAPywc+/uW6rLRq/PYNSjViPwTff9ZFrEhCYzmQkuPGVyre9Fu3C0TUL76KPVE7
/3m/hg58ZsOtzQa7Xu2IPL3aat0KtFGDIE7g7oKtl9AnmM+jU6sawARO7c6nmytw
25m16OBjwnw+MCgOMKDpLQAYUXxMSq8tJOnYsQXnvkCzGdzEMaPCg+xtPjYFlPj3
Hq29S/AUKy87jegusCmQOpyA1D3yn+ym/uE8dPMN1pK8ZZhY1ER9AQeIRDFpMpta
a+GX1d1ZNnDhiQVo4jJgz7I/nmY/CpG7N5jk71Ap7eXpvihBKlDweL0yJrs76T+P
H7FPTECOiiEb8zbTF9PmGZ1VyiZwmhyfSA1uL1YmPUVP3rCk5tvfmxP1FxkXl30w
jkwZl49EQ8feSnNM368hVJSug8roVqfPUTPqx6hL6B0NZoNzSGpxH6qt3C9olaZ7
KOu/lmfJCwtGx2RttAGdyZ1/7wbCaC19jNOBnEygypDqhf7eiUBJHvKCHIzOmnFE
r14qHcHVQ9G79U7xxIWamP9plt1Gt8B/WoGN0JHXJn1VtXf1R6okpm7tXZv2v8wJ
7R364Pq4u/5ShB65J1bQxaEtMq5wKk8K7YKyh7o6ELZgPi5kBwfSGv8m6qfldQRU
7bECVjmp80jZ/aoaRpcIlN4BBta4D2ydF/olULz4Tio/aafhqT+yKuOIC1XMfgJm
JNu6iPGep171DrBPMYkBIWClnmQH2REKB067STSqOtZntXuLWvidy8qAUWbevUKj
rQ4oLyb+nWN9DLBQTKQ0OY7+enei2Al4IhNZXNFoPUJRSuclCZMcIeOEzE1jKr1w
I+WsMNHokVkRTY58LPvWr4srRRmT5ez2YLFGiJ4v8358B+knU0rNav4F/PV5Oqne
X0KJfTsi7H9bByZrkzZOhOZKC4+NHO0o5/9C+64oqFVBBln+iNr7kT9ZxRLCLHFB
0y8ndpowEaYerCMkQfFAGQU8KHTKzlrP42FOwKo2ST4gyOlK/wBL9NGTY69MJlA6
htaDuTSAJIhG4qsPDJkeRbK9Xkgp7Z7Na8STcVU61zKUD8QsXdnLh/CJ+sK90xpc
fSr+B0cTtHs9+VqIKTR6MOk8JaeYd5Z0gYuoaQGwrxlztEuJyjbHxtBsC55hDh/D
gf/zrmw2KD3WhJzqF5/DS3wSAJanbzxy4rMIQ86H7KJ3c16tps3dEykHB1uRRruK
XNhDDCq2mlmjfkouLTiNuLkIawNRoPqiV0gd2fA4y/PPRg2jvJzhnt6TZ/Abj75H
pm0BojFNt24mDKg+ewPFQIIKluMIBjFNg7m1cnvPKBdOhkStfm1OFT4cTAPe0veM
xTHqm11CL3463UZV1yymMP4bWd0wMngu6QqzzO3mCykWZ0Hniwxn6JCyuxUtPbMM
Yu69To0bRpdwr+p1IJ4WqIkP34Q/2Y+6h5Wsg13BcqrmqbsYKaKcvZuZurVzu/IP
HehIPBBHHP9FG6fONXLEFH2U3D2iGsstt05ct33ILWVhtVJxJlI4CCGXWNZay367
zWTtFJ54U1IQC0gN/2worn3U6MMC/1i6IuV4PwqIHI1Ygh4oPUq62BCm4Jiwb71c
nAKs8+ziqqfKyTou1rdMMBDmmAHui80aJZkYAFpic+ttQYWT11g3nHyBniEs5xqH
HbYwehs+VT2sFs4KRzpmmxqVS1rQZMpWMFflwXsxHRSnMt1r1jDBWYI6fe5Be5e0
bAPxeH5Q7bv6FYnevdqGqa08eWBSd4GrZ/oC8GtA4Vt6xKd37nzK8UvUUsM9yf8p
CLCuU9Z/mJtNRsEluclDi9qGLiwAJmmyqw8Oj/2HzjXOD3gWYnRQ2xKckDj+vEhf
4Uz0s3wPcIYm3pyeHKiPw57pwTQUmJiKGgm7UDCXZ8Q6Y79cZlflyN2SjscoB+CZ
mt9oxKzDSiL+r5uaa+FzJbJZMNeojYzCWejbkRiksTdJ+n5DHeI3o2PVifneHNIV
hozKMBjZoo87+6tIwYKGugGLK9L/KGuw7LmNHmtfV8i5eBQ7Ktgm3aJ5kZnp7SbO
7ulcobbjSnZzqzvkXST0gYQylAzP44Qmv9fr7aFiP+/yU/9aL1uS6quXLQ4KroX+
46bIFjMtadhy1znT2Ej2xXKyVfIRRgvCtZ2eGsqPAiOyVmwQ76QIXY5dXdRhsA/a
SARgheMEuj+C8vIc5wdR9VQ68MTUos4i5NkmAvnKIBajGndu6Zwo/O5vXJp3p5RD
6wJEjsw/70ZHbfKnvtW5hp/BAChq0j3ptvXWEp83wzrWoOTUqHs13jPqvdYe5yoa
N0xLCQ1qs2mZJ95tyRF9/Dt+NbXfNeZgFko97Udh7FTvU2SH/xHoY+qh/3pgzPTd
JJIqVXSWL8RVleuJdQQGb4BPFhDQpglE27plgD95zho5I2HlXBQ+RRbWwJOtgBbw
ZTkb6L0NX12ttGDgL1tQQa08ud/r0QZheaLVz3QlRsT6LaXqJ6wK5EySGzpDg9Kn
daTE+k1q0dGizJbvD3LZ9cqVNnyl/CLUFD/ETjC3nPOPsfhRluJHPlykD7PBGf/p
ZjajQiDeYkag8y+yEKjuHengMz7GCErjrMkKA1uiozYIv8K5YDDwoHTHES55Twst
VOqj7VRPBrTDM27xE5pEiGr0uwjbfd28MyKsULU5HyrgH81kiAMNvELg4WV85Myo
y57F4e+K3VLgHx/xomHHsX3nmNKLaNFcci4eZhKD9a/CiyATCNE0f/HtbAPY5eWA
RppmtmyI4+9IRd+/3EpNzkqVKN6uEelv0WdT0k0S7QaB47dcW/EiTbeL6Is0lynQ
P8NhhT99AIkeOEcl2Wj8v4AFV4WmWBmbPcnNPKbFmrvgaTuwHRUKj/yIdOjpmatu
OpILXXR4LeY2D2wncC0H/vnEaIdoMkxSh6o4BNId0/NllgZXvWw97heI3w4M0YRr
FxD9JO+iLmPXqPONS4BQqH4yhB7g2q1UmQPLIFcERivGndzFVJ9kcWRly8fiebsu
WQDPbj0L40xqOK8oT8Si4MUQ+5sk6mEv7nlwomTfn3mNai8RYr8PvXr5Rbe9vl0y
XsqeXLx0fFmvOGJMfo9KwkL0LejaSUK8e7hjx7aRsvdgWq3QQzn0ALz3LD2MC3r9
sbZoL8WdC7prRFX7+PIcBa7i9sqC543W+x1NKTwfln3AOMKJD+suWgbKaq7d3/k2
5I+6eOhKTai4Wcy7yQkydeHH9+/aogk+AK027zfsB5b/6X8yFHgojWzU2sxocqPb
FF+sdLPPq51uB3j0yaF4dcDTTpBbgy08DO1V0abUAhkeCKWEnyANNzAcPu2SswFB
qQXjHYnG+1Q7+3e3vCKBTL6D4RQPdFg7slNvyWZCbkJg34GgJtOLMRS0VzoJT+38
OTwInS1PIxkAfCqKEHhFcZNMqAELbYq29BlbxIIB+JEcqCzDEN9QqyDj39ays/Nn
qEY0Ub+S1gYRVkgiCtDNllFfi2S3h4dzDydT2OeAVboaWs7ozBaCH2DRrlfmhbFR
jbIAgGipTkM1PRq/+2fw7lklokoy74gOa41iD74h6w7Ep41sqaEd4Ffwum7Vi7GH
Pi+yRVllwlAedkd2OM8zV8yGmlo7jhWoMiVPYm3FsX4u8e/rZNg4+W95S8VAzzmw
Zryv5/2A5ZXOyGQDhaqr+0fm2QD4s8oVoqv5GJGB7l/bytPUXdUsi3qnT/CDdXeA
vl2yEztF6VSastG838puKzGA64R+E+hqo5AXt+aQui7Q5oIdZO9woT6IWwxcqI5X
Er2YtA8LQLfb8uX+uoK/99+iv06Sxpd3P/tiNCeSZ/CZz3aXVyUuffo783Ov2zWp
c9OitII/JArKJKoP2Sq6OtmUBbBez0fvdhnGo3ysv1R66YhOj4+pV5JGxGTJ/vfE
eNnkHnzinGq+wDMMecMJwIXKUmpNsA7pn+okWc5uyYo55M6gqHcGaHRZGjUO7vXp
2EVnab7blsy8zEdNmm2l3Xg6Z+mICpMNSKcK5vQlGJsBz7A1imCD17jTqS0eHFVG
Rcoi/AOAyfaifnI9YhX9hTC2dvSBWdMM4wPCpL3Efcn9I9bCFzcatxdViVcvyeQm
vxxliXO7mY1vvblOGHFN4tb54S6LtgTnQYdhnQ/U8fiySQiDI1nf1VrVZ/K5zgp+
9JevjI0naDMZUgROwK3DZhREAts5pMs/TIkUBwKRKANfL1MwM9qCMRpf9aQZ+6Ip
xrdROOsmV2B7lMNjbh2bQyX0LphTWDAJlAiFJZBNDyCf7RFGPdGyz80IzkxVg3i8
MML+31JkdLgqV2DEWwiRGM9Iiz9QZoKM7Adl3Y/8KmvBl5v/z2GH6ejdapJOtDXx
GfJSbXk5C3kp0Dbk0TFW0lzo8DeA1/9lqBU/QJZjMjuJ+cyZTAmoSjICeQN/nReB
mR7WK59XepIqTElbdOE7cSPRNqsqNn12o6jxnj7d5a9IU6DGhcami4ZDwbxhgeXh
wjC3wY6yBeSxFEOwQ3vhLDEnQv4kHZ+zRuWugraucxfkFzjr8dunAl6NmqRi/lgA
GcOIhar8cruarf21wx2vLEYw+0qeHYPRrH5vSFI4J4BPF4TWrTvgpCKIGU3vSe5/
a/1Uzm8kUmgnLPhW6Nyu9FFphsxNNcbJp/uqEgcP16Gl379OnTN/TRnSpVMSLKaa
6OHNp8CNrECDyP6/Yc8jyc1oSKfWUkU3WAEIS95L3XXwhUIUeorAX1CJS4iKKeX1
mo3FgyWLYSkkAKUEvYS4Vv2/nD+RLcXrQOER+QhHbHXjkeya2oGda44F7CMHpCaP
guMyZu/khh1R328Pk5CrJheH6RRoicCvibAETosT0ti6ylkVQ3R/6HxUM0dU+ekm
MQYO5AxFjk1rnXBFw3C9MjajjHt67Y0M27nxKT5PzqdKWkviX00lILfzhjN7qJah
YeympslzF+5O0Q/9N0VyHqKNP+Phk8tRYlV/V2GwcCaegwFDoHaPqPyTYoeoDqRp
iW91mXK3/+n6OfCqBTd7PtAZ0tAXJGs6IbAThfgPSJCSlba3Kid7m+GykyxjgLhM
VdIhq/ReYiELzFrEJQYmbV58OljYU5weLMWEYm3M+6AHFcYavNpZKGmcUY38964N
1wup6YSfOUKLNqGM7iFZW3+voE1EPyFRfNjj0CydhzGLkBnOCu/FW7U7NDfwJn0m
TYFVXtPaWPO1lg0kGOiQ2HtJU+1c3ilKzlyMPv81p0q1T0MZwy5TRuJfSAfNdAIm
GMhFA+P41d8PxEPIKiCNU8hoOJjUO1yO5L0uxCkw856hSiqg+lgO6Ywu3kMK9If8
RltZloUGh+zdcUn7ji8f+Q0B8XA0oryht1RFO4Wquqv/YcInycGHRB/C/hbxD3GJ
jrg8EfJhxKDlTj501LswqKCP7rizLPcB0DHzgEgyz5fr68iv0TsFVDsLplE0+/AK
5+vCUdAkQmSHj2E/nXjLXvo8Uf6/JVW2icjkYoY2M1lFSaWkVABP/S39oYSjYcUB
XQOI53oDDTMVcLRShQoZeYOhW+43VDy0YHWcWK/X2TbI7mkmEMW3SgJjyiqXlwxq
U4+uVu0xnuLLzIe6cjrTU20/U+BYNmNXrZMm+3g/VWab8y1sqF+5bOzgr+Mdrlou
Q0J97eKyD/e8sNewV5I/18hrmjylKos97rWc/a8t8h23F4rThwdKLdFbtXZN3//w
GAQBJsLAQQJQ+GDyAJID3A1cVvhpPCmAZQ3LF0rM6gHT4Vk3t86amevr/23FW2RQ
CISeKcZKKUrxmkSOAPXHYocP/qmQ1J4B+D3mlS8g7qjvYPZ/NRckUyhd7YYoeyVc
6jHnFv4D9F3BPTdkA2GKnq1r9uSU4rGv24iKqEE507fNGQzaFu8EehPUO8+dvigH
z8e9T/RfnwMXc/KW3u9i2LjkDqWnEVYTQbRevMagSc+imThQ/Z7uJ5ols19LXEC0
WUGVGMbKINinIIpzgvLdjeHM+VMErxPFk4AZWz29bY8Z8E5apV2sW34/+TvNlYLU
DG5zwNHg8uFDjxUBNp4Icfu+Zw8nMl2/PqBv8kd8K497GxtmQd40v0BLj9CuM39R
kldw9ACNsIyWv4kCamo94EiQOUOcJqsch1dXj7da3cBiYf/Rze8vF5peh0+ldlxl
UUE1fCtTbFAPQCvZ5Q4iG7Lf7iYu9Y+adO3ArBOzOmsKOQDVx69P5yr2YwfOE5Ww
2FlgF9Hyqb5q08OATPL18hKySHP1qc2zsR7hdSMr/jrZfoYcPohfFpnYkxDIhtIz
YbILJfv8IjmNpZ/bpi3KY1qKNe8/1S1ZrbIht9JNJa84nYp1EcaOrpIm3d1n5YEV
NL4u0nRX8YTyEYeDKmOjAQCUUCKU+nuy1VqAssNbdDqbaRDNgKun7TxCb+hZ+vRF
F/sWeU0r1qXnJF6TZ+7XcUJuIUG8PW+ZhrfqV/W2eFTL/jhAB2/EKxuQPNS/Hl0O
Nn5rHbUyDiEF1Ateaef/vMmt7GdNLg5I7ZS5Ap8wY2qJlYMedS9bEmpBJSrLzc9i
2Cg6Q0IE0G8UY2gvOsmbd+untleJ98Sm+XYN7ezIapUy+s7ChjAjGQqP0g8A9GzX
XURLoAfRzVYV+/iyA+Vu/MgqaOQXR0geUj59ciT8olcoDfsvQtbS/rr9wco6G4gC
zxWUWB40ZIO997oGtXIcOhad2k+6pl2vzQEFMn9DwH+M9MpEewOZJAem/gF+Nzcx
7RhccVZNAuHH9BEgIscO4VCnc0C1NPTDNu6daMqwpwc5uUTFVQ1fJpwtDBdyy8Hd
M4EWYv1FtBMb+2nhmGnTURNFY3jDFS2LU15aJeh6mq4PtCLdxG0x03n3CfSzxpQZ
SVOzsyp+tNN+0Ma7sW9HMA8wNXRltRY3gjE3o/LDFrAnHYVWDPTng5c9PMdkVZQb
VXoPzSGYCmJib5oGzYCe0WY0JtNxDMgJQktmZdHC0icuPayZds5ObyZo5DlxQ0Sf
lDWk/9bjCDVyc+qaYnAJqgL5FNOAAoZDAEf7T81FOvwAT5PyJH+qdVsE1Nh2jdwx
Amq4CEUVjIBi5C4rUMLhvyFJKOXHexNQ22rgzidBwB2S1PBGNQtCjZc4lZRtUHCX
xCx2soQKr0/AoM6KsFeH+3VCiisoqxT9UonzBn682z16XjsW0DIvoN8q472EuoYT
3Fc5epayLmtVnOmQJiTInSwSJBE3kPDK+NztXfoiBjv6yKO0Pcp7tjSsXtuokNXH
izM3RYyVAw4ckWkTygcYXH4ciRX6QeCHA3WNXnmNzVAPo43BzmiyV7whOiCtuxOY
lOv8bC1hvhZGWlwOUJ9N+UgCzTcyG2p9qY0iaOK+w8qhVDORy+o7g+B1g3/cHwo3
qgL2oldMnHxJc8Y3guc0tr6wPRpn2LqDGZD1PzrokjJKEqh0s8GOY7Gl5lwvrotr
K6EoX5un+YUtOgld8aIn5FZNgAVE7etkhs4BnKkZxrRSpylJOS6d1Ust8DapRzUQ
Bm+znnsNICfIAM7gScq4PQy2W7pL+WAnOFckmx2cVXUvGgZHp4E+u8kCo0ZBL1Ra
Dq8pfM9QPSWw+rFIzLxLb4rmgv4u/CYLB633+PnHFuv53je0gqLLrR+TIMk0jsN3
pd+6NK4RufuWKeywIUTd4p3alzc3rfOXwEH5pbxTB9Z34wnIFhWsOJdqiaqk7Wge
HHezR/l61n4WpbfnqAavQcN5UtgQGfjPb3aujbO/Ski4tNcbzfb09SWMljz5KojJ
DsHiVC0vdi0qnFTxt/1TTilYhSoNRhS86cyVI/q6UiEAKdf+FP1sn1uYpAhWvb9r
o4T4ZmZxKy6rYPuCDPQn10+SQ1CBcoE9QQ7uREE6+bgVCcDg/6rvxWIlWJVUBhD3
gBb1+1VRquzoQYY0DrVjsamo5ty24qKAxl0sHWOho0/iJwgLAmrzQ53J+eGfHBFw
tqDi6HTNnYsfjx0Oc20mdm83iei03R6fc0LxLHdPm2a8Bq/Tnap4jHxtcJpyryFV
vkxzev+GOkumrjXGq5KjS4/c91OJCu84lf73R9I316NtDEhMnEWNV33zZVizbweQ
l1uytOX8GaG3MKeb3KAJFOS84Ieoyqhkom7j9t4qE2CGQMESX69Hu99fCxa4Q0dK
vttbU12hHpI4Z24uJeHTD2DjPl1NUpAfYyxoO/CJ3ChfyXWBi7TiHU8F3I12711i
7f/fU8IXw7DHCIqMciRChzdXJvimuPWnjE6dRqXgPU7sdqtbux01MLp+ZsGFWZiz
wtQ37z0vmsSqZbbeALU1dtPtusEKfMYnWBf4OJbZU2aRv3dXTI4Jb9Sb2vE+si0B
ZZReWi/+ooT5V766NkYvDxG14hnCz1uAfXCzAXPo8iFUu9/Awgc8n5M6U8pVZa0v
SqHa8QFy313/rgJR8dABc7+ReJV6FvtLg1ZGcuLqQ69q4MP+gqaSHcAdjUjIbO/A
QMv7xl2ru2JnYjtQ+oY1Rs/vUUJALV/u5kYVzXiuqqf9XTrKRBPPkfZ/gX+94StD
1XJ76FrYxI2ITUefv078AWmDlyJzSlyUO/FW9paQ4W7PrhS8G1I25+K+4BWW9Ox5
43HmeCinlNzR77Zc+lIg6W1UC+JvPwKCMVMKVblZmPfiDv2NYU2XvRd/g9f4mLaV
KoaW6reyr2aokt3bzKLPzZG5jSfuSPbgZHnuuEJdd5GlK7zcP4TW6ezzYDmH/NO1
XOl1tpOPnJTabM2Oc+2b/4mEqmnzp/4h59HBBoLXphwTempWoTefe8DIxlgrK3D+
2f6ogfIqHLK4zx2ttlHjWRBh4G+Ahq5fsRSbA9fk26mIBRbL6PwveWH+FuG87ow5
vm5q4rauh7pA68IisSnSYl7sb4qVkGqhVgAmBrq88yMt7lLoqjJDveFcnqDZtf8W
nNfGIh5DPpEINpy54cEGIs2DvrbJKwaP3uqymPQu9XbWwKQ84xyPEFe/s48u17wA
DEzpdhFuisnXLPBFMgcQbp772vhF9u79KLSSFClSvl4QPM+cWG1hD+Snn5mjf2aZ
m7ArFnAciIzRUgsRJG/jmGhHGq97B88ID6EBrttxxn8O8UOwQt/GNOmvDRE10Hq1
Jtaq/Ehrv5Kzo1UnxGLcF/x0JRAcgZJtCdA1NXT5ErRqc0gLbXEVoj1kKFmtOzq8
I6/f8iniX3xS7pET1VC6umUmKFj4TmJSJJC8YQlP7Lj1d3PV/NGBYk9WdifavY3B
8l98BZuj8ZY3yPKywPzwWgZHER0w19/XJU2LmrmR+0h9CB9HYiHRe4Z7BwwGFt1L
chfy3u7O8xhjoGPUuV8fyZrqSHnJBQ6ohjQslrzoy6U8CrRxuNq6CMXiNqLfSGN1
f8irUHBNKzhKK6dDhLaK52hE2B0OHhdccd9GexnKuQrLP1n6tB30lw4uFnvOATVM
M7pEMRffkUt4MVGrjoUPUoh29Zdw31eAFpX/I8VcLKohtU9RdZIHkq1c8zYOQiu8
5gFjWyyWCxRmofAWwaTMc6b99eCPDsfjTbAWgvHqkywryAgY1GdS/9YNvluI/l3b
rXtbb0D3TNWnbOKU+sDNUGCYaRz7RJATSXEDbiQRjfWas6RkH2HRhN99LhQB7KBF
pc414Kx3Uv7HJSLdkvtX8wwVbHGigLTjsHvWJVf7BS2lrIe5WbryO/hXHv+FSfPZ
v/U6qN84y5WnughzaKxO8q9QW2iL1bVOeA6WPDeXADwNmYBLdxuzoJcuLAgeApLj
VEwsbAsE57QLkklUsHfH+zAhrm9nTiu5Um84rA9oVqzBKnjWpxBczocEip3Rmn5I
Ql/KZPLWBGgfMRJ9iocAUPY6suAp2gNF8qza5m1kEMJcl/KRC8gQJgat0s9psS4L
mLfLBHVPE3oL3diS1491QEMFmTpq6v/nY8B8UvJDi9aQo4zNY53pB39gcHI/Eie0
elthRirmBD1vY4RLT0WxcIiy7OqE+Z4qptjdoEmHEDVJBK9NjO1ZTIWjBHGAWK5e
9xQgAk8IkIXdsq6HAbo35TP/otN7JtOW36i+MgZW/GpC+10Tea356nIw31xmo8IJ
iEoL9KP06CGXzF1HdBKCLfdLkKpd7xtT1R0yGTbxosqd/ifRfO7SX+nslYvMtIMV
f+wZ8WE3ouvBwdC44mcTTfS8yNYBqltNZIxbVIf38cuC1VujjKZfua/7fJVReqNF
STHHuru6PtFuHpf6jrRhBx+TLxfJL7uxKJVoeh9mS71izGMbYZol3MB+BuE7tbUk
JKNy06cRcBAMLWO+uqxRFrUuXfsjreKa90il5KG4zOTX7j0HOsfxR6mlcdUHqDh4
lxa2B3NKMOfMo6L9dtIuDYoICzNBaqIBUI8tzkC8nE5PjujpPMGlFQk6RMdk3c/x
iCvIY0jpUh9Sa9i8ljZskOY1BKj9yRmliPgZBqnS4vPLBtbMVaqS/EtI2XrVVaVr
jAVD/FSBK22xDOTHUNuF06rBnqqWH/A/o1P4cB2GEZT58M6PCglAaXnJ9R2KABfW
Igxk6AGWSTbR0GdN3q9JHLpHCkpzD15Wn102qbvM/q0GbQIZpFNFlVkef+OIhsdg
rknli7ck51NJQGBqSk5FdhYQUMvl5W7VGdMxnL2M8fz1Hr4lDP0h0DebYlZ1XrMZ
+RNNytX2S5M05+Al8zb4S8Ni3i8gwAauBsacu3hyIb51vKOv+jO9TLaCn1RGpCY8
W6zr5E4hRr4VmR/1pMlDRyAF0mVqZlIYI5OyLlm1NAD2CUEma+DNkDkQqIns8ZCz
YpRrY/16RdwhvA7u3DlZXJdY0qHAViex8ZsqyYEanp8wqigx5NzB/wIzA31U9Wg1
rbiKj1+7Y33AEyjIFWaGFScp5uZcoisdRO1W137g8eiVpg2XqrF5uanV5GrWIs86
xOtj+fBi6LkTPsYjJQ22IKpd/vBf1b1D9JdCSJkoPRRgjJ3ZJEnmbEE/1dD9B6lj
e2F2AuaoRKzbQS3v6E7kEUUkMPVcppAfBo8YLc6sIpivec6NxgiPCLl9I6+091zb
UunYCVoK3OgJKCNVPPW6QUbR9qFx+rfidbl1s+MrmL2+q32vUIoW3Ske2fziDg1Q
SkHcB/lxsiKPuve1By5YyGUNVB504WH6H6bW9m+8bKUbFT1rT8ujN4UAER0n6v5D
46lvLMkizHzO/Zjx5cySO63lXOY/tEDevY5N1zQRtUlcM9CiwdPt9EV+dJ7FPJDo
4vU8iWtKmMDEky4FE9uHy32Yksh9151zZBwqss/UPNH11Qk1z5hRiiazfbueMTYf
J9nLVBvtVQmZhWus/EhvQnmzYbULGGtL8vFTGp9629n17+M0AF9neahO/iejjVrZ
HChDKHnk9epl1uAdhyzMpGvsrd5wCnV7IFImCH8yhBh49zQ/AZICSDB3cDzj7VZv
QCo7/dB0vAqQ/mikcHMzZgXBw10BhaAdMr24s5vd9IYXsUjzkZt6mok5A4FlVrk1
QGnw6YVxozeEHVjXHgN8JhUX9GLzFF2uUWaqjCnrojdXzJ7vuSckG6NvroEHPBMt
QUUstGK5SKM8Ya0Vhmf+91S0j81pQbZYkT4w0huWv6zCW2ASaoxLSwSdg+8PLHzR
PyiQwu6UIupr6L59HHbRoBCX5xyDMAZYDgP9leU6OamkETluAWzIG79MfhcQ4KJu
Iz4zsbEmDql5yAP5R0L2sXOzOw8So3jGPBoQdvCwyX5vmOIvZIMDmphaqTqGAg6r
cKK5Ki0iZFj/M+yHYoUUVRpDqC0bNt/33q2V1gnVvJdhl3NhhTqnYf4PmG8ct4SA
7p9dxIg3EzvBU+UhY7eowESwJPd0jjpBJnc5Kauewu70R1O1cxJtJawOUbtZ9e/w
BEy5bVs5OOXrPaIu9P4slfiG3TQY3Olzup0bOcb7ESg/230nIQlr/QiQ5xiVBAoq
MmIl5kjJOWrqRv16v/chFHR1C6fBUgD84ywXCsxxqo6dEqqLQ+86NzsiBrxZ+B9n
MmIfjjCQkxaWCfdJ4U1qYa0+5oShT9LDIE31m0pWHJsm7Z7ZbYwrda1eWnWdI9AJ
oqRdCFEliXlUF+JOGFs7ulpSPsTCb60NVR8CtboNVQx/+SIyLFhOzU8ZOEwBxrNH
dauKERRxP4fbDJ2dinAFsVtNDwJJZ73lECHSj81fbl1Edmn4SYfdNNu4Xo2R+k8h
h0cP9kVLgrItrtXhTfapwsevgXA4jiOcFby9re2nzqO8k367C/5D29abEWojw/55
iJZoPUu7DtzKSj6bC2w8fjcdV/HThHH2wQCF+oMJQ8a3gCFjHpBc7CghHCTQq5dW
4vOpPUtLOR0CEeqo0O0X94wOu+FlAm4nuwFgA0VTNtaXnj3HSoK0T/Ny9qdA2jcG
IPA9iskpIVvNMIekctFNvOZAbcnoy2tWKYiwxM0r9ec8z7FasIvlO7SzIwZ81VtN
A6qH9tTbSG8/1/bVETCD5J+4mAz0bMNloOXDg0rqn8xK8EmDi0cdW1VpSxVorxnr
ABt8GeMA32iJu2r4uPz7J0BjnsQWRLUmhU46502mQLsoePgRpRzMYE5WdsJIhSLq
nS+7z212tc8cFMO2pY+8Gnoe6k9x8J26XSmhNuGodNmAFpDGFAQ2p6hNhF8183qx
BuMJS9dY2y06+SERzT3XZNP+/figEk44c0ckMspvdDUYmdGiFRdpaegFIrNxJGEQ
9JS0ERyNAqCav3RwTgH6CKV0O3GfHJ2snObMPfujwr0pgWtyfqDn7KhvCJxuxmTu
gUoVVBopXWdwMl61ZISQS5uy1p68XR9akH7GEGTVsA5bzVt4o6KTiQdWXHAEzC03
ywrXz1idJU6VdkWT34yHl9Bd6znRJWEXl7T9MMc1APTOxqZey9or8vPNyvtjNEFI
zpi4cm+g4mtj8ayCdlXFJGAiALXsVTBkJxNCgDfIZmm95tmvOkvUO0j8C/XwWRmQ
zRrJLibpQWMXhLOW+NQctUUKXgxaPN/fUir6KN9Vv1Wps3QqA2JeowRriqxafJoB
Y/CiIhGZSotaMKZfmjb+Y1K4sd/p6OX4qMsUl3WnEonQqZIEtZelCQW2ImBlwza+
W1kpJhVxt90h9drnhVxC2RNucXTZfXZC3LPg5GWYgyKnyLWHbbQU+47Bu2cfkzn1
ms0L2ihQDBYgFx8bLFWrivAlXkxTJlh+BH2zenIIKvs9Ozgk61Vd4K28ISNPLV78
sqPaayIH/zFBplzuJCj+ETcHDftmWwZNXbHCz90+COvP/pDjIidk4m9AnEUH3a0N
1kJgBRKDTJAyZ/JfiFbv2e/IonFRwkXMiAQ/6DmOHzSH1fFHuvUDOCV4b/X7FfB0
zzggJYjjSbvZFn6HcrJCVycrhbjldUrnLdUrsrIQPEB3ha+5qYU81DqiZwD5GsXn
bOfBanuIGGtNrOSQ+KUVfn7Dh8BD2Y3N1VCq3UScHZX98gT0fH6L3KeVBwcDLPxc
x0O7SrmbWGhgrG7iypIT4yCJVeTny3FVNhuqoEAjQVCCf5EGsvJXSPRSyEaS8Wc3
xxEgAG0nmWzNjBHBCb+Nup1Hx/S2CE7whbUe2EF0zp4V/P0KEiuss4MR/JNr6gWB
73rk2zgnLZjvvDAR+lR7rpYRyhcywdP2BVHnFZZkKfwf4QAs3+xlFgjPb02JDElO
S0Hjy5/ckp7cN04RwMPJXVhxEPTwRZ4tQKSgvAfgQbVmjqnuCMwytA6MrmJWZ90Q
a3PjXPvxzo6gfLunwliaogGg+AX55z/zdapgL1tQYlfVuVR9fy0u18wmi7BRnwX8
I+ua8/TKMSlphQtjkyAtuOYjJgiIfuQdU4sdK64A2fxEaxnEVIFiQA1ix5hvKUKx
857XCwmVCTIHUdXKe0P4Q1fwycJq9rs4LA4OwMBmhw5d6AIHtDwESoNYIsTcdr9o
YZAiqW2NAn+BgduDDFmEuPIv4VzuSlN+DHA0Mk0cN32uxH9VNL1+D9XomgSmgRNN
dzqf3EoEahSmX400yFOUDpNSzm5PnSfF0bMlI2sTwin0RGZyaQsVEMgyxt0z7lht
fLNUPqaNX29Q7nqlq/ldS/15EypPf7L6UlRoQqEvX8MjXp1XucBReL/t7tV/w/MX
6QS2ou0/GFIDay9xVJVub6I09mnBuVClnEaLTNFpPi1ZcU8vMD9J55DkEctXKDHo
ZNE2byLdIV3ggglahguK+REWtYaxvJ+wPyeNdrPN7vLYeEDLFBPgNhxPzZGqpevF
p+XxLdmODR4p3agfTwZEsWeGWmorKDJxqL9GSK737BzpzZqjxyP9gjfqmm4OV9T1
ysOcu60rHAvD2ShguQnRyK7OKFzB+xN4WNgXQLwqAYlnYzw8uhP5nffv1jtT+e8E
vk78j5RVsQk9BmI4D3lMMP2tnJ5DGfrS4eVibkasWe8avgWCNMl+M5kmew5MCfCd
qds4Ui8AsjoMgio1SwimdwqPaYdxi2QJ9nih96mSdvLvnNQ4vuwqQY77wYIc5BsA
qNx19EqI9Zo+B/c53h5gaQNLZdAhahe2Hi0bdF1rplKAH/QijZENvv+WNYcaA2ip
Ii4/+RcZoXvTxboDdVHI6CSjlDvl7nxRo8IJS1i9evdExkuLXlDT3uastH4sBNoe
CmvwyX85/Py7t05JSe2Npb2Odgrdhh6kq2JXJ5Jnk0tZYGWr39QIvSj4VchvdTrn
sFaf/YAmD23jQ9gUQJ/o6n5ARwTdYWWpDZO6Ki5FRaj65fQYtzCVF0lFhR1bxZJp
crEPk8ONWiae/0Vfx1mywOGQwtFwv+qsENSs2CiCq0W8MT0ywqgzrlvTF1kQGpEa
Osiz4PXDXZxVIbt/6XmGKbBIuXPCNkSATKPK5lz5zVkXxcmz9r6C2pb/8N/WLsSh
7wHt/0o6cJHeNYTHpL31TIMslNrtSJI5bGuONak08t1J3dwXTaa3onXLeHnKSTuF
L3GnjET04CFSezyR3Bl3sP6NHh4euC3OougKO7n3PXYDSeXdsw5y30UCadYCNGNv
slkhosENLs1/Ou95zZd6ReCnydfP3pIjoSbFKaklkCdaT0fNeB537G8LGYgrvK0R
UkwAOIJSz6xRuBYfiokwwZLq6FhDB7hA7RXMqGxoa6TVuar7cGhiEqF2Sjtd5EU9
T48VVQ4RvmLW728V2uthLp4k5v69ZV51rmB0Ag9NS57kg938j1VtWKeTn7ISfPba
sDh3LEvadtgI9D9UwpcNw0KPRcbpC/X+I+/MLdn8OwaYUcMse1YaeqYTG+C80Y0v
INudVqSwYzvmkv05CRZjWRGk71KPpmDYVbT/4FRVVLA2gPLkN4Xe8OhfsEHa2SMI
nfzixeyYkVvwUPXwjitBFSyA7Im2MaSND8FIcM+DDIOYNb0RN263Qk6eyH36fVom
9yITcZOqTUcANrcIXrQhEMfkoTYdGy2t6+Ymmxe9qUr8q1QZuN6gIwGgKLtKSdib
5ku6do02skdw2i+qOjTReWM1QQKCL6JITydlGKyZQMFi/wbMiUdYvcN+ZsjF1eMy
xK8u+3cmzC43A2EXGMtg3ptXs4Hz/C1lnNzOJzhfeh8Hz16+MDnEvVfNXCrHj4gJ
JvO7kBfRO+3U2rpBKr7PBd9KTrGkWfEUsDu7Y+mT8zyOF9uH6TuPPWyrs7hTDBPD
BZE2jtRyrinaXBHSHkVs78Ndri3PCg72+yNqlKaZVU4zL02VP+iP1err5zEoBwy+
YTVMHIb4mRDo576x8c9dGXm13GM+S5UWoLYm87bBpKlUzH/NUMQ+3LvdmT+8AkSa
8JCedJKa2J1Fvpse+5TFMEZIZAShV1WJ/bldkZqx+kb9VionO8XHviyMd7rb0DE7
GwlcNzq5Uj3aeLmmSpToqPQQov3K2y/yr4Z465gOY0tgj9XHYeuS2Ktg9+0pVQH+
3AmhmimjsYXFqFGcXToeO2wyMIdA/fxbVxF8qEaZ+LTGbAh/SY32qs5QTTOX67Cv
G8rokNtVIZswWAu5NP+9LqeDMOqZiRZQC5YnKzoaj8Xk7esJ23rOvtQfE18afhH5
AfBKyeo+E3yMyaGxzTsKqVtWaUT2BjVo3lwbMGXUt07P7+pg28z4Gw920+0LgAGe
Ky9C7bo51nXTKY9CErsDE+8qJ9y65VrlUH7cs4P45nqPdOSXWUrfbYgHfye/cTwl
rik28/pTIBKuHClF/SKR0OSyVLmCyjiTGoXMWYMuvP5m/7f2bHENTejqMqcxOll2
Zhp9WDXeSKkyQVUSQg0CFdz5TrTRk3kSTp/6/xpdERvKR4cqYS2/pslaEBDx7bv0
v5aGfJRYdI0R2zgbQYOkyOoEIJx2yp9dMpKy3wpUZ0Ojo6G9cD+KxErlQfTYmv2q
DwCJ/QsovyvE0Ky9XPM5NOUsFMr3u5jJmDIZ+/qsmtO6lsLyO8xepxZL+V26GBev
ptYX4p/igu1RNZKeIHevKEJQ9SqSaGwE8mWFXPRRgQocWcy2bEMRKu/6wcvScgPs
yQU1J41RzBKGNxIEezg6Bh54i383RPaJJrHgb4kfpFEMddDg7cko11oRpIm98pGO
PtpgilsVNqhncd+VMzYA6Nu9PNlR70SxumebwquYT043Vp8ATodhqSdCqygkJqu3
FXmwm2do9LQp6mYLLOB7lXFq4jlu4OpBpLGXkVKkoT4/7ZKsvJntpGcSRxMMDvPh
m1RiH+DguP52LxXVSJsq4NG1xX0XLVYeNLmrWgCHbyqCfausrc5uvLCs/3+67ifS
b7vaFuvzQ4YpVlNLa7BKyPv2hnjF+y4qT6iVcwlJdpzGgp1SjpIE1fehJA4NawG5
rMlAaylkis6AHOfFOLfpR2tA2nz8BAvJI8E3HoqMfK0aCXHHi3BOJf5YGP882+bi
n6cvEoeqDAO+kcj5XTqifdP+OQ3PmrUQoMmSknLpnFROW/foB6kdtLWT/jyYv3MU
UqrUVMoHPj7PCVes+sn+DAhaWLE8TtJrP+plCUuBM5/jyBrZmkOjaa3iwIH2rERl
38DrLe0omTMFG9f3sg0fht0VnNpExM/bNL57Kmsa/2L1VYKB4usbzmzL8IHMiH8k
p1tQSsgjPc4ZTfFShA3ntadqXx8npvgiQKQt16OhlfmE6j/MVG54zmya0o/l0CfF
kWSc3l6j7jXpsHQKNtpokTEiAA6RGj55UcXG1Tx+JCQJ+F6A3Dy7DPcUgnC0oKXU
qOgXW59KUdlSD9kFDzYDFA057dZQUx6TXQ/I/VVbrNwaSJ0n0pD5KcVTvqnWEdvt
KXMCnBHCu52+JYrBdljgiXwVrl700JkggglmRTsv0MXMBJkyEcOiOOn9X3CFoeCq
gFabR0eOIvkZD5o2PRxG0YWSAR+Nfei2IQTuwQ96oBf5jGXyerYElt3EEp3G+xaw
0O7Qr20Yeq+GOzY7RXlFxuv1q89Nkhf75DCSPwKWAHP5noXwIf+ymUlF6/CPGYVB
jMSQlW6OvhWM1AlnIuThjwW6tcW2LikvCRL51LWHFBNx994HX/jYgbwUsvDIM/vI
k6oVYSRPiE62z5WOyKKJ3TXnU26Nv5+UqJWsW0tJgMmP7UHX/WTQiQBPMF5Y0DGJ
NtwfSeQFRUkDEEmTfM5MMHl+SijQMl+7JGCR/eUBKLiNcwcIBkoCbPAO0STLY3oK
sdfX50hS8vJsK+pnIUBN0L8CdZz6TRfNc1DxMGS2motKunOClU0bSpvytmOCT0fI
giozCIn62R9PIsZelibblyX4j/9YbvEcZpl5EEKrVS2F706slXelivXVAwv5qSgD
Rmfj6VgDOCddhlpG9kS7VJhjRSwJ6RcWpZVETN5V8XmGPGiidf9BrypNF176kyT+
JsDZpd3lIYNNa99Vs+G3lmbzKbtcnIeM3uWRP/LMAfOSJcw5pn4NmwPEQViebYwf
mOGK/HaJhu+g1zLj+DV7VI3dUzFtKJ4B8r0wGFcmqWAFFmAzzpkMaKKmVVh2Sory
eqJ+Zf/H/PS6Ll5vGAW9/ScA40JiDMI4LMyBCAqQoctj7IcFJ694S/yCy62jpR8m
OvU01oyeXgQSH2+XsdMNq6KiTHNBGd4NpyAe76JZfnGSHp01mOFsll0xiGtzfVOs
xj+w10MyYyucSsW6vXtBfSpciplX73p9AuwRzMNd4/G8L4r02tDmdOVkuGfwa8Nn
TiW/SxwIlvoRSh0gT475K/xMt5820ivGt30voR7lCqfnlj0jvSP+orXU9t1efLyV
2/tjULaQJpPIlPqUPdnr0PUNkGVfjPqW6H4TJ/KCP35sdeaKEOwS3Zxi3bfkN24+
8bUZcIAe57E4N9mf5HlCGIHTL+crrQ1rcth6hQZBQyMxIOqwYog6S7qcDcQ6NoI4
xn4vHxMmRL1KC0PFS/pvu2TscLp74DRx1OHY3ute+nDMitoa8YmLdVWHO9n1vr4B
AVz5v2TI+vZsZJYCNlfrWCfBhvMwsLpqAiXsaPtbcwGK1DT7nMouO9ODr1nX84+7
sMK6CLsb7Amy9H0V2mTsZQmPCtJpHAKdRuqrfB1dxpjQueMX35vcixC97TIMPBSL
iu2ClRywR+e2erPnIZnq4+uZ6yza70KauIdas5cTeUUmNiuJOcCJUJo3i149XCoA
BM+XrEPylvfmPT9Mw0OMgTwk8+sy7LTnQtY3mo/Kd96FCQfSTi/+KKJ+tdevewjb
iTeER2ph0rNIz323urH1Zi3vYrpzDNe7r30DQECfA6Voaw5qcuUWFwZ+F2qw9B6B
W91w9ygWie1FGeAED7Dz6QCoO2DD3Uc1XwkXj7vN/7c25ShWfBBuUpE6ld/MxxuC
+iKfgl3khlO8XT6uZJ6xx6zD70l8vygqZ2pZP8aMDDVJwZ7xjA4o2ozrcufBusDG
q20lSk+E9aMdirFFCYFK97er+khs2aaptmWYAO2elApF2k9Ke1hOg1u6vCTX85b5
vsLhQa8YsJUYdE7bRWvYinJkEGBNUu51ooFRg4NnQUA1gt0qFWMzQumQWIzcHDFr
LXtKfA9Ki1bKjRRpKfHZqRptOp+BywXJzLXwrv8Rc+muWDqqyDPM8jMuSZ/+aXYQ
rvvs0H4MeVj2gjYGXA0TuGlXTLvLNi20PlzCl92ChtYfvf4zTLaX3/1FBofhsiwK
AZgMwUYeGiShglo/vchD/oXWHVg7VO0WOaH3DN+HITyC0jOcnfn4ti3uWBC8f0+W
SocGi0fc1MMfymeiSFl/1XMgscr2qOdV9/1aVibZhkaNtooYjW3hvrJM0bUx/eWe
thkIee2Y7KsjxQzF8Cjgji5UH/OjyHpmeJhMjj6yqdT3sbfV3IpejS5aht3Faezz
EFp3lh9TTC68mqctG+SSU78I/gaMWwDZvcZbQ158f5MgGn0RAtW2StyIutoKx9w6
EcKj/vFwEakVuUOvNj4Nui4vaSz8zgbCTj7nIjkF7ms1khXt+NedO7FQVJaFi5ey
59LvT8MHEHuD4f2dbTAruy2eMF532rgrPI9VKO8Y1w/PdiPQB8lLqlspdFPD7T2e
RaaZ6ErWCVAzU+Z1KAd1Wt9BpDY2dDq5fXihwueuhd1jfak9WWH+vv8bHREqPzhS
jhnvZYS9Ui95g20A9TXInG0VTVq/7Yx0pEn5A+McRTy6dDisi0znay9MQPmmdb+G
ZFwM0PhJk5wU9D7abHTvupsGxml5VgNG3jvddXFwjpR3+rNNjABlNolO9jWuDml/
t7o3VmUW4aEdUwmIdXBaGTgJufhMXutoDeyWg0OA0CmmOw3Pl/FZe0ymrV/ttTjr
wOwfyAnM8IhbVF3bBqXmugDmrjMHaw+0FQwe4bhzH71O7hsOd5lt0WpIggBPGAD/
Q0N6lpGzgvMQRDOKz2uEUm8eUkEcE8+quyuRqseb6eHijLbyJMXrf0aBNc75i/HP
fWmOgy1G+ZHJ0nDH8cz7xs+MWcJ9PaNduWJz1vqyV88gE0/wtHw32uNfx1u+NMKg
2GChRwix6yT5ORbUxtfgihbzABQM+owJXeZO4GjnPjullqeQxx5YN7N1u7KV5v3K
peBhgkNX7f/FkFvTRvyN/Iwr9AIsVb8Bm/CKlDJkEquQ/z5IVDIhHzvsoIrckieB
eEKlZKH/H5SOlBSBuANXA/vsX4ldYJnu7A3gG7k69ZT2C5Y+IoF2cBd3kRTd9wG7
8y1uQ/kjVU56DrA6dws/LAc5CScoEZK2JE1/cPae8/vA+4xyyKVItuB1MQfo3DWM
y4R64tj7xzW+6FerZxxT5SyfxoReFOwhyNhWcWcF/AEU4j8yCBuVEQnyUBnJrdZa
HG4NHnFMio4pxDaK0VmYrrHrUvhNCmlTDEwzsaAmgr7wa5XY1j1m2iXRYq9/y6LO
0/SZTc4mO2jp6mytWH+XTPGmCq9+tFlF8irVtg/wl6HhfNIXxJZeFJ7aSWQVd+nM
MW92QNz1CehA31R2r8wlhHjWE9AqUgyEulr4sq1HyMgL+2A5xxmZgwe8bCdPC8dT
hb1Ri6UNowhqXe8NpnOmzxDVjY4+ylHbzrFPnUMlWdFaIPo+JlTkVQuhbVLwksMD
Y+ytLJX772NmOLHBQFzpmW8rPKmAorjZkOyqftXpNf4MI/ps5zg4gbCSdZ2WNHIX
TM5ZIAlr2NFnPzZNP9fljRvFWiG/JIJzhr39sfqGex1RHSju9EVpDZRzSAFoJ6I4
QuGtQ5oETHWGAFcJuj6Dayl1cGlxmYjSZ6tqhkMeNIE0DoO0UjxFT4jRQPxG0siM
IIE2XsV+FMHVf1v2Ize66QTuCt4eztFjhLvci+PVZ0OtY/eVI391yeOFh1pXY91R
l6vaedrf1DdEdInI/IpZyufnNcOJwg85BBPwzJvVnKV1mIfz21I+OV7Q4GJOZ39S
VSQxbyv0hFy1HThIxThE3cH+1ykRe4WWmgqn3PDTar+UXx05der6YdoK/wLbXWbM
9dwetQ7H4TxSAFjcNoztaKZUXdXaLvgazaFU3eOqMMvNochGRDX9kXXua0fhsbLv
9k2FU1Bq6qBcD8rB6vZqY8kbP+XzwvkEoQRsU8wUqV1RMuh8UDx9x/sXkwolIdOU
Mgpy5mnovodgqSsUpNf/pUFMp2lkTl24sST/gVsJsy4tPA/uSNsEQQXajFETTEtx
8tLv3PGKz3n25fT3jq9tqFRRG1mBYSFtinPeg8OVWE54Kv/uNxxNujhouHiBR61a
qSld5oWFfAAft3DAoZGxOqyo3m5ZoNVCV+P0JrZgsmh3dY9DSQB2L/HuZFDE+V/o
YJJhDoVG6Yw8xmwpZt/gFbP8lagUiYEv3bPkNS8g3fUOgArX9sDboUEGhGbEeQwo
xTrgTA3yCbPLfj8b93m6PDeABvtY9T48lSqqKL85xqqLtHFkfI/SeJesCcDsxPFD
llA1Du7BdkWwsO/mm22+6ok97+o9gJIBfFhf2/OmUnyooMtRzC+VfkKVtLm38Rpu
7PdsUpKC+MVw40zCulRccCSVisRRB9jJBrYoFMHyujIwzv9T0onD9ermNRp2vwSB
+NN4XUKkvSAzDHQgiWHmjOtuHAJdvzdJCSOh/4WoclXPLYKWbot3KKRiCSiJL/HR
H2vxcxGL8UPgmtWoxXmJ/nfo2w4XfplykY+Xi+Xs3qKXl+emhjR+3XPGygfSjxV5
wIVtpGyd7sax4gS0tU5rSg0VQ4iHrpa09jvsdlUUPCUhE8BjZF6JE/Lv7yUEn2MN
FZp0aLK5uR5OL1EcT91/ZnFdu5F0AdaCYhyB8RoJ2FhAShSA2zqXc9HCxhFO6p5v
zIQPdZ1KuLQjHV3xHPw2xm2kn3zJE2T3TED7eEFJKSP7arHmxj9UHwKEInco2v1p
XIG94YKLNgoG5ePei1c0RhKs9vk6tK95xYLdfUO3h+vqpVOWccVenorLZ2aOOHQT
Zno8gcsrKibywqeCO3LDOk9rvve28XyXiSJislBOwAnd7CP4sk7knCdMjJ50E+AA
k7UE4KM6dTXB0P8rKP7Lo18jLySLEr2MlaAI5QXw4+NGCIx4KMVSblknUqA82V2B
e//OHHZJgtEwAd/XuOEqahMUIzJ+Ox3Vp+mnTtGAIkfLvGW9/W5hjCYiiqLvUWWd
B9mkqHyw4AvfcvUh3M4iNfafJ06Xt15ieWK/05TbvNgh1VUXvU9oCLZIQOhLyYDe
EKSBBUHZY+FmxcghlwhBuKE1gi9Q1P6xJT+BTMMTXKNXUqvkWMViainKJBwEtoPR
muktHrR1ls5IrZKn579M5BxsJY382ur2QFi/9fyGJp/Xo/TyxN1uqp1gEfLUn8zN
E5MA8DS3vE8+EMzfsUkLibKrpdykKy3CeiP/3yOk1ZXeXYyYcKqNCbNASpzUzklX
giUgVTGediv4JbcFX2I8YY1lWCkys664eqxZ49DlKdAybwYEdeSeqsa3pdTT2PIQ
LAcw2rA1urjEo9DKO1urcp1AZttcCN42LoQrhvXdBNoJym/69OQspVouMiXhotcH
jBvqv+A8IVFG2m6Wnhxe1Ok4MMIVv6Csw917C7SQemsb1hsymkP8cJLTPGlq0ycM
hVbJlEF2X0DpJl2/v9TJDqSapnK3rcy9rL+ZN4Gf8dwX/Nh4eW5mE3mRWqbVVRWs
GUF7v93CQtsKZ66Yy0FIzWJXj2q0kxwYDj1Qr1q/STo8zbJZpdFf3yJM+6WzNm/5
9t/p4ztFl22BceBSP95HaGA8mjj2QLZ9dQ0vwSIjURnJ85KmOenkNywW8uOdMOFs
Te1jQHNQKRtwTqelWXxZCwqFcGB4x1Nnev7dWIfW9NsLmslPmAroEL4s9YCHMuep
k1nr8LtGRp+SZcQHNWnANCSEGdXk0jhfd3dE2jC74ElUVAhVBrd3+2jdPOTuMD7r
754Xqi0rbsYNlBBzfWDILq1CoZvZ3RzgZf/ku6ebdiHhEgEXa2gJnr21qSD7qHSy
9ceoRk/Kj1xyAUT+O1O7OTRMveFR2KKGS/kIigLCYcWXbB3SKTq0FH4kezyR4j3B
GdDL19tN5n9hnvrAeAJRzY7XZ0/8CqjHFNufNfYdDWKzdzCCJK64GsWTTS3lMUPn
qNxVAD9zzeyA1/vvSvkVDVN0ADfQH+WEg4EElcFji23tGBbGVhX4B3CTzy+k3QY4
YjsbhfYlkDaIHcGVhKEelLTdNn5wtIGe605UCg3EJ70C9aRupJIJFzkNpHDMMJwu
3T9Rw4LwmFi5WuREMHbUrPQxvgnpFaMwk+wy1/z8yR+jLBCHphhgjkJF3e0FIsNr
Y91ybMKX4qY1utSPOwiJDwEI3/5nbNP+0axXGFTB6O+OUakIORRXbwgK+ldizF2h
QVfr1i+XddJoPXZJoseKjML8JDw1wX9Ro634g/7Ix0rjYDpbeIOL7DbHVjsifAsh
HpKjgsT1wU2eZ0hrbkXg3YkNceAcrMAnnXGVQGakgLqgmqoapq3aS67Snu2IgGTw
QbHSi8Zo3HsT2D/byWQe1cmV0+2cjI0b9216hkzraiyCzAuBPz0QXmnFJly2rP6d
qdiW1q6s302DLLWyMJMaI3QSshJoyexaAKp/+cICeETdORfgEywvfX7s9dbutSM3
0c64kCrLP6+x3Vcnu7v7RXns2tWeecMRlKpdY5z9pnLXLyVgCvD7CnTu0Zxz09dt
JxL7j3frcmkpn+qv/WkbM+GEAceNVD+nA8GdoPnMTqDftvgtvpZTUvbTl1ByiPC7
37RnxhvUqTfEQzneXj05bRzpF4Kxmx50GBwEqLYCriJG+x+p4AgclMR8xg65U6XX
8d6j2KascRyYgFLvNaskpMogPaVFM316k8RYHzIabI1tgEiztsC/HwParSLLQh1Z
An2gYbRFhqVY9RGQd0kJ/9cx2vb9953LI0qxGa1NBC9ipjS61HyyVM8Hu2isX3Fu
79WHARbVz6i+dgZNYfkBPzt9K/zYyA4i6Z0KJ6ksyYklCHPwtIBjQJnBivZxJw4a
u375RI6v4KBlv8Q4Qet4HVLRwtUgVPogoO0alxF7OrFt1M/CfltLlxMsRqWxSGgc
YUTBuUNFI6grh3U49xYSDhcIFuU/xlb746E/Cod+XZ+/l/9XrqjmQDMKZOxqHmqp
HQb3Z4M2/fxyt1vD7raRqan9/NM441X6OyBov7ni2rbhyMY3NctccKXSnKPcUMze
qToq8WkmA3w7IPaBLYzGK4KVv7/tGgCKh6hGAsiGmchaE8/dq+wSWGD9QZ664ivv
eDMjmceMV0/ckqM88wRXa0QVpGpk7tfUz7bl/sDMlTlBhDKewrSwYOEZjPcs/CCs
RWV4QHuUWUN7wwNSlk+U1q0Q9x2s4EwGJGNsYvhFxOYLBRP98Z6CQfwk0Qd/EoW2
4T7d4S+46qoNDSMnL7hKUlIUFnWz7lSaeLH31VskPAy0PB1Y+wy7yH6z4XOloFtD
Riknmbu9S7ZulSv0v8zcOyO+SsCPkgkfi0fHBrILYgxutcaoAySucTGcVLk/Eych
PdPYf3YMYWoUo8FbQJSsBvbM4HRZ7z592XgmXF9MY00F6dhNy3KM+smZ7Ya/abTJ
vQGPFq4DtlpE2EHilO2A64p+m6AOLRnKRUKPTidiuajZfbZ5S5n8I5gNhIoo55kj
rZYnLeBrfP558LqErYBGhk2iLlQqBgmWPcWRfWYIbtq/YeDtGWm/E1Ub5f/DE1Nh
zmrRDpZeYjkljj4Kcfwf8QMrt/hAg9nPYP9iJj/AMAA51ECDXt6LYjf4Zy5Z6jbZ
pMt9enhSfLd3WNUrSjnAkoKn2vMLTrVuEOQIWdLwPbu6n/1oYYUcKb/Kg+SCsiWk
m2Xtsp3Ei/01OH+DkEhUrWRm35VRMr/MTdf4YVo1Lh19qwR93YpvfZCnIZpCMv8S
G0W7bO97L8WL+2pAu3phpoGwu7YgAok5m1avJh/I4OXkPhftTT7bbI6w3d7XV350
10HMPQKgY1dClxuS+PbDcxx4ce0UjcuVdOYwAMjvcWhwQdQrSSoXukbpT3tTOgLv
/UyHPChiH8QXJde6jQ2q8Wb+H6GVcmXW1FF8s6zu1gYrOYWEx937FV/OJlZ8bpsJ
dSMyPjW4MU3prRKBVzlAiKabEIz9T5MC6bs8K4TZ+DwNlCLopvCRkP14GoXUFgUv
mWXmPeyfbXdi145YGnbVWaDUcIV4JHgvMRZTH2pv0A5mNGNaiA0oPSnS0Zd3VrUh
2HBjR1UHEDn33Bk7DfjEtVHl7Va7ODoBJ6H8/LeMwwRZcqbK2xgMNg+vVtYjjjkn
lwXAC2tYXSzFOm84RZuD9pWaccGoPZdYtLQTuJplhRKgrQfm5K/KipZPBtWFy6Tn
3zRVfgVSl5yLmg8YjCK4VZ1YkU2udqGLH22OAGomxcu1cbWyvo+meCDOpASRqTWa
xpwHRiUUW0iFRKjR3vftKiVbovaKLm0OlC19CrtJlvsRbQMISvBip62zRQ8gO4MQ
S1k5SASFBsvs4mEuxVHTAmEiDbF4Ifg4hQdHdxJ2szRQtsgg9i8AQNevf7QJ2pQ5
a+WsLFzXjawWzKVkeu0XA1UkXJp1reNN0NxoqyRtOmFo1sHSDiGFBMxVgE7E/pm9
Jvst5QmH5JTJdydgWnyaL9VhnJttr2Bn1qd/tnxYLKTYIbkJEAM8IZo88JI7KM8O
p/jKDaYUHdEXlMkYq6iJL8LheZN2sJ/1NHRIVJr/63GkzioYFDqOMsYd4vkor3kp
7H+439wzf3M4T6rMn56QHlvjCoTo8zEj/urVPIt6mxYsnd9kihtDVSuAMe+GHJ3+
MtZvXYlNKv/fuQAJ54Yre7BJhL+J8MxZNA1MllAZB5VNW9IM7U6VsbOF0+EhQpJ4
JPW72u7HlacJ29iFtejeI7YtRVmaTl6aQ6C8doQ4Uys7cOJE/2UVoY0xeBrN/4z7
Qf5Wvuv633TcSvxMvOOuwifdNmsNPrCIGUzo+vSO5ZnI/UxyCJu1npEpwWwOvIWg
JZAkgZnjqS9O+k3J0iO48VZLZJ43dHpszQY53Jjdde3nRkYEGqT+b/OcksFksETo
SUarxTYiUcSVGtfXpUAHOkSEntS1hoR3LqPdTYN1ayOadqMuEdRQO0j4q6MNisLB
kQUgus0Ro1OSaPsSF6D6RN5e+5ZDdQ9qIP4Q2lAcQ7wn8bbLVeHL6QE69blkXlhP
h9pgn47b4qKOOq5NykP6uYszulzxhGdbkqY4hK5uD8p5CWnpDQht5TOatYo+bEE9
o0OepGBs6anChyw9+NDKoooq6+iXvg7kfr7aAwiyvQAEuE2Z+sL96DFo6xHD48IY
0y5v0ZLaAulWAfzprzZ0ITWmVy4cYEMeU7TC3spmoUsG6h6NeQj045zzgvv1RGA+
XqPeRlfyGmOeOMK+g/UGJfRpyeSzpQayPh0blN5jpD4q1hinF6TVZK2Ut8t6Au76
86dh7kFWve5xMzoh4w22PZRSIeQIUGhe4mKuvgRu1Ri2RRnC7Ane+OfnYn3CwjcN
VMNqUR96P1k+PKJjohz6w+XnB1gqXR0yxaWIAMl7FuVrfYQnZqfOgAiREahLl0/M
OszRpw/mU/c+5L+vIjLFEzxTS6PxxHXBBP/BBlEbavEQBf/fF/WSEYTshp5Yp2Eg
EpfFMrg4nhuQ3XCPVjWf5BwRXVWhzczLhcZU+Adbej5usTalil5do7LMNpCHZl/y
vMUv09ZDnhfHFfEZO01gsU57M44GoobQWxqBLwZTgoExY6ME4Gf+bPTGX/5oM0Lv
+JoDb22XwxPU7LdQuowGrKgnXBKh3kjipBt5mebuaCvcE2v90itHBpgriSxltzVq
eza3+0KpRSJOHNwEec07gZJCSIcIT1yzPCHS/Tr+t3BblzV9I6GANYFnFSMeDk82
AX7mnYPd3vSxWoD6TkNf9UOSBpvyrERJkJt6hMyQEZj9W+GtU5+TceBfHuvJXwVS
0BFvLoU+YOVzD8LstpTgFMClojynlGmcR3B395HgvlCBDFBwlDLjZ6Ms0/9D02ge
xANgxM1HPYZM2yl9M9d8ksaU5V41lQo0PGAcD38c2JOAoPua13hxPx6LpV2DvZU5
wL4i8Tjmv73VMYMgih1pZx5ARe4lqE1oo0SsNCkUezX1sdHnkIgU08QYetVoeErN
lsJSeGK8o4ROtjWKNpiQiArjFDqr3h85yr571ZpM8w99rPdYd7GNVd/K3FpY+IOV
N/qPVC0MypM4Ao7F9KOYkEOPQWvpddVS1vUnJs++sR23TTvciUPi99zIm51W4NBU
ya4epGvo2ux7Z9ZfErMTxd+kCNNT2ncutz5oY3zMqAIJW68zPU2sDcvFjLcG80HW
/dmPCdn+18CBRT03QlXibpdmsv3wzTvjj5MsuBUDM5MUZsjXoMc+nUfGQ4LIaY40
fygYGcF2FGJxjgFe1lT56c7jgd22bCB/t8Uf3YMW0doL963cJB6ztCDg6S73MXCT
ta0Pl4e863h96i8rU42cAYsbRtc554Hvxfrkv/Ji/+3BGZKkSBJ4eRdUGlefX0PH
RtVHCmRtieYUJk1eIk2sM3SrxknqEyL/DZ6hs9adhOUKGmyxdwkXeENJw4b1a3jf
LnTVQ7YtjvlWs+57byXMehIQruw3pBdfGJo0STJ7rIQZTLU0Xy1KZ+qHYhIRxfiY
l51CkeADXEl5D+/wqlrGMLGCGuMuyUuupBzoisFLaqxQVLZR8Cy/0ZcIBUMNMbm3
WpXtVxg4DdFWSlktjQ4xdzXHDDuApdfQHmKeTnijVUHeNOBJSbVjpISslw8jEPhf
36N7BdtGdB6UiFMuqyMRuk974vSvWsM2pKzrL0/gEp/1FDAOfXc8JZYi+3F31UCY
4Jfln7NZ9j9WLh/h1JAmfNKH2HuhjFweG2f3snozk+QAEGXtkdnUmMavekk4NcSF
a/SpBTFosFpqtNrajvCcfZLJXqDDrB62tlQnGrJfc2iP3kBMKcrseBf+6wT/hKDZ
QiJmJK56Rc78FCOY1lCoWbXVrGazYicrY2kEeRyaG1Bm1uhxGS3UtTcwHd5I6VgT
byRH/b+pFXWQn5pMM9Py9bvc5rcWluPZhoimRCtQP2ulhSDK9etFrGCU1Nyai7LZ
gTp9iuR7wQ3AqZYe9svrv3EyJmHyxqWncDCslVB+4JwCEkBmTYC2Qu/hJ74Q0gw8
14KRmPBfjwPvrIVJzYXfc8+jrrcB0KLU0nkMVqII2mGDGFWsfwk3Bg9DuBQMXOE5
lAdyjY/g9u+Si7JqRliK79SLHvKuDX/cb4DdObDrkK7pfp0d5R/O0fn7vjmI1aHg
Gh2ghrb74l16+ssLerC49+PLd5VqeXtOyaBI5zwWCR5/a4pCI/iKBQfLy1C+H31X
r70EGCu58ybI1guhmJAamoJxMsDu3dmltbwVDrcl3AKqtxWquQEWgjLlzJRL43pE
hgZ4rrVbsAclK1qaaxk+LXtd+dArnxZ12+pti03FLqM866XibUIeOapt0SJq3nkX
04a7kQZjfxkpLMPSphlIEsclooivVI52bm2EN+jPRl4JrN7aJ9lYSqq6toowFoGP
Q+ccfruP6Kq5NM1puSYtD+Q/vOpy3mx/2Ar34FVT+4YruIbGSfxee7cUWroJZP3x
dSWe7aoHi+NrmU2hlTeJReT0jSTo1+myYAcNcgKazKdblFuCEHbDMwbP13h6jPwG
/I80feBvwM72u7hsgdUMEF8H0/OUtzY22u1GKHslIntNDWWvW96W2QkCTlP6DHgK
Q7jZYFe4K6zYaubeg4LHHF+N+FYSFo3YRVri9NZhe7blJXWqIkJ5f28igvt1gkOP
7Jc3vECE48UA3Jlch7KXLIqRMGXwcKz9VIbFbq2phSM8SrzK01GssA5ZJZzglXpM
IUtgL4wxQaHxTqLYMS6hgaigKpX8OX1Lpk6rwz5DeIGE4bUiEnQFif+gw8uymClY
ukG7aU6Uw7CSYqofn/aE1bOpGO63c4qFRqz6CVV5JulX/PbT/Jv3PWZqfB8UfIEy
TAgOit2xGgjaK83zGFAgDhNJlbdxaJpeyyq1W56ympecVKZK6FETwUqIL1ctHi4O
mW2eDqrI/fX2nPA+CCZLu9FP2HQYvKNbwrLrEJ7cNzb0XdKpbwLaezK2ZLNRjds5
WtDjBhjGqJjSsrokUJdhTWVPr2s1YlZuRZy7mJIt/gAic3DIB+GpqV9qjocor6XH
XjkWYPTuMAIgrQ1XefSQPrhCd0cJKQDfV2Mu71zOfa2bREFQzpevR4AmWo2aeKZq
2X6dpFHYHc27SMAOrcxfY75AAFOOGptQzXiYZTKZpzoMRzH/6TZHvgwJ5X9AsLIt
n7buJCCIJoy7WNXrxxk5qaOwycqwl9K7AmgTiv8zCsVAGkZDpXsYap52GAg5q/Kb
/sV0+snshJxehaN7gpHRqYJY3EEb1jEJ0Ke/NaU6fXQNmfn/j4pBa8XzMvMMgpLv
4v/RdZ9Pd/Np46qZAAMSvSI6mGPejodaHKj25dGm2AW3n2FaAPI+YMuwYk0vacJK
d5iw62Y1ZEFywiKaqxK4u6Ewq2SV+w38Hlx/FD611Jw9wFzSTwaptjXJoAQ40Lvk
eFTs07JkYjCDIJA3xYpSr+5cPmDJ0/XWKrQHm+Y6ra9dsUc9ZYgQycg4ulVeRXg+
EHFIsTJZQIQadpRYYXMLlC0CDDeAovi1rlM4E8G6oseShx+g1/SUwdfd6WskaGMe
JHszRbQe4RSwc4ZTf2IRALH7AakwhtEEhPs/NhPujvBLYua2eGSNjkaWPLeaa0ZE
uDFM8a5Qq4b6dcKt1UkDix2d9MGTrNE/bh8L9NtokILfbogKOFIWqr4WjPDC6KnL
rbGgllI7sQVn9S1YIiel1SC2VgcstO+WOnDHu0HBPXiAhA+Ca/jCbzEEMVuWJ2co
ztCUtZa/llct/ZpcYY/6Hjl24zEGxmhNU3OUs0B5nK4v7ObIQSeIbJ+FyCZgxpC0
VU4ZlCymHe2zWpeoFOicOBECMmQ+y2bW4dPc9dFnmbRIFnsZssA4Iyw2Fa6Zz7kp
BJlZiMwmEgLyCAOo/9xPjktmlY2RTHbezczmwhU88JjRqMXqtLstkUpdJHL5Buz+
kQZ5zhoLpQiC1LOV5CqknPU8FuZ7At19AtbmKzkXoGyJmjkVEtYbI8wnoK4wooHk
9GHonxD0p6mqAd3cOGXdcJ+ooWA+1WiN15XmXO8TXp6MIeSfHNZWYTvzrBs75J1v
wYg3SyfSqRNR+4kBRG5BIQQvK1SfkIW8ps3Ae9BR2bMERV7p7lMm9NYq8U0KjPUW
8BtDGSDQw4sxWm6pg31JUfTPZLrPDUvY9Hv9Q+ixMsLwWyp5o0J5RfWh1+UpmZHt
V5u+FZaP6PGfZsHLesbW73gJm/M/z3+4i6a5Tfj7TFb3VPwsXmJn5XX+/jPZRBE8
MPXc8Qs8ptrkcg0QfYy7hE2nBHrrYcdCvuJXrdwyFvqSw0+ctBW/fbGggyPLFcnB
hnLVfsYF5tM0On3HxGaYbIjMmODbANtOZFBNjYVTTrDSNMJXAkoEb/lqZOuANcua
C/VHkmS2lFlEFUfbZjoGJ+4//T+gelaZGJk+l+JFXfrBzGsaKXqjWS/wc9xVt2GG
LlwfEwbYlniVfWU5ATCJJs9mIepoOv2bLyaK+n/kNRPN2D3FwT0yYRMcAuZq28MT
bLE3Gt+LK/jFPhlKoIM3mXunBTKnsriNizNAG/S307wA+9Xhj+B1SkKZEQU+chNp
MfLb8d5yQBQH3o4nFwmjuCIxSujTg/LPIkzk43DIEzZivvBg2CtDp15wrPJYV6FO
eIfpMMJbL9Nkw6MtBVVlwC72UQV84WTTDM57PIX67SU858PNdQsJnJtZCeLT3Y/S
YpzJJz+gkm/v6WgCbZXBNciTM5HyZxysgg6YUImN6kiJNgpxd8FyndNHhybLgAll
STaFNArveSb9u1DWyKFDZoIH8TF1zsj1Hj3mhqTLFXU12r9UipgU5ODbvPPG/kWC
eV3Uv8XpejPt+x+BGRVFNT9Ajo7AjMH5m71rrB58dHmcZ8km6ebJHclIqgjU3fXq
aa1By6aSQ9em/kW+8eLueV19Ty/+7nwIOKv4fPwhopqXZBvlLkCbPIgEwknmu6v+
IdqbQWhg1gyzcbFpSD9nLmfQImDxI8fXVR8eyAIAdMQCZNks4OUnebOsbVtDXEF3
1Go0WVnjKL521yijTM29ptx808ZHb+hxtPjb8v1VF1IScYZNm7jSmooOQlOEXcLu
mYfhwew1D8+Ed+Q8MRaAM1kkFP8qXT05zPGFiWOK/H75+eGFs3pgATF4kjVhOoWE
wXfUAkWd0LQQlnP8RXUJ6+0KkrbZoGnzhrjqpVitR3jgBC/hxr1oUNrIVdIqZgUk
4gcy7V8WahG5zyvRFNChvvKsTK+LHc6O5TTBqoBwO3dPDUrA27YnardqqrdIByA9
1QpvOMjCni3kfbTMcCwqpg+kouuXQj6br9A2rrcco0uhepTnlJA6Asj40TsAXjUN
JMZ4+81DdDGbAgQGdXtpyT4F7vLFv01NBuY+ueEDEiw+IGzCuysr1TK91Ry9D3KM
7ue8Ktj7fubxWC6N3Qs1PymNT2tI9c6gpaC9juMD9OZkmu4oxVJbySED9jtNiAfu
dAoSnSaHxc/aYHsujdhX3bQ9+NZlPain3RG5XJNRH5j2f0IjK+uF15NhpuNh7HwR
PV5ObV10y7osz88wcvtv4UP45QguMMTWm2FuWQMj1tA3C2pSTFGHDJPA3OnRVjIq
QDuSENE7E6RGA1X7n5sYfoUsIwwoiXQwLTI3ej86tEVCy1yBSVCfyFMIlHekYZqD
mBVarRacc/21oMcok2nnJBK0ifW8UHV1idHA1e2UJb5s74GpjDG3kwXIUEQWb0yo
iz6E3jPxVkfIkDhiTebpDNhV5+3qE2Y5xVzZXRFtKZYm0fSsxFiQmmlq9QrIKHdD
x24SM4wbPI5FosaGKgd7pGwQrayzDW2YlGUA7A4qftuSodWoXZcRmFNj9vdRsH/X
tYgYjkEStlDttJAAx0NbJ2xj+4MPSdp9ZF44iobn0N55XQeMcdc75j0bWWR1KKRr
fT05+Z3l+psd67Ali9zFtruZ+S8dyQbmw3VQqwx0ZZhNn5I6fOu2A1LFfFAUQrxN
1/4z3t7RlKx6ukhJpcioQc1E9DMqQXgVNnH7z0i+2jKYmTySfY+vcaPxxwrx8C5G
ZdgbW0TOu2kX5ZAg7mZdP3W4HyqjUIj1Qg8XIg677azhFlM3ptTL5YPYEvQ2zq+G
75pTLR/46DMhfOflIKKWqL5lvVWbq5BiSo5Wir2tdz15EE+7v0J91GKoke0Qg9Ky
ZrpOGsKXHjkbLvbUOmQCDlHpHEUwciD6Et9RXMzuMl4yKzPxHo5XojiaOecuuGY0
SecJkAeMOFy35HnwkN15r/uDTnFgXlsvVPDvcVJGawSTGAGNDgR9qRhYCK9PoIEr
LnWHjAw9PVVmd7vMmUzltc5Icz4zcK+5SngJpau73C7q9qnr/3Omzf/d8VX5/DE+
iST/eS4yMDIz/iJlU/3z+NO4ej5CiXtk/+M/29d9lhPBuLtatKwYPlF36QElYD4b
49mGBTtGjJXzDk7Sjj0xNSk6vciHKQGExPMfrmvUQtDwKvEoesmE+ahllnB8EIVx
WuHrAJMK3akr9D5e8wj/dK9k9j1ppEiUzygkOwRAf/f8kMnZd6meAI3BJ1sneYo9
2ln7OZLMuR5DsFJ1alhavAyS51RGD544iRnws4u6tUD+o5YeaCBprYQ2QM4salAo
AhAjMydFeFzpqCI7d9FFMYBjh6STHoopHwOqocFQ+BcwXzGoyLAZXKc6IQVIABzX
x03rG5Apmq5cCFlhS6Z7TFbKhBacca7OXKRtU3vBbtkVkB06usttY7qT9NoSfela
lHBU+JltFvIRWBkiSo7SGuVPl8BNbE9jHSHkUg6iQVdwZddoO2I8cwGo7ZjW0ohN
7ImopwDQUObMcGyXoc8wwG8a0EUDr4PDtucVN55k8d+rNWOFj3XHunIF1axlpZK1
BR4jLLmyonaPzKxWl/bBfJkdsckUNtbLShGQR5qPlqK0kBiK409YzaCxgYWJB5pM
U6vccl+QHC9tM/OFPEdR9tSo/0H4PSMMIUwWMHLJMZCS+cjoIMrHjNrPUWRjrUc0
ozhU9M5FubHAvm2V0xxNrMPIQus32gsGbRtPS3CksWpemtv2sRS5geDvpTJTt2+b
xoVfKHdgVYyzOAr3Lsh80Ay1IH69jY2LGFjzdZR4orD7aoWuGoukYF3tuZUGn1xt
pr6XOuLl2pLmtefL23vEsuAN//8Hl+NgsA9gJLQuSZvc/dOKYTaPmt02g49Im2rV
7VNrV5mNMwg+w9aJFP0h7dC45tVRv/tiG7wORtxYSfiN1N22OrxJB7K7L1OnrCdT
RqIXTr0uiPXDR2U/VtZirjeYI4RgQ19hmG5nuZ+V3dK3d3dfodc3IfcJ1NdvNRgR
Fmt/4skhN4h4jX1LpiI6RrQDsXRd8CW8iZG3RPU+YLkQ8U5Oaw61nBFlffW6hStS
YwSW9cgBpDcrGyJERJ+wITb5qvPRZNJgc/Gmvvv0oMz5Zx/HKOaYCVl4uJ0KO5hf
0tRBIc1Q5dgSDZPOu1pX+PKKJ8tWIUOmdpzoUBkur2rSIC9vWjAHklskmSAGYXbf
hPvsE29D5ZbL4zvoDKfGcPoGBGn0Lyarp4y8KfozHPqd8SCXo8fFVf0aI/nzjvBJ
Dw0CI5yq2KR24B+PKR3ZtBQGkBNQ4WAHLfnv0damDK5WSQ74XmSNrCjnPao0bewX
n06GbqSr4kU4pIlHa0HtVwHUIUgMi+v1wQr2NiBC6H51x8zSmYxOolwvdnuaCLeh
YoWBT9bXrsRPkzQYg3Xb/oswe71WpcWFjOKiQ210Z6VqoADyBOvJvA7fs5b6SUOq
O91YJZzKyUJ7isHZwn8SuPbqaXX2yU2l6E4jmLWTRsK42vE9wFftaXZplb7WPQlL
QsihH4X3G6xHX4+w1/vuxwOqtdjZQfKp8DBz2hz3x5tpKuvNqwiuTlM3khgJcXsM
qY5A+c2KdCXeaF5N5cDzTfxSzaAhUa5Z/NTELXc774rS8FScsHWjeiZpg/OhnRh4
wpvlSHoxc51v00i0k8q2NtdknjH6X2FtGlNYlNR2s0oX3VHb2pgbHlCLfr+Sqo03
Xi6fTT+HVVqxWHr+HEPtci6duezw2jNH331BMiFWnvi2T5/1eoe9hQSklJw844VN
ok5SoTe5y2luEwdIQ16yjW0jBSEXeYIC7+/f5a5ADbHYzPZ3eefTAtzCABa20LoA
m4sE5vJz/J5h7Y1oeeTfiYqNHmMeYcZan3UC0rryGZSltW1Z3kPnTunlUjkGNoT5
zin1pDKx23Ab0KmLLyulOH/8dObGdTDG9NRl8EaSjUIN5D9fFCwC9/gJK+j8yvYe
/m5kVBbBrJHGXneupJ41PmXbnI1DHhQUgKXnJxIe677Mnxaaqw0+r9pCXepAO7IR
CrNGfSpq/iNFgwNmE3LsSdbO4hEgchMgJUTWnTkx/cxyVzPHLtH9rkjIBQxLex0O
bgZSM7Dre3Vzx3kKEZ/X0Iw6hHCbgbIl51GcFya/A4eN18ab+ARiMLRyPrExTgxu
4dWuMnQGllsYwcXLiTiDuyKGRljtrGMdpc3Ar/jIqIm71+1jrrYWh7AR/WIVa1Dc
xREw5XUgkI+2YB7Tr0svs8lvQ9SkeVuKDVmfvrP+rv98HMvcI9gx5Co1NcPA/t5n
tVz5ADEdvLKT4sdtYY7B6n04wHZDJ7nIyW9qioIBKAwBroZtKKAqd9ZYK65seS3O
3VrkzKLvOOMJqNFB/Y41ewUSowUxxEB5GUT+vOhWguKOEWQbysC6CJJYXhPnF0ID
AK0+k3ok3EUKrnheWmBvnWZH5/wbMN3Bu89iucdxXz7qWjHkIwjYyCsToZaY5F76
ePh2vSB6zTSlJ6M+QUbd6TN0A4nUL2WULDkGiJLWRqk+Ib2hT5IWgOf+cK8PKdW0
J6EMD0EGisDpd3uGT7yB5p+dIJX6d7VUIou6AGY0Kg6EttH6SLnZ9wC6krtGzwNb
SKroLFjAggF0uurquEH8koQkZOeNVGOZ+Rh/YBU2wCCsp8AQCbCRies4dUjXY6jT
ITt8a9g9u9orHDhgWTWFLIIwhq3S63YRdQLN6+4i9H7HfsoppaPFVDKCBsSbcTlV
qntzcu2OoxMx1RMPisA3J8Qk8GwOppZjhjRVCoIIWG69S2jRcrbx6JZJYhpHikJ3
D1gfF9ks8ZBcTEp//5Cfz7OMBLQpysN8sPMfxXqbV5Y6KkgwTaQeN7+qFUe5Fs+v
VafWFu43LBnr0jWlRPmnfVqgd7x/g+WpmYEDvjROf++VLztnnDEhAfXiMzwTL9Wl
n8ytL9PiB0F+0cz7vbZhpl5WQNWlH3RvmK0tObCTsbR7nFpRdBTggVuLVImzccMe
AODToVow97TVxU+F+wcGYeIHjnIPVU5WAyPsXepZPuruCYaiMyh6qjhEQGqRBmo/
IidZkUIDLqi8Eu//8cCb0LKqnfzpbAzIqZwodSKeGdrfaAHMXz0VGsBPjaTVlWoL
zHxZ7S5JzxcZ1WXzUahTJI/jcfctrrfd/kO6Die9GMVm2iM9/6OhmIdJkmH4XazI
3hjhF4QKdfZBMDo/6/e96hVjNHp+zozsBeRYh0TMLcabfcCTHxpza1ZeKZLJe5ru
6aAKiLbyLcCixmNdNdw17dX4LlNp/RJG5ZWHZkKzdUc+sM6IDOQYx1ls5bq/Dhmi
NeJNVF/XHWjOvjT8q712yBEdYi45p9hrPW3AMBrp1mSE+DKEk0ZkYnuMQLhnGV4f
7xHEVhWuSb/4mBl+RMWonj1+geZddSwrRyNLWwh6u9siSm+KWe64dVZnM7U/9LCA
Q5qOWbrWCS+5L0wp2H3rjpaXuwdRtD35KJ/UdLCILLnXWY9/k/yyVyQbymiocCRE
NwAqAV3nT799rdZ6VlS6/AEdkFlHvJ483iPiGBVIir9rjBUrfDfZDUtm+AD+gfvf
e6PufJ4wDJSMndfMoa4/m1Wv/BKMfSnqLlhSu9+QgSVRHZdWItgj8wBvhztrsTfb
NweiKv3IgnzYu/jepQTkXelN/jQdlIt8oaSo1H/+ZmDOlDkAOtX25qQcqGaN210U
YvvJte/xiUWIG5/4qCBhwLvLBTfb+yLaudZw03OfB+B+14iWD5lEFclWdSJuF1tu
nAnE0j/lNG4HH1KpEx3VXzrbZzv5anSlM/oedGSOjfBCC0Spbv4L4EqffqmoXXXA
Hl+1VQUXy3L43Bju9ofoaII2FV+vtrEecqYPCOdrwdBemWLncnqwSn6VYPQkKIQv
RzUcCIepmDb1jq5yggfXMhpam3z0hKl4Fu4NDjSqdsD7poduaAiHxTFdDuilfGNg
tczq1gj6VCiwapJN9tr/dqro+zLykM1ExsAvENKJRAmfVM2zZJ+hHf/UmmeUdEjb
aJu7W/D1j2EBf/HHGcCwH2+nap9tY8a7KsKDpXckrH8dDyAm8SaRQC+iVVaUxZ+F
SHaIferTaCZ3OgUtzgfxmlE+qZZPCyTP/f/K6reeWDl1gcnHlh3c/cLRyDiclbJU
MDrp39zqJoPnKF56u3zi29i3XSjPZCZyqgyFQrK+0i3aZvGke7K7d7fJqIX3c5B/
Ukt2jp4be7hJBc/WbQTnSKniymeSieaZ1hj7UGUc+BtfU0JsN1lI+MdxHH+RfHke
NBeAkAZtmSOBe4wTJXcXBKFSd2vm620krfAsQwAcov2qHKI/A4icimPFOnbAnr+1
3kBM9Vg2ifZEzxtkBzAQLtoPA2KQtlkhOnmZ9vggHzg/tDFc2YrCFM782wJiWGfC
uJMCHW9i5G/no3dU/6/lCf5mDbdwyHTOuJgeAt1BFho9VzSxQ/F9T2lEqLl31EAd
5LFD58GQY8Gtke43nixg4G1khR3vOzCvVmSgUUiF/nEckt0FFSIJVAkO3Kk6RE2q
lpU9oebwOPNuoxcq9LPkqlERva7DfYZoFH2BMomvoGxBEfxDrrRKu7uoexMDqBDJ
4m3XCFHZoDhR4QNcqFfNn65fEvPOQLbW3td5BNeeTaoKPJfF+Q4nwJOBqmUbbbiV
CqU6YyT3/5Fi0Ncq6AI8llkdLSEezPkaJP5F9qWLB5EefUn1u5zMyimyPVGMNjYH
34+hHD5391U0kS/bNMkpq33YoHMEjX1R2iKnwiLFvC/G//IDo1wOnCXvPnEI0wnB
t4vOoWOhvOOM7ZEP867OVfxz2Q6m3MLJSm4iwMkT354TnpyAnUNMoIVDQDw4bG1M
f2X6IgkKwqTam0Cs6js3S/2TZ25Ef9kYBSVE/I/bOMiZ08F4ay7dZpuYpaEwnG5X
HjqqHJhyFesn6vzwldiseToMEwothCnrGOC7b4Gg5NYzryVdI0YtnBN7yBFP96F5
unhO2XRLf0b0/Iokyh/x2i5zThl3nv5MfrneChzDxRtcvzDCoWB0QBZoN8a0j1Iz
28G0vvYi28gEfQn/IWxATOH8QIxQFx7SCLWdjTeEzWfDOwrbXHm02PGOyNyzWttb
cKRhfzKW1gpWKSACMd1Hkc03M8rfq0uz2irw8n3HVBhwgr8gSrA62t69Bo1g+ZzG
VPbN8KWcw7ZeC8qvhYeGCU/gJuoAV7P9ojRAheaiNgZsDTV39kUrWbPb+cSdCEbu
J62TC15eETUW5dBZTkipOuGljrOAAZIFUgDKOKlYeW0KXDm65w/FN2hi0QzdOOL2
nMO6EYhaipHuygpMaQtJCnk9UPsgZ/M+OHaOukV60GS9lLd/oFdOf0VRrBcDJxko
R0hvXFtCpfVOK33diziiwRPhaBsjOF71Jzxc6MbnfVqy3BCa5LvPgkdj5FUNOty4
BB8m1MnrSvgqDVPytNSr1VlcEwfFZYl6/SRgPaU7164PRIooFKsdUCcxXRSi/pE9
OsHbeqCLserbfSHiKnT5wM+aRdkEEV5vswoWIpL4SlyPkA5d+HPoNryrZFp4qjD3
U4XVdag/eQPcZlooBJ3mZ++fqWN3O2m0BtGLpfAo3MPAnQKDJvebw6Xq28cPvRIF
wXX6Lh+CAh36To8Xma+sYOrADG7SrUv8vcpKTwvNeNZyOJ0rmrapwau6GXkcS5+O
2HC1v5vvva+OxU1qdUkyb4vuajeyKWNsNrzJe9exa+u9M2LvcW5vWHTEejTq7qCO
cq2PYURHw8GxcWB/6jmKSFUaHfDlbXSwgoGuEt0vckqmnv7GRW21LJZy5LHy4gXv
MBQFfLUO5l0qq7UmfTfWsYBa6YHkBkQ7FNyPF2OAzG3sbmX55SbehLvhCaH01Nae
b4QLHY7G2CBPthJkLGM8uBltaiPxTfmb/BGRVFtsemq7lD5+gEosE20QcdhchEug
tgJ83O+CdmxPXBGX9sI9d7iBvEvDTNfBgjbs8WSObLOBPOt+bWmtcptaiZ+Edq1d
ezzahLIyZTrNVNNLnTvy2AFwWIrSQb5o7E+0Uin4LImuFecQlP9UXgZKO3wToof5
PJW3ntaaE+71Qtvt1tOblEdcnXkGG4EqanMruJuO+Fvn02wFAXSFzppchvMnyihI
0OTSWn0eX06+zsuoNCJ+9e97p+yG3LwHXdgvjKUpiFm4/EsfwWottqg11Rxqfiu0
FAOJb98fg3xeH8GOH1mD83iGYgtZ3rkLChkUOxkz+V0BqyKPX2Cu04t7xsQnlEQ5
kfZQJ53pUoN03XWtIXAYP0AXNAriBTHa8BJHWFYVUEzW8MjX7Xudly0WLs5ndkxs
V1Z1duRCwc0Hk3vez6rq/LeSYE98cu3Jz+ghUEX+YWCsE+iqwhD2xLCdK54Fvhrn
FtqVTotZGAn80R+SJpOfd5u4LtF2Dl2KkYQUrnapx0QrRj51UXWolf08PayHj4mS
3bpNeBU/JHYu6StCZEJQ3cmeYVC4K+F3ys55BlhjJIcz1I3H+1xqDbBqZFbPIsbG
qaZuzrMsqtTpqNw4w34+LPwsJUHMk+UTd/Sqi6fFVKvXIVr11CtKMeTu9+Ax3W8n
zhMGG5hxEp+bACSYKPSWggbcfdAyTPZi/dO6iSVXtNpuCwkWDrdUu5j5GYeD/QDD
K0U8ujcLM7+OC+vxCz5vwYH/ECc8gMFjX3A6fytpNEE3EwzTGPeBPfmZQaTJkumy
cL70ChjQZEmXFmg1L6oSYaesxFrIFtlCoyKJlW9TIEV5NF5jbkl8VjR8o8USBuIe
0waz+NUs77sA2hJqJiXI8f2pfO2S1qsCYashcsMKYUziOHmRh/hHO7ht/qhP0NpH
LniYzZ7Be2cEnxHU7DSJ1ycJQ962Wvpxqa/TZjX2GygiYNe/TNVg3rzDaeGyyMiV
8RBemSeKuQqjJs/xh/hUMSBIYOS6ReEgOLmgIGnudcZnrbLuFSEOzJcyYBbv3qyr
Ry0hivIEh1NdMcrBzQScEQwdj5pr7Ik4vZHHum8+zPDIw4bOVXi20N7t//CP0/S5
tSp0y+0C/n0j+xqSfUYfLdsR14lIL1L2oi7LYu8o5tT1RVlylNIOT+oDHXsj6Luy
FBEu3kurPfoYgPygjW5emOuqJqZkINgOQA1JMTMOYpjYRfC9ICrq/G5TeGAfmnpy
QufoX48ikynO+ObObvkiiaxTDYbtI2ECQSASweQMsBRoqhPToUuTk/e5crjyx13x
oy/8FmQNJ8vQ3H4WoOH0+82fYKPEFUZaiIy/+AtOEuC50w2JVu9rxRhhKvfhlIUp
Zds9QmjIZMK8ThCzY6cAjL+DnxbNpr1j7DRiOf48x6MX92Qx6mG3QO90JIUC2zJD
Es49ua8JZeQXSz9IOkP/iMGVGeQikLKypGsL2QhUA0wHIL2Mje/FKpkok2ywoVjm
xxo0Zaeizit9FclmkKBEoR3BzS5dK251oqC2eT6+2/fkVPLE5SzHCxckGcaxfh4U
GDdOazD9+62gpim6GKmZJ42HbfbANAET4UON5m37hw5ZBzG36Ijy7WV9nZ+wBCb3
n46wO0lTcbEFCU7o5n50o+9YI898Z1G63ri9OJwvjEmNCKCYlHrGqbO1VAvKYFZF
S9wf3SI2tsGCGU8Ob88rGToAk7aAp+lSVmV+PnogUEuH2fsBn/7BezlOQrTBNvbr
mXtjQ/drzBIhfqDbFAZCEeQPhQR+o9mEr9R+upCEtYzfLYIf5KJnTahxFeGgneEh
2hAIE6NH2JxkGJTXN12ciOktFOJFw19R0ivugb+OFVHq2HTAFr+4llgbsNvrr/VW
MfPafc5LQlOheT2bt4xYudPk3z1iUsBROudPKFuz9w1jhheIzkmKZkW+YCXXdVCe
9FdmSVLDn75+buWxyjCdCckjs9v9ZL4xp54AqXYmGa1hrn/Gcb6Suy5jooSrcjDj
lb4+paR1+wpwcm2gQUJ4r2SJPtBKBRbMM5pVyFFgLjovFx3vqrI4tWWDGOvxusE4
rDXDIArsVh6eoDqmMrgG6hgB6hJSkUonHxnSTkdX+0cajyRASXthrBVkANyDgLzF
IR1C+USJnBa8/q7AcJcrun1GPysRmN9yNjkwha7TqhfS9bNV932GR/olFhr7FVc+
7ncQQaf/wm1w0r/hWl3DgOFzdF0mKsReP51djeGL1LrQRgBsNfgkkzG60mh7dQJz
RnmKcOqzKXCdFze4w+6yF3Qdyykb6RO6NYnZBNBmpRL1Mgy7WQLjCpj4hC/V5a9Q
6VtEehK2+KiDvDvCd0Qeue9R41qvjiD7Oh2YWTMqUMO+eCXR5t9oipUIwMCcRL1d
ZOmbtiBu6098Wn8AyUn3Nihqy9qIvy2dGXB4syzlz7pq/S0CgHTWNHmceE5hEh7p
CavHMvpHb1vZohco3noX+KZ6zw4rM90fgBtihqspeLfyJQ+Z8Emd9UipWAWUr2Ct
XSI6kwHhbZes9oK62wzJvLu1eo7cxz4rdWJqye6HHNNV7ALtVS7N9QZaTtCB34JZ
5vPGzVNTos2Yvd7GBPkU+4Mo/S1vPQL6HShthv5fH+fu8XEd875yf5F/hfIGkzvO
WsXjnnL6O1bVmmi7vFv5cPTv+gCWEcbBhD0Fb5mfU4IMMimBnr1HurF9wh2wNW0d
wSSDtBNk2Ape7Z/UtX5+RwlNmKuzclwvOb1OhkLDdqZuAXvRP56KbW3Oq2/kiGJs
hxpkXjSqK8iFFmqF+LHT4xQIIUbqtrXEzsZBAGYdMuDQ8+EYItLy/n8DUqiT3g6l
3L//Lvg6G2Mg1HitbMLeAf7NA3AttVBwFiB87AchGpvK+f6V7P8rNzqGVnfmmewT
JyPp3HflKqBrx8vATFF33kOcf8Sy4QTJHx2uF78tI9+8Ml+2v2lq47EQtLjIGwnA
MdykuYwcILcJ65F4GEWdSEg4qPt6NiECPHc8xYRJjd4IQxa/rn1rsX7CyyE6sNPT
QbAdyFt5r531xsrOREpJ46OmBzkL5bHD1VlaEYTe3VgFs+DrwGCvL/4R5GDMbl+D
F+r1AEfCO0idV3BjDQhMs/bmdhQn/Fa6zKY0MFuf4xOE0dUpA/Bw8ttTLX2WmVsP
huIML18hFAYfODeWfkYr0NdR1zzWSw1ZbLAnCWFoQ3eKgkFUJKdNg2xde0VEnqBK
9vQSIAi+/pbuddpKqyUqwgsduI2cqUqiYirs+vYWluz9U/VIrSdHdm/xWem3U9Ot
Kdw1gPwsIhl6syOOy74h73mGEVeZQrW2x7MbXOTNpfnoatSwp4wgtKGP8MmCs3LI
Lne4240ZU9HIBhPqKkg/tKXebgKkWiMXT9xaqZz9vPfLWf75o+YhOny/5jyRdcZA
QxQ6VyX3gjHHG9Ryg2VjsWhtSelElf8cPUdCTpoANW66fe3+EYSE8EWGkGeV4CRJ
kI3/p/pjUKKKVdxf/7di1cH4mnW1d8v4YOXdzAouP0gqI5ZEKFlvK0AJ0rMi+5Kq
lfiaxOImu+2f8gHSsMoqH+lRe6zmYmdqx57Msi1f5epAj5tPcykm1P1AfCb/72Tz
WTs1r20pJyg2ZChI2YUxh5w7yfRL2LU29cq+lBKTudUkyGTYIzFBfiuZEuC2KcuF
zlhwjoM3bJGtn4pu3HzwhH6f/Y8x4BhpnjLysP7A8cu8WWdFSlfdf3D5ZD2vI/2u
HEqK0x+6V1odbOx6egG4MFR4+6l67CX2q5YFBdOeCl4u9DwrdSU1KCAfDOE5sM4Y
arTf2XoTtZmiFekAgwmXATBWdNslG+NOVViLLId3qcgHG2BLLdkY9l9CRa4msq0A
veXygr7mBb99vTG1NlxWLDYrL9GNnA7Ell4MqlDIxxWUvcXoUSsiJMYDN/qh6xT1
5pWRu1r6vUlDL59v3uL9mugiY/9dMp6gURh613jsa7GfGb6grvvGxnpGjSdx9HyB
FJ2mdyDUVSZPQBS5DFd3LaDt/35DqxlOfkXSgDrPWokX+CZTDUOCUxXDbanATTrW
aZozLyjtYwvwbg6TmRySahuTZEjCjUjaCUT2qz/3hL74grPVzOSqs+ielUV4Y02d
rg0JAv9SP16aVSIvozPwpaEFXWdIQ+Y6plw5NIZpCvZypV/DgRloFm0bMGoumxW0
lvdFA0VJYXb4sgSRsptHjEEQZGzbqN2LIRzE4IxH93HziPlxlar7DbbBvoLWJ6nh
BIgYHbiSwT9aoGv/IsH4iR5+ExSVWjnweDy0mLcnZSdSDtb72W4XHbCjXPKmRgyx
CEDw+T24t2KvhADrT4UIGywvUxK1pmV/Q20N6MKx9NCTH2zcBqIxQMvzC1DrPyg4
UxstmCwZfezzNi6SHK8MMrtlzDnZUf5gF1CowXCdkSg8j7wm1pCRebsLd1IKP2HB
xHjtGWJG9BDbciZDyPFXjs+DK2QA+jGqSy5c1CBgUXeJSeT9OaiPV2Iq5pVd9aLs
JU6Rgf6PgjxPzPvvzCwUjXKHgS9Y58ZGpDR8wHQmJxns5neKv1BhJKLcxVpFy9XL
rOOCcNtO5VOElGduOgOYEO/HRWHiBD6gwMFoqhn53UWMdRdgWAVfVtpQnWtP72m8
BiYXyiFtQEuB9V9Mmh4zkG39wuOKmGo3hJIcckXz8GI6pX2uKFej58+PJZ62NXxn
Z2h4sHCc1RYBrwWhCZoAzYUPhrFjog6HkXwqekkRxfx4Iyo5MzOoPGWC4C7pvoDt
F6uyk0l8sKMfOXnx6H9cCnX4IwP6ZlKHpxEEE/GgeQec5y+h7NGyX6I0tXTxWwwM
t6iLMa+5C/dPlfzE+KioKf58a70MoynXQ9ASGxJyYY5OVHl/IXjXoXsJIWqOPO7t
B0UyTDyRAn7twO6XFUz2Ln/2d49s7XCnVm7jkKAzUM758EcHj8wR0xrr9bsubj0Z
FED5a+LEcT/6IYZfHJuqaCpwLUg7zr/hAM4iyninWGte/uK3QdLcUQmJhYL3crUU
gErD9uH12TWxwbdzuVodkYgdYOTymyokFmrNiemBlvduWHqxqbtIxpegFK5hQkOT
/QtZhWAp/wgZ1zOrQSBQ42JOXs4TqfsHX0Her0B4P+6/7jEVdAJG5D5OPDFwXcMZ
FVQ80jGNm+wTYdWyp66T74DTAz0WE1iBHws5tIZ2P/bcR2P0THzHi9RaSHroruj5
qs37KWkcQSAf+bCGRgNFJFfrIuVMcqKS2hltHRXJT7akyr0l9/wmzXMlRIIJwazr
tVE5elz2XQzCnhiaqKW0ykV5DDCGzY3jF5E7Cy29OzL7wYzlQt3HMWX/+Lo41dcG
MUOf2bi+mo29rqEwjsO14RwSIxX9qor1KLUTQldmGc/DPZysGeaZWqfYRhGfeq6u
UevyD/tM0i/Q7MLZu7y/KaL3eqpOJ0S2GhUHaXB8wsUmjAnFp568JDQ3iUtIIgdq
DytSqWdre7HlJi0WbbHvYkMJVS/1z32JaSFyJJcSt8fqT+TrX02bGNkb56MeRyhW
TD7afw4CIM+Zhq+k23fAs7hyY4ZIVy6pcM10Avl/st6dDX490SephF1hrm/AtLfw
/NkGy37P0yeVJO5WXtKwYCX/W7NpDxjRK727fI1SGZiLfGxe8s0lq6S+XEld5bDV
5Y+jkOOaasltOHSftuaDTWKzKkRS89xcp4f0nGDtMj+gK0nx3Xi9KFB7uoa0KXnK
GvfcPR808zSBDAtJpeoxJQuvpLco0kyBO2dHXoL1psoDbql+YnYxhvgX2JNHIxeq
fZ7zYuekt6P31e77zWKaNB+MvicSV/Ip6ON6Ro9VJG8IuqeAZezDCgRXIA0upJGa
OFtrLfMOePF9KS5Mlh0j7VRY4wZYlu/cw9H6882s3fERT6BCVj9N9t0oKaPRYez3
huypqvQWs3vrUX0oqDpUmQdruyG/cuHKLxflmCWMmuV/M4KfgXvLL7wufViFHpOg
IM0COP642U2lgjt57NeKTJgV5DgvnHvXsBWCpqcyJdskdLA3PeZhtoNk9SKWUJoV
iwzSEHvGPvnbeyLkiYwyn4RfS+9lp9aGBPa78ZxwbnAUDwkNx+9+ooN9Al7mkTL+
SUqzhqlUlbZ2PvGwh0MDGta21h51PyYpxAulq2zKTDGtKuK+nP+fsCgrryowgIN5
OeYmPTgtZWVeZCIx7Sb/25gOQC8U9crflDESvSO03Doe7Ygq84iVXzRdoTrScKRZ
loYdmrGXbjBBBPIN7NtjlNgsRgM+RLXhEn//XMi81mlaLeL1RY3anoc+/CEfnJG6
aPl2NqOxiK198YGcrBP035gXrhbj7XQVQzWOHauZpHU1aFKjmi1eVslQuy3P4BsV
MdMxtj6P2LpmjK7aoKRKPyk+I6fqmzNhssylVgeb8PONoEuTGmjaYQqXSIAuaVal
bb1UWdu8qyxLXOiSG1wOFeP9N9kChY69b0k+kxA7ES16Di/psr1QW1cmbIw9xqB2
YM3zGoN4W2VsoRQZioWK0c2KUuPInnq3TshRNXnLfjg0y0b2p44pNMuP8I7k14xd
a7OfozqF3VF931+yln4oBSvkXZldA3loX0hpan5oudJdz0Y4fzCN7dMcXQ+0d+RT
lzJn3F7cbltZ9ryfC05sYDL5RLUDmxhc0IwWIsKRdW0Y6/bTJ1MTQZMZHhn04yK0
P3HAXU06OeOL49sZhmn5+pX0pneZIsPi3TbB8pixIHCI0s2jK4iAM1103zBw/E42
ZeN2yusTfCFeSY1hTBqY5OlDY27oO7Tr9eg3Qka7OigYW9nxdFlmhiI49ZqoUpQ9
vLHfZNGnoVXZSGugB6cfUKrXtsjdlNNT8BxHdTYu7ymuHEoPijm7zbjLVYV7ozRu
5UCE44phkAqfuaj66IkrhyYCJR78qWqFUtCtUpA5s7eWns6T92PGcRJDLl8lUaNs
0weJeoY47iKEdixu+9P0qTF2iOXLmxFiZP8MgTEh72m0uCqoqHKc47eJGbD1CWff
u/TgBu2Kv8eyggUcWGLVcT2HkVwBCd+8pyKoEfzA6N766nfV3HUx5NvwS+i1efN4
Ai6ZncrzTSXQ28KWF7epO5/3vY/ZhO/lxyLSLjCgP1Ho6Iux5loivLpZpPBfgEmC
BhLRT31nklyvFkM/G4brvCxIw9MRHYpqotGxMdQphzjDyq+Gvgf6q9IjJAOfxDRq
T4bn4RUVTZQg7T7KpJQ33rEl9lmCoDXt7aW32+HKK2Y+tDSbEeXpXzDYiSntZS55
g9Rqb2IE8Vz8VfkpQ2pT6HzfG3SYSK24Hk3Nnvv+SVwSYgMRAD9Wk+lGDmTEBUN0
ydSmTmtUTksudrd111yiPgv9UFB/lvWf9PqC92IoPbYcrqnLWYUsMHUYiLrYbXYo
xhXd4SkxASZdiqVD0HxiN0DVhc+wzm2DNNmponW6El7U0blyHdiy3S4ScOtYVCJl
cgm9Y+n2pt3kjXPMa03dTPO1/BhMy5NaFmFm5JQclYKja3ZbAaBWAwax4Zc0Hl9z
FGW5X4f9NF8o0kOGKUj4sUeAF0QWwnr1+Ue0JCqYCHeWYbCdzcSAd9EUyidlLH4j
tg3GeQLDFMFuBCTR8nA4cifQY6J0Hno/Rx08M0FxZSEOd36rW2vaijYpaMPqwboH
lRlNY9Z7p26/kMZMu0rqgI3qSf0oXEeFXczYVVA4yDUvzl6AN3jxdoCJ3R32PqVg
P8HRqHwo3z11uw/PqDpcBBSQD7k6Qb5h8aBpCqJ6tg/Pgp01lipi/y09W2tFWuik
/pxgtaxwVrawNKRKVEtivFrG5QHEQCSp4TKgS/ZAi/LZUcfENkWYIn7Sv9zGm9QU
95/qvauS2Gnyzx9YapAkpLap1/RwyguOr7Mb3HRKff3nwpQNkakHdTSkc+SBYAJe
FQpnTQB83XssaqqkK5N/ug2USN7cv4zbbblpteBXwOZh3OYmVr18UN8V02cy8ksY
myNdEUpI9DclmEyjYpUPYylRcDFdgajDOwDn/n+rDmKl0r0ijF4Bij2r8ilb/laE
KiSWzdHKSdiSMJssAhe9pvPPFb0O2OVTb59TCIlF7TZERif/uJFJr3Ol+wevhcMa
r2I73bNznaGbn4EBirqAT5y0qLPIGnWrPZGvtZicFipJAWcBggPmX3dRG/vwWho+
AMlJCGrpVzXTTc5WDx5HYn+F3XOVjnqGbDESzODHb4S0N1IFKkTZnaFD3QzB3r3f
qoZ5Or0MUqvSP/qzX1CPmO3GaX8uB9M3x4fub5C7iuiyM47Dh5+4hGlkt/ww7DUE
foH1aLZee773hviqg7YPPvvxCsALcQo5Z1NRRMy4dJJhwCgAk7djGjtDKA6Hlamt
5uO4mP+MgLmTvmArL+U0cjbmiyaZh/znot3+kRIrE6bWaQN2ZAPrr/avtlvCtLlO
agTfcVlWP7pEaoz4kWkJPptsHUFK5SvFUB/U/Q+sK0a3phIRQohMPAZye9wT07dU
/RlMYi+huVCc3MR7b2RF8Ela95XV2jJpIxkeymOgJDCP+psXXkX+5IoBRW7KT1nS
VfA2/SWGSFgBM/qQPvQgQI5jzn0qxTnRe1oPh67LtDDUKRHCC2Hs0SQxYXCzPyb9
V6MJfUIydMMKFNXOvOd6KbMA25AgUos/y6GgVO9f/uCQd0qo6xyTAxd1SOQRHDi5
8FI/HcwKyKnt+KI2Iu//5/rvQjQ2lfcxnMlxTRuIymkcfUIzRXMh8ZtjKOwt2+AN
d0VrD0p6MjfDtDSKcg486A9sHWDlQc/oD/BD2Z7s9pq0NfdlpkM3cDdtCG+4Lay5
ul6nCw5Dyj8DGec065IhfHXZYx28FHVygepCFppBJRnXB2bompO7UTq26jcfQtHV
/h/BaiZnfoHGmhyJpA16w+RvQUwRQ97ds5quWoVCubUGpKFyIj2gJnlIoYPeZak+
xMtCW5yz6qZScdkzHtTp/dUYd/aETBW0q/fM0LxFWUHC5xKQ2Ng5GCDTXD1Ec68r
TsRlud2AMbiHFzCBaGqPRSUwsGPg3koQdYr4agK6bk3CG9PiW0pMrNIl32OW7I0q
RQ6HrTVJxkDM+eQQTSVMs4PL4sIlt6Ni1Y43FT79P6adYDN7ioi1DnVW4cxg+Cmb
OeWWM4LAETRHQ+1vIM/iKGsOGPJ326nSaEXzekJFUdOVbF5t07Ds1u8cDHyPzrW9
PtwT0p1m4bY6obqzxULF7C+Ycl1J09Qbh65kRx0pNZMeYZtELcenraAaHsnI3zYv
9KWoOJofnUoLC6tTbOg//XtZaBH/YiTAiywP9LrCtKIXvHdeWQpI/VrZlwlyEVwZ
Beav7fUKFK1UUfwae1fC+6UOqmFAHhySC5kXfKRqhJdfiYVFZJnD0waiyuJzmyPn
ASu0HP1ai0oOEyX0lmymHxpHaqLuXItjB8JePAH7jJdOT+xaqGUL1EoP9d/allAR
QiEqf/SU7F+jolfbzktgGgG+9pWOcd3O9SX1dGzJ24I/fIskOzNUkH/aygZ15U3d
3R7OoiQ+Yp9swgUK9tS7libLSATmg/RAo2nqPFvkFZZklbGPcpI1A4ry7P/VTi4D
Ehm2LQ5t0osnxYt1d/RQ/zLD4ubWONfD9QuWqE8rdy8OeKrboDzsvKGLvivfwe3U
TVKBOmNqdYk80cOoEFngQuMDbxn4NCREiJoRLzlUZDKrWr0+ApTri5DfhejsIR+V
5GfbKzc25fg4FLD++UCHh5R3g6G/XQtSYkVVe9WMvIfMnWKi2QFCwJRQ9eGxymga
k8q2yXJdrwl/CZuyYZI1Mb+vTVTxMPWktLIwt2HqT2AfwL0cDE1MvxLus2kOP05d
6rVzRkDcMs73DKJkdU0R6wjfqAHksaM6jxPgeZFnV48XjhKGBN71iJskfFeTI0Ym
tPbGxlEcPxcVPvJgBgqN3L8bJK+7hzq7XXy2h2aJHPNjMGsvd6ElWuqMBQ2wFAYZ
tk7eP5u2qWJOWJjygnQ4APoQYIrYaQ26DKWAts01cLRPlUNN/A5LinEroWx2Zu/F
Fl19fAqKW0N6LqLmE0lOXShLEqkps0/CnE0j5KGzGbR1++bo46SlPLNRXuhRR2Kx
93tYlO30jqVnc0t5AGLMpZId7ZT/S0ioRQrY8B2i30FToQ+j+5mdofHBwo+BBxVV
aGtdQ652Vki3pXxkd7MnEioqzSUfJn6SRN61OqzbH9JYRJtirEhu6OFYYXhhmzLg
PYj/AZUiC2pd4A0wSHpmYBucl1oWLYDDsTOxLoyj7VlkY8aQu2W82e/G2HYevzAi
Dh/ygabVTjA09UsGAEbXwzpLk3c4X/nRT/J5Rqr6h+sTaCrIprJH37KRDlbXUmpr
UPQUHRRJQtczug9/wywult0+DQ4hJjUqpKpgcWYiAJ9gAWd8jjDMlHStBB9JBDV/
Uf8p6VqbtR5Z3tPp4+sYVdhrFA0WMHJGfPV/Hq8v5KHG1tJDmA3JC95XiaaNGLtX
BVCD+E4kR/yt90EhscCbzol4lDFnS4/YINQqVXLJ9Xb0lkHWza4Kz6Tg3jyiwmnf
4zPswFsRzQXSkT6TbwSQSXE5jn33GEgXO62V64ORxSEu72p9YEFVxPIVN3MFqK+u
nXWKlo+/v1sigx9T9LsMOMc4EYjAI2LZhOJw9p9CBxX4f9vcU4yZ4vuj5TMvDrpW
jGF0SxozNRafVZivQKSFUAiFn3/DSJOnfiBscBFYhpn2OLuEcPIEsukN3NxXGqcG
3dMN6CiHwIPU0e4gSR2b8xO+kqlCHcD2/OMFy5bTJkCTEPS/oF7tKkeLZrh655GU
4eU2XsTXK2TJSN0swvWJAxRXHYkEa0ROS5EVrb2e8Zv7TK+rFLKLtN/e/WBb31Kn
tfUUMUABnHkGM8/pNtnpl282QoLaM/pv8q39p55IeqxURW8G0imkel+JC/kqCj+o
fzgifxlOkAtWzNlS6z0O6ExQyhNOpTL/BpEfD2DMkqsn9OfeCGKF0ax/sieRTYdI
Pr/rFrVG5uLuuXxJaXnlE4eGlbsB5y88rImrx+LiuKqXQpAwrrCPwb7Ru7JAHdHT
BVNovwXwzRZwch9m4Z0ZetGWQvHh0w5pkozdbI9HiXRSxSCO9hfTP9DiNpuPhSVP
M4nRu0XMyXOJs8o6L/kOPacsKCkuPPwxEZXBpOFNWTosYoPlt9K0DNIkXFl2Hira
ric3XtbmT+RZ6695S/xu1b7gTdCfmHwRP9orEE3KZtw7VlZaGWFUseJOlh9blCOy
4HRA7FFXf6+KI/nJNdwI9Im1ACWCLhbODLxHTGajDSPkSbI6HTh84dYEUuX91KhW
3CbVKdqNmTHiWGfnlLe/i58DMt67IRK4S4PNGHDYdt97Yj2PBIhuLpZbe0pcc76M
RZk9gEo5vqlmN2sgvM+YsitTwNX7f7Sa+Mc2uFIMi7GyCR2JZ+IvvP3qfetWe91W
BD2xrriP3JpqX+2dcf8mFC4LSEeTPgedcm0InCKOPU972GNmKwRqggq5juGg/7Xl
JX4fZpYmTq9HO/JtNqlUIxF7I93Fuc7mxk1PYKuJyA+1eenHe5SK5hyJKIbBHZRi
t5EKJBesPSjWNJaGKxURSVY4ahWP0y3G0bn8GIS9Of+qNjCUPFOmZV4pBPnUnWLu
eUaPj15uMMd3HH7zMelAePlddwpf9ADGyi4oCKSub8yRrMl9kXJiSAzWmzeNC16S
jPHaHnDce/aCXtrUKGDtDCFZNPp8hw+9UKdlH8E1uDV/nWbtVtYA9S4yCu8Esde/
lSby0yCw0sGE3OENABe0DxxRPhLeNOgOW77CzmPW3rheylCOAgF5wpqtC0bC18Rw
m7hlbrilnrK65nViTm5iks5XrVBiFu4ZOAADcpYFGMqkbSmkn5Cf+vHGGr0rjtXa
WDLKaDJiPgW0R3NRnXbvkrux2fSIbj3tOMO5vmm/GRzjg9Wf/JvJlKvkXUydIsx7
hAHtvmpjAONur/yy3/l8QXDq1EXUeeXXCbQxd2Za0c+WXwlFI5GHQlqQEqGMirMR
SZWKg2tefutOHpjzdQMgs3ekiFmd/KCpo2hYaVjS+JLc6iBLCIy/E9msJjdmkvWz
nkslZ1vWuFsKrbaHOhXs3FQHg2G9ioRRpPm8Z3nDXDFID8eE9b8BEeNV4CuZkfrO
qSvoUQ9/9qKSdBmQqoNglmxPmwKFSRyPqw2QziLZCe75BYmRJrtsO+ISc/+U/yls
6kyo6ljNDAdsxtQAoMS+HeU48Al6IEXxxQbFD1265fhsVQDlRlFjuHkeXalvi9yG
tiqwRxEkcWTQfE2nzIzC9wQtzUdAQ7nIZFCCPkXZeCVkhdp9jBjCo8JBSQ+czt1b
G8XHoRS+mfjD3aGv/vv9q5z2N9pXHm/zIptL41zfsTn9PC0LCWdVZU/C22BRkDLg
gTxciA34lqPfPW+WQiLW00Lmq+JTALhmtHIpwqOSVDXt6v8Zbxsb1vrrsImyETnc
V/6+kqCJrAJ8V7PXDnvY2KsuRNkzeKYBqIx4V0eYPxCgOV4VLHk2IKNXOeKcyMXC
lUzd7IflNzyk/x99zlL2sHccp9CLKCGfxbIInwmgENBqPdOGhxmPscDCdSAHuKtg
bjUjInE5Q+so45h16gPz7rgUdHGID84jcecmpvyV5TnpnfcsXvPIs9sFI6ixwoXO
dt80SdarSH1wb3kSmDU4SGi2ZsHXPl8XVVGZ3kfbIhUre77PQi3PoU5hFmR8Rj7H
Xz/JNgfksnbjYmr7hdQxUscCXcqtXSGAxL1bkZ2Ns9nQIGWqRmg26HoPHQowubLO
m6cNQFeaiS+EAA2GIJYVo8RjUr4+7LG62/G3ioSeF3QGLQ/4HfdEFzUrDroP6+qB
oobbQuVyrrna7YxmNIxUZ2JSc5KkkhNfHosgC82Gyh/xNvjjpTfwT5cRIGwmxM2Y
oP2Kuv8ph3myLZrKr81PxhMOcsfxetxdmob3TPBoh7mXZ+1LMXxuw2GjPelhNuci
PCSdn+uhdI7EJNKPTBU4W57JxKuIuTniYoY7xpujbrUs3lhg0NTY6111oOeil4Mw
PwRm6/SyY2p8zTPdYjzwGdD9iSAKYUSBZYPVWjNpQByqeV1+6wq8DZZeCYmew9M+
jx3kELXGZmPt+M97asHmptQl7pAYduMQtUI4N4kNgrIYMzD5eBAb46jCgFYDdDfs
AjoLgnszCsvwV5betXjZ5WoR4Fmvg1pYYtoTTT1MgffimN4KLPUpzBU8gDcyc+SJ
7cgWopKKRcY6rtjqLQjc/VFeebaxErt5Bz4xxfmJOHflYgByN9kjkZYSZ0fcG0gI
ohfkCeXFjBnXTppFKxHaFe1GompTZutcpiS8h2+8j1hnQqWblRRTUI3Ne1NvzOEq
acVtqPwYr1aPWBcnMlRcKhsUaGCupsT6GQ9BvGZ8stT1BDu18kbQ3bZbjaZlFHvS
MkdxyoXwS5OWsdsplq4nEwudd0lfBeor/TU9vZTAUY1dzEYMSR5TTjRkkmDMoUuK
egGC0Go4QvU8Re+7IJEN5QZIBFMmeBztV80umy0mlo9Qsp1zNuAHMMa0nzznDBho
Ex+r6HRkNzD/FlSyXq+QbD9EavwJtrZV7p5bxV6SM2ylifEYEeUscZrX9a4aWVhe
FGzL3I31mEKYbyiylzmp4+mQsTq6YZp2cZp6dhuiZmNsT2s4mmbCxek2E8ZU243f
RBFc5bIAJ9Y8e1786HUdhJKAtYmUVF8MStO5odRYNo1hM+MkFaEveA45Cix1Vz4T
ATDm0V3Cws65D8eutTPvNih3NiBslgpJo6l3U+1zESzDJVv/+q6zhIJM6EQuAFK4
UGGRVQTCA40TS/pbOKS9dbxMEw2iXuhq2Zv1o1/kgkDSLGVHTs6aAihTwmWEn9SL
pm51MrPPFsYU8poNBSN0PP9NlQY47wpLBPTuY96/EO/so8CH9P7z744I1cWpBHjg
LGPxYr7fE8JlP8S2p3fjP1B7QX7DIbD9zU+EZbJPkjrE5PdOFn5S1QuX+m+gaCiz
d9zWvOcRFPbede68O6NL0QcmpopuK2XqlKjCXUJXtyiXswQBwY1uHX2+yK6MmHCy
qQL/gGNfBM1gNIRAK9wOMh/nF0EALpBIDiKAe7D1CGpeIcUswejOmnmcydrJ+WiF
HnTOkKwbRQdrr+xbUczsnXlsoZOjlbduFod6o1UfPkj2A2PsROzfyRM5Hv+t3Esq
l1cp8FKozYa69XiMfQWOAa6Taastf1wqWjOa60oMRfVesqyr1d1O3KePdV9KfB32
vcHtImPJzusIrBXFaSz6QJV2jseKPpMQU4uofy4RM7nuEQxqDvdNIUofQiBvTwyE
0431P2mEZwayNLTAip8hKE3Smhx4Nvi8mWd6KRBtBBiWJBuY3FoYCZwHu6v+ibKM
cVa7JlnCUglXHli5HJYOrxpw+HmtKncPBIrTLhuUcOgnzCp6k9hEwQjx3n1J8HHk
r1iJSb53D6y0DFtacFZezOlYU9DhatM6gB9iNS3y91k1MHES5hF4HfwW2yh1p/Ck
fIv+r2Rb6py5Try5ykI1THw1x42+mxMZuDEzFMJIhsynqOHmGCaZI85WSKrAxFsY
LNyKg3iUs5dqRqajJEQAbsVhnujhpoth5aYFForNqEQS5N4xsfCJp+rgLBEWSWg/
kCIKtgggNANKbgTX2ZW3FXdE0SoeG3BMqHsv+S8marvq7jWo2i8CbPP3lgxl0EFQ
yvKVe7LKbXSempSDe1xcZrU96Q+P1OU+ZMsF/PfJ3fbYK+OVV9RjYCJyzHRo2SCS
o25ZPN9xFrCecPKWfxozORYBZjzhnrzhdLC7F4EukS9JC74h0lNOl/41tMdPuARf
xUvRxFfzfT3zuwH7grdVdfM67MSTIisztKYc60T2eikODIcx/APEWitjo8v0U7ru
69T9SlGsJ2mE8ldgULCVN5+S2dLCoS7XkgJ9sBlKcKNU/g4DsbcjfMmniJU0f/n7
dkr6NfZuAgV4/KmJv6eLIOTlBIYgtNZJG7jfzhz/z6YYqRNV4qRYqsV+r62GjuGy
07C3ZUCctgMD+XF8rPW+0D6lNfDNSOjWjMqlkUR+yH+24kxN/PGtpIO8zXkyF9JE
yqEcfTCF31V9l+ghdH2ZKYKyD+8mUL8t3NhidF+xPoBnE07brAnl2nUzalE2Liwx
YMzrhMgqhjQCtkVB9kJFlna6hxD2l38ZY4Nu5XkfxRN0xIFDR00yOWRvaRQayZf2
6VYvnz2TTYZZKap6MnvjJvqM5vWEd7rYkWDHV7xskqQHQRBfO9pQeZjd1iFn0ACt
HFnRCQo9qUl+agYZr8b9noiJUpBGP7hBgMN9Afa4NbS2HT/QDuAI6dOpmPC9LbzC
4e04YZ2+8ZXpWlXt1tXnweUpBqXas2NJd6sZlyGmqX7BKcZtTn2/jF7S8T5o21hT
UFqRRiAXA4Z2c8l/VvKs6U8teTJk4asIRYjyxFXQlZOQloZLuCunoykXzO4EMPhd
jgpXDW9xG4qxS8yzCtnuI1e6RFnZyPKaT1tXV6jN+I+LCcojRPqfIsuAjaiScTPp
iRJ17lLi6QNikLBcUN/g/lhe0FoYrLatjXDffWgZznrpgbgXais4Pvs5o37WwHf9
Y41nnLcK4MdpTTPZp+nIC/xRi21mS7Pdjrvp3gbx2IfoM1ZBCRbKBPgqusqp/z2o
OifBh4BTQ9qWF9C1q+eCueMqlVY6Jb6Hhl87lz/XzNycCmlKA7PRO9KCTJI0+iYD
3Kq1Jhbqx0REpqQaGObkwubFj2/fKrNEy4j8sA8Kb+KN0njrqFWhtmpG1FWe4X3S
oS5yObvjlBYE4ONxYqSjbgaGR9jd1akk4sBcBVwI6bEiEJvUZwoK/4DfMbRMCJTs
Hv1fvQxWx8pdDpJ+9KiHl0WAP2f1HfXcn7QgnAANT3KcG63Ge6QpmTwd1MX+VxkU
oi5GztWqQAv3za+5H4pwjdsBMTHX1yER9hYVbCeWOkdtdcmxqNbP+psMZirvrnSd
EfcS/XWrSwqFtRks1HKDjdZgY51GH3Vevm9lrAUxX6bO3eK1sz6x1Ku251Qkqnok
WMk2kCvbVPKR/umrJ095G7G0sZXQ2byEeE6g2jr10Kw5Ekq4v6FiKu/es/UodLnu
Sr+QGPgXK8GVs+DUPJvGjxkqeHTFKSirsOkULJ73o/odSGQJJOfzlC9VPcWObTBT
r8iZv3E1/m3XAO9uMpWLkdDWIXjk3aA4/8WXvoGacPmhDPoFElGycjM0GtVgKRat
Aejn83GAd/7yGMJTAGNONAVvObZZpW436OVpcCe4BW5JHSikgco11tLHF2Ih0tOe
x5NlgzCWzI3JtabTysSHCxGYwvf3iCqChUyboEyLTn56zS1NG0XkStfWlgNEpTqS
gaEem7GKDeLDH6KLpCGgmvzrLq88gcGTFb9xCi+QxtnLqYMehQqRiV/vWGMdcFU5
58SrHCxn5E+Tcyf76V+/6R4Xo1g2p6pysWaL3cJqHwlseX/U0ELthvCwCh9qJtWg
5XBeBsSqT8HGGkNw2RrB0xuOAJV1hSJIP5RNElgJ0ppTm0qIKUSvR+g8xnmWbfXl
piTLWu/7+72Hwz6u+Ov6Cz5zLjKpwuS41hO+CHVMoDcGN1vjAOPVOL+lpE5CHoYy
4Op2StuwnA2r1EQ6ZsJ3k6icmQMaIxVUFDNsATGDwVFqfcmZKUTO+RqoeSKf4a07
jRndEmZj0t91GXmaH22YpAV5W2IJb3Y/e0RdFp22+U+oOMMFHO+5ewzEF5sJJPps
0IAMI/yzZawDhrkolBNDLq6DSqXbWRT7MaoMy7HjpLHZsKULK8uiHaBqua/8kOow
1EAfpSB97U0ztYrH4SKDHMD2JrBRwk6SvLh5axVqXetQgiZ0uzD6hvzicUsJEpMH
Bx8rs3Vuc5i2ooUummm4GQx8bBw2QHBF/KFDc9eSlObxf5OpHutQaXLhCQllv8nG
+6o3Jw4J3QfH1KXioB1+tjZ9FaKbHTqEBp3l5+AjVBchg6Z3vsN2rKPgsXOKvMna
kT0436SNX4+zFbgr0lY4oHwT2cZIO6xESHZ0fNeWeGivjVWzjjPX55AL15k1mdKy
OFmsHUeoix4kHXfc+J0+S/02cmugrLt3NPp3+nZkyF28Ws81lqCXyOjxrGxpNZZ0
Dwwv5L22z1wRbmf1RMq7u56uxc73YP7bHUIJ8AdQbeMZ0BoqPUoD7mNZjFvWvdni
0cuZwKLgfhFOpbtzeK5koHWVyvyCbLB4WGQxx1Xz83Fz/nGLGjLoRFPOv4onbtKO
nxphDGx3V1e4IEzVNroIQzai1c4tX5IaAoVB3pn29Uk9uzXJMXFji2la1Lzfxf9J
lXtKO9AezQ/+Lstadpzg2kfEy9Sy7qHObXGxVPoJIXmWac9a4k7wxEZSZXKVtYFW
ZVX92q4fYr7K6eNUrm+dPlN0o8rNTZjs0sJc6gYp7Si0fx8tuu30PQgVG0q08pb9
kYFqKsUbtHUnSMNIEgz68gTNu+K6b6lNGAZgFUI4UDPF4nJyPzjxLYSSyd90Viny
9m1v3E9MbDpGph459uGJyRbHPro0AdIwwkYzQ7bnrbEAmNBlOgNkbA/Do0zKS3r5
NdVc8LCz6Fdup3R2oTupGVPVtjpwhiigZn0AbKH4stRlJgfORgCe7GpVL7rz5ugj
40m4Upb/MmVFdb5j0QkwfCz8ocNC8/qY/EMFsYM7QHavmB0MNoxC80cwWDXJ3J0S
YrD4QR8GbC1plkPvMfefI1mUeI0FoRHlm/ihRDaxUKKcjTBmupgCJLVln53HyK/3
KP0U5LrYvGFuiVjMIptuGpBbIovCxcUfQ4kgzlba+I/T1dX+VW2i/1KecSNpG1vn
mPwbSyr4cPDhtno/dRk40b3DW9tXN0ICqb3av73UVZMv58bcAvmkAGxmvzZNCZ9V
h4om0RUi3ro3bxxbgaw9KWMeeaB2SzHz+FRh5J9G4wN+Dkl3n5oIUt87j16MW5ME
Mggp/nHirKl4xf1wQ1w/B/iivYl92mrOHYPq2FC/fl3ZXmEiPbIM1/8lq9j8Bw0J
SoiTAvyjLJOCii/65Zegld570hXG70+F+XV4arqIvdYETrWVt01Z/2/UcXDivKSb
Gd9FqCXOi11RBJy2ddM1UrNjZS0QIpMTNkMcplomVzRhKKRTGMaytXCgkuTJTBke
joaK086bgXO2TCg88MBhoJGPEx986ZuJNqDmVWrA75fUDB5UlITfCiUo7Ca7GUPj
7eAtYN680TRNknybTySVUoPO6XwxnFN1DmKgCZwYzn6vL/LJDYaThi5Bjaobst2/
JMBlMqNT1dlvg5aZZZ7VBBzpap1pdrUVT9YqydU8WQIosGbecxH6C8YoAw0n7fY5
DHDW3KExpUWmQqNa/jPQTYU73hBZ+/da1KMSkCM5SQq9s6DxKS9VBi5X0WaiRUJL
siMSy4hC8TkoRr5MFTGirJ5Rh65IuTwTDbqjGjZPIo/iQrH7OFUImcuvS/K5/aul
TifKvgyZ1Gu7gzxW93BUCkSs4MftwOXAIa4TZRLU6OPg3N4yoRjYF52Qgh0kcH+z
61Vrq/0eYMyMSTatgC2Wd6c/E/qojYOOFO0qdYFf/g6MqkttQR3ZwKV+lRdaKGmw
wG5j0W8NZ9ULFowTE4JZhz0+6i9HKjneUROqhpFVlcjJ+dbWSnMyxcM9pwaN7/As
c9Ysptfn9Rxc3pAHF+2J3unOsDbrPlIRPy+4ludENy/z7joVOGXrCYwut4tJZedo
jaO3LFfUHMAP0vMAEMAPndxV0V5rkkg+ONFTE1AB1zB0SFsdcXY/a6fESSGt31rj
Jadxg8tHW1Z+YpKvDTT/pdpi12jXstAbdRpn/iHd+48DAxZvBtcDYy0yDSRQ19cf
CUzyB4Z8xLyAjyB3w49vrTH4ylonR8HfJnwIPQGdXSRkQNRv59BZVbGN1NEA62q1
Wh/YvlkMeP9X7qB2a1G/umrXV9cA9K08iIuo2wDIPMVvNPGP4XDcLFYy7V9BC/nT
LNZQa9vtXLjudr33mU6H4BbGAy3VYd7MPilJ/L4uG8LVHnT6zN67cyBEvrzxTSWp
59ZdTfXI29zcsW8vZGmsuXwe3LaVnEERc1y1rFmEkxVaaEz3wSDs44ieacHvTZHb
0RAY/aRdtqZ+joQHqSmaQCNQ/mA+w5S9es57FIKPzK3eTBY5yQjwAE833YoczZhe
GAfcPrh7HizXHnryrGPEtLSMVfG0+fQCuXDwnzJY0Y8IIt+oqZAdAEr41+Qy3SjC
Z662JppkhXGB/nxlrdo3tsBY7/3hrRs4iMZv4hVFBShxfmjaCDhXqIdSJW0QmBFe
r7RV1q/7eT/aKTF0fTdsJRWNhjzezZOODA5ojnz60oFiTY+mtP2v+oNiq39UYMEF
Gyg7I1QoDIyDPUZFzzejYSzfEEdELMU1D5KDA+dI8Ahm80NfKwIQABR04e52aC1G
KuQCjHcmNplFMb3Cp5c9DLR5Ic/Gfaf7KbvxJ4JaY4vqpsFvadeL0UBjVyASTZ7A
oENcwIARf/LNqkDZWbNjw7btuX8PL+aTHONfxxAK2ycUxSDmxrFEVokuuGbeARFZ
Nfbw5Y9tfITwUf3EupSJtQPR0QZDbihOJp9y7kN20GcImAlc2YEbpdojYGzIJ8bF
S7UesnQQMK6wtnD0goJ/a8j7sOhQYMlOgIQ2iz4jETA44w+anBvtQAPkIasKspXq
nx9kTmCElxNUdw4mOTeDeQpvkgY0CF9kaBHXjfWNEEWhgdjbX/gxJ/+FSFkmoxdZ
Zct7rhA9DwnXK7MF5z9SJOEArikuLTsOPDroHFb+hqpKXtsmoqiMrMGbdfg/nufr
XElGYwWMpztK+l65FHBQpBcvl5k+IHmUmngl58pm+IiJU+VffKT1Fl+3qL8+rjD1
O1HijeGH2hO3NPcMo2XFIl2Gc//Jgr19JzXcs7bnjvIllcdqydv9YxhVy6LJmYi2
zck2MVwplHgzibr7Syc4odiYij5QkKquDO37yc6bZWwnFZG3zyfT6hK/XxTbiQLb
+yhTFV4g6RiuQKg7orKfeCR2SXKMXFMtsDahnuToVNNIIrC8D6Kgp0Btw3Gu9pej
HU/IYtjgPhubwWRLy37rYiPTLB3RwatYfP/3ra8N1ELu5Ww9e00JwGOwlFYm/A+8
WwAz2O27q15XUd5AvD4cymD7eTeyQgwJYuFgqReMKWNfKstyww+hNYPPPYHljYcL
KL1UIYSjA9Q+1gjhbPvNWbx3FwWi8JxrqPvCy45c2XY7Aw2Rgs3sxyUwe3Cyvejs
8fyYiXaeWdUXR8+uk7M8mL4FQSWR364zQFBjpveDSotsLzaF+KOsZo+QpgdlRs4L
13dq6j+41eBeow9eoPmON5X2e88i2y8kkiaRkSJsW4x2cl1QwnPZ3BPx1z1WLAdz
BUGRSEAFd/I4RzXY37EVQgwDBjOoSFELyhCJuZx1EujVtzwA36Z4h2255RFfMQzG
14qjekzB+dpelEYsa6iwpttEs9IWXxviPEGp7uoct6yS0BCvOJatJChTk3sEGsEU
JkkceG43PQ6lpHvuujvnTzXjxxEs2Pw8TYJPyjWPz+lf/eEMzA+SKhayIiQuo8Po
srejWLVkzHoYCEnpHrhG0kZjmrkde830OmYzyRRKStTqvSF29JpljH8Y7b8pl4Uu
DXeaCH0PAQBndrZFqxsklvVU/UVmr05izZqe6yJmsUUJVWOzBySMVDMS6julwsgb
FIHsl679GweP7ZPGmmu0sV3mSMvZDXOsIFyNkyKqaqeU9wQ2A0pgrzXePuuJwbIj
o1QYS0YA2zq5hZQuyqttVrFxR4HxiNUmDJdiZlm8YZ60rB8DxnvAkcES3kRl+o05
WcNK76ZTccw+/BQa/YWAvIDqSfcKLOGErqW2qdj37Eh0bxt7XSBPxsQABy3DeX/8
mAfE6N98K3T7QANgPWnqgau4yjdwcTNGxceNghi88Hcp5ZqEBZwsn7HJPD6t9jat
JZgpzKnOfbtsrH4ScGFWKVVOz8JCHYBgI+85b353cEkMKHbkvDeXpNo77yDu4X0f
9MgK0VBE6H79JoZYz5QTP8iBMJwdH5S6bPHVe0Rp3r/+7mT12zOuXvZ3gfojjyZd
xpqGbms20/plCldYuROZWqyYvEGLlJG0ofexI2ueyrgUsr1tvDSh26XxprwR0BT/
ufHZgKgfB+JZ9ewwGxsa7ZTCzHW1Oe3SziwdXk1kIocywCU/U3OrM+OONwCLtWHg
fBfRZ2hlkXpfWtB21tKIJz/OSfbvGWvzM2vErQND8mSQ0zCbqD+9k5sRUwSPr7p1
oZy2FncHtTp/iSL5vyJ6xI+qc89WNux8Urbl16QSX/ZA3Q4k2GLP3u8VadHWEedg
Dl+BYD5rDhGv1rKHIWOhVYqmNqE207Drubre/ycfLKfxkdycSkGx2IWE+z18Mjso
By8zha+kVv7qPU0i8+ona5o/BwnNUMrmnZud+CifOLF8AmgdYQ2C185x7VDniXHm
tn2OcyLqPehy+ndrGQXLq0D241rICWeuNk6L2lGZEiqPNL3q0r40SHMOzHKT23ry
B9FJV4BNY9xKmsrOM4b2XB1kdSY7A4OfTZQjqfBnOBQhJrid2Jd2eFVFbLpvayOT
rq29ckeOyf2we4Z3W9WP/epXGHK1BHhE8m4Lsd0w+HHju3ti2Mh8QJt+AxcfKNFm
Nw9rzq/7uzD1jmty43Twa0VU3E0DO3XnxC9Vg5K/wfZZXWgr3uIohoFWjKvNriKn
QdEShTs7EVgl24BPIJvNqVcLhnPjLKildtpriOKLGxKjnlWaSJ/XzwbxgZMtp8rB
iRX0njMFT+03dPcDW5gFr1jHPSKHDMo6riUc0maLo7+hWB9PFwlJTfyu6FycqvN6
S1IYFhY/juXMnYkCltr3TQ1yNnTIXmg3MSbH+DaJ89WVNGWuQ/0NSrJELN5uCo4o
DM8yg4O4VFZ6rc/dye37zrQrIAma8WUxX+zuM3GwuuHOynmoEUlFVXuIYyjfFCOn
PnnXz5xBCan5BabsJl3B1Dut/LCyNpMtP4x4rLFt//aU/zJWKtr80SO8hT8HjMoB
vI2O5kzjZefPCNg7xitAiLoa58Eqz3sJD6Mv5ZZHoasPJog1hnwggHp0G8axF+jx
C6sxNb3DcXYUockzLBjBL1BDZcufalTszGf3Pgn8+Rbnbrln7dFuPRQieojobDfp
MY/6mCueL3NqapAnPFk5ZhyPd7QV818+WczdPiOOSsTENEPK0ADHwSuWIiRji0Oj
Z9jEXI1Ta7q+cp6UE/CMBRuwjMNZmkBEx9sEqqOQm+4X6x/tad8mrYHe1/nyhFsK
akdhd5LD/LuUmuBlI4rHM7exPSZPc3vh9aic2nK3pStKHN2vkHcnCB8Pxnv2jdRS
+ctmvZjZHEvbrlECw7rfgjlIsmGqBJ/D3m0Q2+CcRvZAWcoNz16gk8Cgvm23hoyX
1RX067PMVFg1TLiwFHYLFdT07dOwE8hSSoltA7wtOf5o19aeODNxBbsTLfQTc+o9
quoi1bdL20q8XxBqbdWqnCUa3USbjeLa2a2N5iqt4KVh+obDMPrtu4nLBFlD751k
n3siAZkmzZdRB+LnWz7jXVygxw30Yfzg3VVC0Va9KYlV1CYQu/gQrYir7Ss/mSSt
o9nJxgilQL8xhi/VBVxe11Gfua9AVnQ1K0W3K9po/Xjg6FvpeJr3svRKoJVJEQ4r
b6Coe2Vx/OI9o+XSEhisyQQ8fk8rH4Dsm4bISwKbdNwoeICecA8CRH4u6mYWboWX
Zfw+OfT8Jaqxa54VIw0vbxA6hm3q//ThNt/nJw4In/CxKOt9xDdTtCu13Z2/vv8L
jAuekjYlDDFpK5mP0bUnoL6ktBWFLWHntKoTBXgEk1L2s8ZHvDU4K9gS/KZYLpge
YXxRxA6jXgXhFzNIpaw8WL0ls28ivIf9S8GWxpQNaukm2ig4ocbLwDjorRJlVW7V
TqYbAenXBG4tngazQjFyaZvSrxrInxvoqt0+iMpAFfK8EQpZ/Kn1Uc9YET+wtF4f
p0ZBxRX7g7ijPxsU/hiHr2yPj33XhEiYrRwquth9SE09NKWWq14NuKoEP1Vqc6zw
vennFACSbFlqHID7iT5/q9vuErqPegCPa5IM4gZGHAu5/MZxSI4u9zsAFpV1QeoL
80LCu3AaSNp3PXVe8Fqm0WYs2LmWbL5cOSixT+mceVpWHOV9JitEXZzImR6BZdqh
5qevnCEoXIQTtOiR9zDzmsqyQDfh5QtxpNdxGQnHj8rzxVA4pWBbVpWKDjSgUpM7
2IUQtntp0eKUXBbNx1RObSHcrCHBUiWB4zEmRkItMu96/qvJEjXLwQErLwK7+ZNK
sggOTFTKxH0bCflbwxn/MojkokTS0LSQobWbS7uRsI+eNr2EHE4cKgtDfgnI8Cbr
1aXYnwV5Lrx5qWVGYQb+eci+HlJoXPaIeKPVMVrkLgM6vWnOBXjYCjDf2bk0LPSB
4pHW2sQ1mAQaOt4JZTM+Lxgq2bmfqcse4nxekfAkDbB/BaIinPSCz8zmlokAWuGs
Er3jECYLU8eYUF+QrOLAOW0G2z9YSxFVpaaiMaVCPLFmosuxsCpDmmEJXv/8y3Yd
Nrnh3PcswEBAaoK4cxlBuncIwl8tMNO5GxMv/bZ04eN8KxHYvpeA+0kyvWSXhMmF
NvRaj/msvlZjMLB0Shhxe4T6mSNYcXb9d4mwYKJ2foEUy8IB1YfnfizTY1HdAMYv
ELJAlbH0NhgK+HSYQ02usJrPtw07BpJZAibtaIA6TXjjJYe+gi7FIihGoPhIpUgm
KrNwbIUxVc/Xe3ABpfKb14AwFTkJojKr5uIKni0omf6AIERe3Gj0G47taCTlqzQY
YyGfBHys/aSIs7Nf0eka1kqAFh4IX4bDLqL4Ad/PlOYqXsyfCJIfeWWDAR8dlxzQ
evoaaVofHnsZx7fE3d6zfu3HqMteRWLcctBUVGjP/Wf1Uni9aueKI2tXakrRQse+
STrOwz7ah+b7y3fcoAOHDCF8P2HVBuSyLPzDn6tfHMdPdTauUBjmiseRopMLtCRH
tlCZqO/MxOcXxDWxOBnqP/f1l6w+XZYhzDnDpfAh+FIbR/skUTjmVGEZwSiKqmVb
0ldwTJ2KKVHapCaQAj2LhvrM/nCj7IDZ4nmTxs7KCO2fCyMGTsoBAD7uhDZmZgZ/
pK/f7OycCp37RUx7Rih8RjDT37sYDDhGN1TUTRrSUJgZ4oAq/fjVupysi6XYfDYv
Fkd1lqz6P+jgYxwy8q/oQn7gcUG+MzhazEJZJSPinl1TgCQ+Eno16IlJc/h12bTA
VSqIpJ4Pkj8MNSuGjLyYvYSgNGIdR/eEgkzQKXWPl+krZPyNCwBwSsJaiIUwZ40n
CEbFJrb7FpB+k2Y23JYZ7JKo2/XkegnS9Xn7OD1Xlbhrcy8+MzaGUGRTxqQm0Zzd
gmC5nHAcZ9E0UFL5w2h3K3cbByR9mPOXm2qkmvT+qLfv4B930NInh+zAnvwWByR3
S44rXLlUj5z381DeDhWSCV5xOaj5d6fLJgveC5RK3bIdYnUUlFbBcNLNsheLa4H0
3xfXzq+zB0nLdxpdFJk/kekttlhdmS1VqouOFnC5MLCIPc/KVmOIVlz8rxHSbpov
PXlLpMgaV89SfE9+nGQMMwk4YB5ulbLJnSJS9BjjNan1yG5Dv8PL2Rk2IOwKWwnB
T5J9hMaXHCAhQjsnzR185v8m7UFlnTNzJ5imkW78TtWLgTpfOijDYFfulyk236Ka
0ZXpKkFhpG0JiZ8xBd9SqQWNvGvCPaCLwH9OpiRxnEqqYnZibbkYP1vB6sGODOUH
c9zQOIQ0kwc8ckzWYy1+urTY6YgEU1cfsFvB8pOzLje13ypK9YKokaXYUZaMvLfr
LCqd5Fh67/IlIYzvbEtZ/Z4gdsfoPyuNcWwIXCjqGL8Gy7PoR5nOq1jr6i8jnkLo
9DnhKT0l09GftsbVdtz1MNPl77/DUb1v0VDRCzqG20PXbPkMZBFHLPlAXcCKnpea
BQbAd0TUmHZyYq4g80cZbfRC5Q5j5l0c8WJD+5Js/LLSBTJr3H7TcTIFr/pIiHyO
fL14ux3v9Ion/Q2pK7FuX79qxEwHfswhAGt6QTNNKy8/J8JGE1kfD+rWo6U0C3HP
o8hg52+1sdOo/8DlmZYWhbh+KyARIxqYgrFQ3OUgpBISr1YDLSuh1qYC6182cOnD
YMbU7wPs2gyXt2EDXPQm7fBLJm7urlO6txklBCfdEJc6IoHfurdCrpEHcNPMf1eb
SvZxtzVdQabwnatYmP7ZtyOF0PJksawb4LuZx/ndJHGYYzMwwAHqDSHIFq78Tlwc
yXfJ2O0MMwSc6Y9OyMBJBMciP/XnNMmsZoZAcujmm+sLcHWfnWep+aTFpsDsFNxF
MJ02s1fpq1vJFszCS3yCXWJocc8iBGmUWt6A6CIGrSs8k4U9HsbWtqqf+ZvqSD82
MOn+CCF03nopvxDk9rEzoK65EezZlghTbjxFakKuLh7qx1/BQ5AXLRQG+rfalSVM
jb8X8uiRJdl2R6yZ5fXWyNM28qXQ0Sy0T32AmJ3in9pqSnPZO7mt7a2GJOgo022p
7PLiwct1jNsAJ4hYRqlx421FLgIAc6+lbQSltoHTjLS5moMNwtoy/gcyj6tiWd3W
og4ZAfqFYLRRjyBVfAJ3TsUSsr8qFJchMQzMczu8tevWUXHldk8MZOpSZE2/HvCb
zROobjgIZfS3z5lj6OrPTRW2ELMeKZH7rwgq9sJQcvNhRndOJAmRTAXvzhw6zhut
QJX8kXeawD3ZSQQSi0R14y7WtjWeJwgGXXlrNYORZuWuXIRvGshHf8tTzrWSDQaT
BxWOX3wSfCxjGWDxzin+PnqXSJQz+WCCEVC/R5/z9XubPhE1pKA865QqME96oPzP
bMzChqGVrf0RW7wRbOAuec1Ru8PGNoesMwP0EFHX626vMZRVa+6wlVG4YbHXG/Aa
p/LgnvraJJRa8lrhy0tl/96V0ILJcU2UxkEXJiRsmHYpJpsoI6CZjIJZEbMmRqAQ
loMsBxnl0uOsV+jPd+5+QHRyLatycC4R3kT/6LIXE7LGuIRuOVo1OM8U7IkaS5Hp
wmVAwQmgTEIkBgabT/J1j4M9romXNIvozvzaMA408+KnFAus/zw6QkrHssjWZ6+0
FV4xN7CZX8At6c0BOidQ6JRhXhWmBDS+tE3IxYgvdhbi58ik+kg/WoujUONqx5S4
qXNEK/0Hi+ld+tYD3lU9/i1QdLBbos441mK6JZrWROjk8l68VAvNk4qEsQ32+0Ya
KTIwc+oKMQjjZ/ZtB/uZr6nhAE9NJu7dlvkn1M9rLB5OVNBgyl102zyi37lW1ElJ
jRt93Gj2xmVAjoG+SSPOpDaFLpQdgQ2JKFtu48k1bFK9uyT2K8wTpUgx08FPRrVI
Z+F9T0AJksDqLafL9zKAhqP56OobDi/6KYmWGgGzfYyMt6Pxtml20awUCraJDJfJ
Z8ey6BknOhg7OrkVdFjb9jLizMBPn7yGAItzl7jHtAULYHQU3zgU2+6mzvmr4RUs
NJDcCp6uqEXl6aoE35xJ03VVy5Lak7fmljt4r24/YaDXOnFCGJRpDMd84c3lF9xT
Orz4q+1fyquvsVxzhpoqazPcETJaz0YrUIgC7U0WjJvZ7ofclIAlUNBNF1StZ0sN
izI+Wu0ycUZBEcN/iV/1kKaqp/UEyB9vDGmkMHw6LaRo/LGgQIzl52gqAyTPCpsj
03IMwFSTOT+VzU/hGAK/r8rNYYcQbhU4uO40kbxQsEl5win+m6DP20QsMv7RmUxC
AKO4uJCghHVH2pBwUiKewBBORyfHYZKt4psuvUxUNvsQuSqNQQFIPOIq2NJCWM3z
8b+UrAlHFlw3wtD0ag5jpj7RahtRImhAe1eyumMXcXzOZEjhBQn74zuH5nmj2cPs
ZbEnEO+T2wYnW+foTbYhPDUkeetn4y83j9whCFBCcSgT5W1ntVtHi+1NDc0knQaf
XNB2dW48j39r8CLqBq3djzEef0ldR6qODjQewvCpf4FdmHm2yThzykt68RumTl/W
R3fZcn+zlvj2gbTikA+T6coLR/NPmt+e7MiAmmM8Bnwc9Pv6/Cj/yF0bl7xhISJu
/2fc4HzZCB5q78QlxJAEPkvwfXnabG42hdGSwGgN7g3JeLYFXZvsWXzN2aM0I8f9
EEvZQ9imq6RMPcBDFQgTsb/H6QwwSGBJ8U98DDHpDaNOV7z4I9sCc8kCiI77u3RO
WHE78xAG/QzCg7CqCaFB9WEb7PdBhZiozaj4Qk8BJGB2nSNMcasvjtWB7EUMoCOn
o3syaN/Dnac0nP0/Cr2Pfvr7UMjf4FLHgJpvIrCZZKqmYwbPPhWnyuud75cr43NB
S7VpJGxmA3p8L+SbfcMYUpMvzIj2w/KL0CSXO8/wGyIhT4WUoOxVQW3jvcN5tSG4
Ly4LeMb3ZUXn9Jhkt5X+JYymT+YrQdqVGfmo+/wSfsEhy1Z4lUpA4cDMo6Mr4dR6
e7jKAKT81UpFW+ynH0m+B42aAoMeLHY2mqiOOefoNeq6XK2PetRq2NDcRMgxohjm
qAE8ejCl48hMpZ4w3+NOVY3Wjgb3aDSWZVGqe1IHk8CFWL0tXSywJsMqNihFYwNb
5zTbKp1AzU2qYmxU//H7o7G1BiWfVzMnIsnz3Mx+WGWu+xa8cdyLEH79GD5YlTsY
HYUgGG8geSWazYlgQYhJ2vxNXddLefwEHvx4lSpET4u9FcV+k2lsk24uCUnbiyQc
0wSOMuv4NFrrshZRhG8+4w9Hb8fcHIwcH4YfhPeSExW0M49vSR6uo2cS7Yv4ia2X
I41LSziq/NaB2CmlIbhFBYI1I9RyDl5fBRv8P/5v91yNuwH/K2OIh1Tg68x+1iRC
sn0lGJ2aqUh9OWFdX2X08Q7uUCgNconBfNQyykDO9om8gl96Vp0zDEl+wLYElmDR
yEVknVnXZwgeKa86Si8PQmRRWoXr/bkF2ZE+GduolvdlEd6XXjAypFZHlCuEMlK7
0m3NT4y2Fsv+0ylpYplhyV+9RBO+zttqvHt9juHaAEhwEpF72bL4QGfk0/8TrRTY
X3/q4xFquIOqTUGNXOjTJnEvwhwa05d2BUsI0OrSgYhQ0+dCf+q3yIp4YEPzQYOo
URWspA3/iQdpYj3I0pvWAiAGBtFE+lKn87NdsVKlDVN/QH0Trili8MF08kdQMDO6
JBavYE927cySHtSEG3WNwJtLIxmEFCSfOI20du7p/shNm9A7vQd+8orNydvuMDcV
7YeSH0EyVoqYYgkQAQf5XrFHElpvQF7fDnJL7OuuKhmxZctwefdhGjVaEduPRRqO
CG8ogCUNhbLXoZUbaXsxPrXM/afGKukCFGA3TKQJ57xQIAsqRzH7oThfu3b9x60R
tQPM13L+Qu4PRj/7jATndKv5cMSfzebTIM3lD84s4t8x0KCb9o53PIzoaB+zTDcq
Un5Q8CVEl7jnTXtEgYmrIzEry15S6X1RBpa8dWdDd3576idDKaow1onDLOAwkFQd
JGp0VsF51RSQyXP/4nDOyX5bGgjbKtfNH35z04LPBC1CuTDWCkjQ7+QVvIRcSE7R
0pvI+DghnfXA3DtFksCT3ydzupawk6VnXYB18TnsqEtWNX9XAz76sBVEh1kc/y+G
06WeTmXXqU0GzWzuxzzv0+mHWZopXVdO/QZYwONYk/NnvDSoC2PJk0vbIfpeXWV9
XmgMKCGwTpw7Wy+0AoJqmnSTG5KXMxEB590O1KRIAiU9gNQp4FKfxghZS3LGqtAA
kzyJtXUtVlS9LarKY5jw8ao2gw9Zn1rVd0LwWsf7XlNmCXEeoNnM2OTGJgdzFEYD
p32n3yZuqm9gac5o3KW5brO1hwreSSEcg9FOpyT/ElNKWH2vQfVSPsdAtPaAJ6V3
ybMBnxvmtXRSqXx6tC5v9VYaHHt/j96sSxVkDMh/Urxub8Xgr1cqqot+ZFgRYHYB
ZYaGWoUDiGCGhsoJzqHpEuEQkTX8qDdhal77PDA4p0fQi+2A/LU0f40vwi6HEHJI
kdLAOLn2rn0bMdiWuUsx/xF4g8CYCHpli8X9d+4opwPR1ccPxqgSGAT6zyOrn/Dh
x1wuUr0IEVa/MZlX9alrDZExC3f1XjteIE0CBXSpkT5XefDwzxodcP/Vwa6+G1IW
4c640IaVQCY9jGvdFUS4Z3eBnhIXI/CUmxQGIR1i/CDjTlobmc05OpWc3So3b+cR
K4P6yhFxA5IfkMEDcEDogAsc+RPAgg3T7Ae5QaI78IkiAp0TeZitRJQlPoqQtTTZ
r1+9bMR99iB80JykLMNJXI46cz2e8BGxiqzK6PpQ+35GJGjRQAm8xSv7iGiSqfrr
eC4xe8ciEMYW5NZ2fl0srh5xmd2BskXg7a0fngLJ7fZ2175Pb8DnifU0H003c/Ce
LATVVzRuW/6/hUn0XwkwK2nw2woOMt37nitKMvhdd6dfCrpnYC7FS9Xj2j7/83Gd
jw10PwUINdnK2y1RrE32h8KdFFb8UtFiFyeOsq16f4eSVqhoqy8Hayzk5ZE9p07T
ohFOMHgLOpmvSU7m/gGMOKBaSgCp9FCsdWOyhDOXIeu47g+Yu7U8ih2LIg77uK+R
uFNsdEdnieJrPGXGz42v9OHc8X6vJ+NSds9n+TJT9PoO2VS/6WBC3EVCcrjXv123
Ai/InFULHHikYYw53SAz0sJJxo7/ox7DPZMGbfXSQjjv3Ncb56kzAzwMjJQ04X1w
zMS8WqArKco1IF2W0Soiam8WjPnbQsd/bxjZyDpapNL2rNzv8uscP7XTnX7/08A9
1MCYmC4LKLjtzS2lOvvx39HnzEYSeYNhMKlw+0VKhboMpNQ/wYmxuMhberfMToq0
d4sllaHPv1bgUHJPBKpPXU8HYdgry10OgYv+ZPS2aJyHDKJsp7cbbuZBiyef3VDT
TRd1X+OorW6/hnx6w1PDBeDjh2xvzGkKcMmpU/y1GpT6G+QTXpzLcf+9t2ybgkPa
T6c7hkujt2ohEiBk+WC9YgyKNPk4vaawvyxGea8V+xWCjsuGEWUydS4KCDNTw0Xd
+OXhQICWmAp1TIMI0R5fpIzjqX+T9q/Jo+kDIN+hhXRm3TW5qItRM0kI4gRbPLYD
MG9QV4fOlmzsvZEw5XiGM/lmkBVVhqGbfN2kvNxsgL8+N+Om3/Y1MdsOHWNTcNtV
9tnwq5BvdKPgFfV3oUy3oD9CADwBBrcSOnZBzNHN55IEMneunVbbOgjAuTYhOnPN
PSChxeA+AeUNP1CDla+mbGGNP1w3NZxBo6MN3M7Tjx7LaUT3A4vTMWXqaKITx5bl
h4Yal77NPzT2Y762HedoqepXQAuEor6eHnocbBn3AwrwlkWz9XRcDTyGWYWyFfQ2
KHoFr1AesSdl/LjmPRyVT+T4CIVGXWVNqOy+IZdDNng5cRfEnRVBX3uqy/CjfXH6
iDczyL6D+RNusHGdEYx7CHo4Q99G8IaERgutBeB6UNv3+fBOv4E1rhkaHnlwm/x9
FoYSlCmsQCK2o7yA9CFF4nGQ11AOxnCHUNMHCSoSlklaJANEEwPBXdnhNz6AkDt1
ydv73kfkBWkKrxZNGF4YFdp+UNwg3j1rSP4m4MupWHPm+5+UWYP4t8hhSzzpkYIi
nfFf1VCnUZCoiLQaKZL3VVL5L5fzumXa3PLX0PuhdBL8cEcJXmPv0KDIjfa0Wzal
QvRjBs/J7FSpFDs1qMe/M1u7pdgqGg//ko+WT+gESUdsR0sU2ockprNUaY9PPLl2
1kto8EjbR8l1gskXW/1QVMrz7jT7WShQhkMJ2FxUXswIT6q6hOqo7SD0l7zIDqYA
TQLknfRkPMDq+GjqFDLzfs9wxya0s0lw883USY1B7P0Smq3fJxBS0CNG4hAT6jZ3
lxM9vTCaCLg4M6ldlI04K4/aodYaOda2YkNoaoDYA2asywmMLdAGAXhZXdklfhUO
VZVoX4yVd3RW9VzzSGGJXjTpkbC6kfOQrwjAtOa4QceOV+/xW/VAXLZdw9MpaYHA
AJdO5rvBqGfRhS/lb0sk5Dr+J9+sxGuVt0hUiFYiotMFXpQHEEOgMcf4omjbSCr4
OIRg/ATaVcCMIiX9hCZnDjRUjpvB/WG8+aFeAR2JjAPit1maBLAB/IwpL8ioyu13
vdxN01i0XktZHsduxpfrvb3IzfMCydFR5J/sCxtJuQb9PvKo+61jEr11RHzKcJ6E
H7ixcKZ14tSWoPK/LZQScKj+FKjChPZzgZjqF+mUr2h4EGr4cOZNPaNeY8vgjrte
XtoSlNe2p3+Pk039lIu0FIkZnnLKNS3BYXn4VCWBXHfK3XcqbbwjlZ7cFZDuzxWK
488OioiP9Uc4LcPFae2lPed/7JHufqEPFqi0/fy1VXwTyXSGFwghtC4aHSpCF9f3
olMZ9qsdzT/MUqBFtuQG0DVAC98V0hXDPFpsMDTzGkd3MQaP9jAfqur10XmCtTg3
mo1opb9Gs+7sjEmSRsBmPVrAgc992Xz/Di2xHUjrDEHyBeZAelVz0gCq8/hglkMk
HWcf17El89pQLPYJmiqeFY4izI8785kBiDp0pjNrpjiGhZavEX3aBZ/KGGMGQ1Ci
oOB8TsgWChc1XSbufENdbKI9igCHzyJmRDUecjJEJOzmQd/DwFjsgWXxHIzuZfJV
E1Dz2UrmPfblzkmTZDkrltyvR8Ts0748qKAecN5dE44tv8JCDJR/RznI5V297+fI
yM6O0mLjZnZBMvUWy/NZHvSYYd3a4lrpZTo60wvNBSfm/sBg6oYptskd4RNDhcFf
YKMwsG3DCyZoT2NlBqe8Co0/g7+uvbjnfGB9KhVpFJY0daDvKUHBxfI5P9MzFfN1
QfFvvpH52nSGjjfVqvaFVOJgbuQ4Yk1Ggk1mb0rR0prrUvOB3BElGKNOKW+HzXsE
hTNLZoQjJ6uzK9tWpREX4YWKKVfB9oP6ZhWRrnnJFrfx7FI1qsqZmCEI8l2G5hXP
5oEJMLD6ETqzW9SXRp16DXb+y/GeReSTtgBDuVi6oEoxQ1rktpPwl+BvTzQ866dr
aYU0IUeQe2tf8g7eFka5KUAMTFehrz5Nq3TcYr6rO6CgrBUXiWL4i6XyzFz18lCH
fMwszlHAGvtp3LCAz9YMJEhc0NscxgZlehXAGtrrKkB4LqvYiI0pyjW26dsvL7Vo
HuHvNm1+8n+UlNqCwA9e73eExFjDFB3A2YU6AwiZGseKR4BUlUA6G5DpHy/Up0G3
oDTp/gFeFL7+0hroV8+kkE+WWMdOG9GjISf3EwCMoAlXvtVQaMm4CmFOpKS/wu5J
wRp9v3IuSRTeJ0u7Hf4SDQWHNPmY8HrBbnU5MxS03QzkKFfoGNldRXGZLfs99fFL
RMxkqZO7NTOgrzuPW1kU83eXzLIAIIGOz5uk7Ty69Ms4S6KMND8bKgrsw2KiOEDL
yTGpHHMvkh8qHhGgUgkja4LGNtTWHrwsvR+o3DfFBcTJT/rRyg1NgGFU4jzfvB05
3MN6y6z/v+fu2ii7Vd1D545emAd7krXSGyDw+COzAL2axC6OjOWHOn7TH48nNxKd
PPkCiWxls+eYSLYPmyrJ/rju8jzYyUNEvLFeHl1nTggqlD9htLYp1nQAqC9+epd/
l5kSQ414Jd8vkKfW/SQEh6V2G9Hu41pBl2HS9EPsfGfVNs7oQgCABLw8R5qpPMhF
HyIVtrQweEVGVmAQOGtSxOG3UfrV9x9vtm1YOSHbawjvtzFwI7oIMmCrtAWXlfj+
rVz0uqoCoEx1Uw1KEgDwc+v+ZBKTkMb3uUkSsmDJQRiNS0a7inIBroFP0CHcJzhN
oh/L6EIhGR8iXLQfgvXbCZmHTjY15Wp7fQchSQZiQG35qMqFyiP36qThgCNS1tBK
DXTZiSlLbT6dwo3HbK1s6dBB5EEXx+wBJIazVPzilEH5NKZxjkZAtMK75gkI5j35
k1ztQbrueY6VYsbPjxOlD5e50x+p8Ux8eOtS++MzVT4hvtoKalfWkUhzPmX7+uIx
U+PHJf1gGyctE5BfMBxGSlcVKiuhUXngGBiFUP+OgdxG/fRi35VW+j7up3YkhD/q
N1wjZJukxCwtdtRVTpXApREi4VDzVtHW8oLbusTmn2auhyeYzPf7cmozJb/owFXf
anzC683HCbOmjmgz4l0/NLh/DhjXLsKBDX2o7kE2WbTYF4gCEcfCTzJr075v6kQd
Xvg4HMuvjnV8LDbT3E8SJWjeuFTYmoaJ1B+4wQlZ0z0dRQYvw0jGjBpZ9ua312Qu
QRBc2EU8UPKnosdk31j0yM1enTDiiJT2ndYrW9EWZo/QS8nTv1Qde+fPFWLJye89
DgfXxWw8nEEVdjP8SiFYDWUw0CvCEAnHiDOPNZnm5TFqwyn2KOz9N2nJWh31IYg6
Vjw+DkO4BfNPARqWfECkLIZo3Fo7q7hfIzAkltaQ6DtrdblwsS5ro81CgCzGCVTa
G8VY8ov2TLFy2Y/aPZlckpTnS4rliCDZBDmqS9aCicrLkyMxKOAfkCRzZEoidXUn
eFJPvc8NuGCI2O9deWA9zTuS7vZWVOnBR9IldEnm74RTJJYsWWKmKHSops+Loa3/
ShgR/iTW11dTK+BlaC6B5wu2cgPvzfqJxubGhyzJ/3mOOEnvmpFH70bYs5YRghlg
V9vJE/70/UcyU5vS98bhXQE2N4m6Ngqbh4M9V4aJ61ZOWjFKQ/O3aslwi/qTqZv4
azMPu4K47UdZ6P//26ceVfa2NsiMIxA06K2/ED8UANsS1MJj2wiTOautY4m/5yE5
2wx220tUyPsxko4cAcMkJjJzBDS7JfEnTL93Ck1WpRKwCG5S+PSRNiNE0MOu2Bup
Ey8klfI99oDjQJ4Xm5V/DIPqMuKbDe3ZpXxqswTaV8azRa/h/zd6EsCjazkKJNhc
VP4J61d9vSbfu12REHVoiXrSPZp5JRozyWTsqFiqEXUueDSZrLr75OfKZpyUc5Nb
udL8z+6EJvBgr2hoLzha2qAnQEzOiuwW4b2IYDVLo/vZH+RuulY3l9lZdyy5UKAx
pnZSqRjOgtULyU7qZ1bXNOEHCEPiM3/Yy+0Rv+x9VjkWe4rv/iYSGzkfTTYJaAsr
fHw2SoTrRz8TVQLbtRdzfeeyCy7WCR+TfchV5FD/NokIgcqaOQJBa9qBJHjWDyYv
BahTleWmG4lo1AjSl1kStrLIZ92nC4tb3XQj7aSoe3Q6z22WP87ER8xmrK7reBlU
8nQJd2Zcxy3PUQERc4vDCbGFlbG5giy03yqRo3nlG0Y4Id/yePNs7liwRDpBePbK
ehHGcQ1t3zjp/xtpXafrLd8fLC99rLCICC7wWebKKQoX7eNO+npmEkr3w72iqIa+
73k91ETXJe8MRP9XTc3Z6TCYDAafRdL0dWOCdqFmDJQpbokZIe4Rt94p+v4CK38y
S7W+D8eapvobgYraaQfLWfx8R2/VyDH7no5zjA58LkKT2bPFZORpUPAdnq3LjPa5
ZjXVNoH4/bUrJFgclHKfpDjd5b3d3BCe3snO5RlGxyRx1CXjSgagpzmUxc/dWNyh
I2QNnyi63Nr+IP5lEn1oTUlx5XiTfm2BeGICp5oLSPSrT5eG43rD8mVjs+HJxCTA
CmQBn5p8p/9X4gGfdJYdzWtfaWn3LSIADwgKC/ipr15l5wRwfr2qAC4wYmI7N7W0
pY5S0iBSnICxHdCygwsVkP2HdcnJnLmf0sg6sxd1h6WGnlgiMIfIi9txUA0rVZF0
o1GT43vMby7UQasnkz5ZojxRXYMdTgud264w2aJVen8SXZQuZtZN0mZJFo1NFI8/
W6JPS0R9CX+bfP5954mmQ9DwiXFnW2MuPKLYTzmbIqcgEWUKsAng9M8nb3r5YcG0
tPaJM0N1RnQRr6cdwb/2GF9JVMJ9s7cBT+fsN6h0UbuMqEh+G2t+/IC/rJPU+0NO
tS8do6mYnLQaUtQ+BUeYfxRdxE0ofd8kGEQaI+6fnLWg+xzWXx4fxyKH5lqhDFA4
jCA4lP4BQIxqzj/VvGM+TLOLCNljNngPn+2LjcL7cNpASSmcSy0a6+ATa1IfI5ZD
TYhgHqFHxLtzpFHOvOfFlpvJu8+Vkpf1oIIyJHXSS8EFozld4zGe0xFzSzHOL+/m
O+jo4Y6CFd+UHBObSmgAybZOI9fWCYEARq0b8vR8j8FOSAg08qNQsQ6hf/WKOG4J
Rl1rJZnBrplYCFdsfUhQMBxTs8SqGnc1DH6l3f1Sr4UWfpImrq2ChD6KPfIrfhoS
9bPbikY6/3QPTU2FaOtKEmvT6oEenvDFyoRFRPvfrrjMp7n0nH8hP7Je//VBKHgW
DcjsuzS6+/nkXggLzVxdma708yffj9wwaDC5UCgUghSRUCVItrEX7ndehcvi9L8T
GJsQKUQvD1NIAskDTYoE14PJgomb9Y48xTrkwsCJyEIfHrt21mMjPItQt9V/sQfJ
vUUUfGesQvOSizugvU/iIUoPNDT4S642y22heitHfCrcVwT0WqcaxvsGNYdWEScH
UFW+XOamuXh1qmBTPV7AIk9WRAbLjyxqrar7EIN1paUlb3abQUzlCdWPdpLU8nYM
cL37Nvrl/H5HqzRPBRmuHjCrGsLIhXeeXqDPY8qGgEmOmIz/RcwBCpFsT4xnJm3o
x+bXirh/kR6ds2JLvSx51EPGjh8gtfM4bu5LqGgsRz4B+wgN7myLV+38nBl6fJmF
O/aCa4fHucDcov2zERpDogV/1RtzrjwjGGt2qV3Y6x+dpbRjTETFkzE3Npn559FQ
+Why+aSZjVuB17IRBuKREadZI5/pCmS42mvZRNt0xcMKN+vtaPUwr76Wzeu//pYa
ZH2OoDW5hX4KKbMFSjUAB2w0/co/4a3uxEoA5jr5v+0cKkAHxhcEg5P7JGozvf9q
IJgLdkOOsdbD0cS2dr/kDYEXYLY/hsyIry7g5g18j+qGux9h+G7DtuFcuruHAAVP
ggG3QrdRP7HvDUdxtDmBV2GrgMl/Qzhtfk/t/QSt04lGJUjbFIU8lXmnPj3b5hbQ
QSn5LnrNLy2zFOYCd1h8vcIaZnBequcl7qP484YGXlDvhWYaa9448stJEFUmwFby
YqPErWXP73+RjWKdTm9DgBSuZvsj9N/tguak+nDOiJMBvTUynBOKhNMthLrKci6R
1sUel+MptOVSmLutM+aFzs4e2kZzJbJNMnV88e2SBFGM83Fp3l7v6KzEsLBg5EU+
Ol76jBPupbuDjajvkzCGJL+Nao5E9GnPFK2iS8TjN5rHeXr7pzMzd2F8oVjel7pX
Pl0Phi/Eq9kThzaAoYfxmQkHCSeA7ugo0ie1gYiEGaU9/flQqNXrN4ZyM9Z+Rjja
yP2NOCxC5VT8xLyEeF8fkJ5anQFKr1pRML2lazit+6rY3BX1L6hB5hbJeQxlmUM/
QDOxxE6yWnXE6TrN3Lhik/J+j3ggy8zeKFyV/cn2fEZhIoZQ//hY79vt2V7ICUa3
AhAR0iym4p6WF5AtGURil99bo8SB81pG1LnAV8ZyZcfN8kLjT1QRcaQ+sibCMBlc
TrF18ye/ixaNFDnIR5O4TW09G1UG6lECX3R0lDbiXTJszAfHytJfJ7X75w1u5Xo7
a3sTC8bs5VPYUwAiBksxYdCDm3/H00c3zTk9G8XYgGMbkhc3bMkH3ZidVbKJMTnS
fa7Bn5Vijaczo1K4HyIydUDMXXHPNTi+/PVqqLRKVeSomr/OpDm0NetNoNv6E8zy
J0g5r0Qqd3jeW7IZQW+/c6zz1pbP8FRPMUbSbLa1+r+qACAeE192TYg/5u3KRSA1
shOwrKhITein7yL2jJ0L4nSMCXlZzJtbWQLTfdHdZlLy1G4G8AqXVh3pc32A4rxA
+qTyB77KvPNCGiYWn/v8ke2enJIt1WMf1tKjGKJBqa1V5p0k/xhpAvxd2pTIseTa
YhVS0mtwMAIOcsqr1gOVuNmoU+3B/7VloJmsG7udeIcgZk2VI1CIITP/f8n/4log
1zoCvUPzzWzfW9JVl1IRduistuQ9VNOgAV8uaKK558uZg+Jql8DARn9ENo1ijbqv
x0rO5UZvhxgq5Cq83WZH1D18yXZWWrOyqEJW9bj5/IfIEma4SEtzbSoOharlQe1y
8xP/oM7GbIGji+z56RAY4oeXXfzPZ5q0cNgL+bLZKVfXdhe0cMX62Mgn0BAQI4VV
cSd7bnxz73gz4hRAXB7e4NSKfgVtyOYhVVrWhujTEIkGJtBjOVObIVaIESNyzRFa
lmrbmTUi3sN4EHh1DVKzArX9EWYqzYyQJh3mkG4J0NlbOqCpLI7aRymPR+MkjiC7
loq6M/9/PgDLeQQBKPoaudjzUr7W1XOcfMI8acfX5QU5C7kzGRscVgEnNs1pXCSc
VB10kHgK+NDKId/gdls30nW3S3JB6mIF4GpCkWnB9Pzw5bZemeZfdDtPzWcuVBbJ
vDWTZP8yAMHHD4TKWnxOg6OIQqPotSQEne26YLoj4EMGQ1vTw6Xva0TxPmhrissO
KdZBd2Eu0GLEO2o3PFVpNFAVPYtcz3DnRy679gOJ5aw8ZoGDpL82w3od1jDId+i2
fM6Asuuws1bEy1ervvF2EgtQych3L5tc5rm79uhVkFoQXBKwSHRPVtxD15I1sSg4
V1tqRA/i1pcpumWtZQRg74dpwCimjCT7BPA66SipBCkePWz7BILAHZVYG42YYIyF
tpvme9Qgq2ZwSdXrW/UrW0aDtsCYbJq59CY4+kuHeuM4+xK6X3E3yYLIYadsP5jo
b2ddtx4ddlobWOAxsON5g7s7/3TBWxO6RLVyTk8pQ40jO5k8p37YJ0pLtd23bYbT
mj1gXOeBJ8fCkzY9mBOpuMxJPjTmpR46HiaRNorq/FWxue6piUNnrQ1IUN4twgR1
WHAlAMdNZ44x2FHLj/lU8qXCwkSR5XxMUV74hlNPO986HMGiGrvGfwTCIz3IjTCS
TfOa8vT483OQfdrze8vEVNPf4U6EQ9jJ2Fy0jNiIP3cRhDww5rj9654URPqp3fCW
KQ0R53/i9TaOhZYz9kVCWawB1T+vLSXxm1vIqXmP6yFcz6i7OLQ4vFjBhFstVG8p
u3cejdOZK8NHlK17n9GUrp+tDUQrczqMZIwUJBSPLYpyKv07C8mCe3M9k66oz27e
Sp+BsWmKasMWIv4IupKM81WgqN2osEnKUvftTatK33vBgsyDdeM3Cw4zk4g3DYMJ
UlFTS6cw8uVAV7OSXsnuaODE71BKA3yFIGnmIffXaHAHOd9kBCcIWe7zeVJlk8oX
jOsWIUUSChY0a+roqS0DDZ4GVtuXYbTqrpCiTCvMVpMw1pvpZLe4niAq6MovH9hS
21tpj0s5iDC0QJK5Z+Bibnjh9MG7nxhzzg2hRBeLq2K/7lXOLaB+hV99ejgIk5o8
bagaTMPqCEMtLwu15GBuvv1j+F8zUwBsy5L1u6ZmXPykfvDeffaR8PM1Ax3+jFMX
NDgaEh1qVUrSsepo0RCYAnlE7CFSz6G7n9bYYmqnZ/hYQV4eOZ+42JCXMZAKFZkA
1/zoVCax7SNARP3zdXRwcsTPPdIjBByTqTN+DoELYwPr6HXc5xPDjK3bGp6m/IIy
nkb/IC1Myo4oKupvB0nG81nXIb1DDsgcWWSyZvXySIKUw17Brhj52sVSRyDDtXdi
9Mrnx9q4DAk2HNFJkrhiaFsW3ZxkNEI7sS7W6ZsOSSrb//GSOxxshM80b55wxyeW
HuXLF/1o4ZsDIxwsxXEp5QIKBaoAanthyAYOJc9dw77UpcRfHmQj1f7buqzzIA1+
nrVjgWvak/T8UUxXxav0KcrJekBgNjImEO4/xjRAQwQ+RL4zO2i+FnZuF8KYuKdT
1Lxn/ZbfT4lWoYq9l0S5KUYf/9H8HkoxrUtXNVxxcQpMNNftY5Ok9h+q0HiRpuz0
wECpn6V8TSkLHsRUenyOcpDufTJjYn1kKJRcCqmKWMS7nOVCzT6yj2WQLTECOWM4
MdvOBxRwUg5D3ODlxBpTEsW0mpN3CDMlZN70KA9qCgLxa8qjmMW7T84NPyy9e5i9
JEOZ2IpqoYar04Heue5deNYVnDPE5K4/QHSGRDLV4HANL4ZwdGJW9qj0CfDS5Nqi
OM/hZ33vhm04rTD8Tf/+lD/e0DmyjvONxgVYNV+mSRADAgStIcjcplx9I7n9Ynsg
vd4cBzZBH8VWEMTTC1QVMd8f6KLo48NiFmsJLKsislKWA2Pa6z22frGgs7Ax12gb
iA35Obl9w9F4DgAGQV2iPfTn6vFUUr+xB60Oe1E+MyV4A/39m/gIDLgrsChHoGpv
YjXs3TAjDzsR9xQiAt8zJapDEb0ffdTYdpqswXiTsp+i3ViYJ3YWsMhpeDa77LEt
flJWm6kSmcojkIbCLRiRW0ezjliF4j8NG5otIXXHOZf7/9JPEf2NuL2dj/vS+ww3
C6jiudFAlq4oMJZ6lB5YMAFyU42hligcXATKOKuS3BhtI2XLR5DRwYUD/TwtcaRI
ROT/dOgaTIiNUWPSbkBtqABNMFXG6aLRtMVAcWYNVtxZvgClKatht3AcJfQ+UwgX
fNCU0NF9PBCpOErycHZ3jrGjHRRx7Py6uQb+R+6X9kn4lr6B1uyZiNADVuUSf43H
ElHDEQ3DP43GzYLqo2pCMmmKwI8Um9Zn27PUmErCRJqLnNJXBlL1IIFrMm3JWHIC
jL02s74bq0hjo4w8Xy8G5BoEKZhPQKU1FSDCdRVHbJg71l7VRAeX7aQRbk/Q9416
UeA1c8enY9QfJWVweO4A4wu4cpnCJCIWuMfAWt+A3B+rxxKfI9TGH2LmWLtz//Kh
vbepH8qUpdPoUUOLInPtqw4OZToqkjG8hvzOqJtchoVubKZtVVv14FlIRtu+ldhr
u4/mg5uW6nIT0kCx61uApVtQLOjLtgTnNetS/6+7N6sK1mi3LBUJG9CcaUEZlA16
4FUfhOas1/M4dh+G/RXyrolbKaS32A8JSgzO0goTtOxr5iVAqC4JqLT3XK7qb3NH
Igfy1LUzlDePNymj7W4+nqkfH8/t10sE6iUzI//hrHxXcdNukbqiuERn4qiNuqVJ
3eGGTuNhFe/BfoDTPmmN+YcZ/RIU3KOMor+8eGnurgXKnRx2dY5B0HB2cMu8VzDN
kAiCEZy7tBo5qF2arePONJgRcu4Oyf9yHSUhG148jCApYxDiOXNzJ8w7Da+3jQEW
Nn+D/IuEQjZOArNTE3w57ASDnzUIQnnpInNZhK8Xs2C+8jGR+GKrAd9exK+zceO1
CMTZrbXHyBQfF6xgbiDCpU+JTPxdzZqCg39BmouDuarpOc/DpnB/9cuy0wTNrBOb
6bNIJgnnT+/wB7jkyue/tCAxFJb1Jg/J6YJ6WiKpBQFkzDDeIp8AVIag4BjFdcJi
YPM3prHdSg0JUzos84s6SXSrfxnJtfNYXtjCQVzaofjFJ1sdW+YyN5YhdN60n+SR
/XxYHAvL+6uRHOydV4YAtEPEJ/OiVvaHmJBFEzPBifBpWHeT861KWv3Jz/+orJmI
OlwOocIkk4VqqaVTedFQcFB9HQq/3V0Du3k41JdmNlz11Ubny8R6QC0AtMwXL+aO
0q0qY3yecCZi1qu64uw5Fv2bI8nargojUjE7k+mKouvt4wrhvFuk7ccFll86debi
ie5LR6jLqWRX5D9pZ/VbW1+StuQU44fE3yfuO5bw7CspNTu/dpTcBmTSiqU1sUl9
/9yfOHN0WJebUDdBKKfDoTTkvAX+kdYjcuPVvvxxR01OHE8DvvezezidpDKUFeou
Yuh0SILLlHb4UnHcDsbh56DULseE8UFePjF8J/P6yCmV5OfZyHpUC9GxaeXhPUzc
7xHGjVIJpY6nS7HICQJHeEjMtIWm+qPWio1LQqU5+tqBzx/lcj0wFL82BFx+G6yk
DOBsIoURHMKCw1lrhS3R57iYTpX7WdgpRMm5o37O3nIR2K4OgmMaJtYm2oG5cJJn
PJnEkGm6iXddZ1uZLaO/iRKXG6i18UATD5LAR/DFLYagfLojwCroHFdAxbmtEeHr
6J3Vu8iGN00PgJiCppIpa73sZxlIrp5fwo3AxOTAtMdj5fTKXonTZ9UCmPkyofA0
Crh00tsTQD132Um1UJd/qSMZB8ZkEoEbR69Bq+3QYLAYl+nIcX7iISjK6yFRdIeF
EiT8Rgsj+Mk/rOUtWRJd2HSLL2Lah+1FrEds54+EHIt0smTv1J3iN/PVrqpa3eRp
vASFC//Tw6+2P7fiS7KgkWebc1qr4KkydhIBZh/K6eGAqiOXbUm15rOzudpOuetj
rnygbxz5Hbp6HsJ0kTQi7r5LjSspGrOccUbIQc9Zk4Bk16B/etaj/f5pxOwtToNr
xKh1VPmh3PLfWP8A7efd/fMGEwb5N86xie1vcpiMawFVqqqlFfwYEzxXCUvSEZHH
MdoLJJgLswalhK81HNtY8EA2iz2+6u/EAK9i3golijqDyqbmeZthsJijeaxWN+28
twVTNmvnM/Iy6Vhaz8piewBHqVyFMi0WjXl1++GgW2GD8uFfvlMFGk2Tb99/5o0c
TaKM1M/tokeLHVnRwfx3BwsnAkjdPNgR1R/6cLQhcO35W6uwBrQndWWqusJ8qT4T
GQ6K9eJIbc5uKDfZMBAmc07zpP23WRJxb4KOTcouo9kcUQBXSHpAX9iC9pDmqFe5
k0RyOig6TMfwA/92Z83coAEijscFvNbP4V0FVks/n54GkoH5HRCl+17Lm6f4cST5
HFWEqSohg/FSHTWbsQg6+QnGF3O+NID1HxpNrY4YxkkIo4P+zFNfkZUpIg4dybtF
iOAfBACTv2X6TYw+HV4/evOe+52+UeT8PJOSmDumk7Wo3OYPU4Ut4uu6AEEBzPo3
Fn+Q2sYIz6+nNEVBXosfnqI1qqW8FXoOO2oebccRXCp3PPdWAtOVue8HS359Chr6
YvzfcXo7gXv2GP3Y5t3S7fryF4usgtx2TVLdsUGPVVzqEynJ257kk+6wyqOqRG9Q
RaFf0x5cfRoUXfcE5WsiDDeXn9KlllYGog+6s7W1qi9vim+qNEWAtNRmZDHbbpFH
Hq753T6DtTVt2s3J+QhlhlqP0P0MoA5oHt4Fpz0HaarcEdS4D9V80/3kK1uJltpc
djA2zGqIwOklM+OamSRq9e39DL3PUzp0x9rfDlaOg7qUssf72wjDvFTCY3oNWMts
gRPW453b4vF6j8HuMFflE8POn3ChsNjxA4MVOg5T4RmIWKMSmSGIM+eErG9ndmiU
zvDM0S3O4zGhmjrmMvBdT7wAcqD0PtdPZ9r3gC36ta5q+eE2JpJUZ6Jk0n91K//s
Nj+W5eWFaTK7PRnzPg2sVUawPU4ERnAH9tSyj9kFglVN2iyVKJz22e9/nujgqOah
uLobUiWi9+KYu0BatiR2tIDaNPZ2yYnZVnCoLx/P3T6MBb4M04XJFtJcWqXzNCeU
b6HEpabMMPxVsYFRkDUcYNyng3N9Zk2dDvwElUr7gsPB7l+XfziFFaR7gluO7vAk
h0owu4pOB+HC+J031finurSU8jRwA9vnJvErCwPr4nwKpJzdf/OLD7O1AVgLD5a2
Je53AiPl0N1LCCixoegaIr297sm5PZVhell6FhmsuKwjKzQ3YsPR6XvzXV6+fccA
3hzbPPLDvMFpkmAViDQM4aaDiaktZm52+GhpVKX67rlsWrwgaQkj3JryCc8gPaYS
ms2WKqInDd26Z4Rj0v8a6cag1jFU/+ki3rcLuYt8WCMa/C2Ww889GbSZL3zgJqoj
/pJ9rEUb8EM9KiPwEErZocgyzBJ1lrHlG+s8iS4scRQwx5BYX/nQba1tQnTRVAUM
GW4IpufPwSGAgSj/qkH8/5BgmLU3vVpIxCD3V5BvBxsG0bPAuafM19RW3Pd4i4s9
M7KdEfe8t4aQDmiammIFnrCfSojlq64xYxxtndXGYhxXeKnvfzvmWf+5GjuOEotC
H4Hde5n50Sy52Qr4JOz8fKdaA2PzKEPrQk9mxBLafV6bGjUbIlFZVdaE3QbD6OJX
vuFfxTcmuJOr40UoV6N3gPexeZUQCnorcfJCDz0lreL/emqiI4LRIul5+At9+gzR
xmppufHynVildYfbq9GZvnhDEPBgvR9SlYScNRtOVk2ZI1iZfbRywr81MLuvgIu9
WdPdmov0sQn6bJoRDijZ7VP7JDk2PjIuRmyyL5KKcAD83QN0qKzks+9SXlHqPV5l
rxCOkG60t0jxPYJGRDTkQayRWvlH1AFcinYbtI276DNKMsP4/46kYZTYhxBHdwjI
PnH6gQInVAcjVlQc43PTn5LxsneJX4dU1MikbT3gpj/m1fX4sxHjzZy5RyI8CgWv
QRlagNmldmxNyNjmivb3RansB4U8sH2Qo4jVwr82kKyxhwXVlBdLSrB4g4s2XKa2
fRROvgTsLuMov9yecwAFk18whmMsTz/yN08OipcTRL073BMA+iTcsY2EJzPKNY2e
6DLzAmgH5+ZYGCDo/Ik6wlJe1AADq4ecfcuL8rL1UAGSlbALHgLQjtA7QccAnSn7
FfqCFaCUmBE0FgyKz09uJEV+6qR+lSjCVkB6aMG2Pn82YoeC40TqLTrQbCpbgp5V
PLucu+3UQPpIbsca9AvhYzY2EG0eCHa/t3cChDKxBoJb7dUhA46eFEbN/BF544wC
gPwWFL9v/YVVMG/snTR7n8F4gZK2jqgogM9swNI/e7mvBez/a8MHW/+jtnx2hWE7
UP5cTQXpl9t9ZTlquMxmLQ00UXuqCl90sAxHuSbC9P+JiK+beyhWrCiPLPBF2U3K
1GavzKYst+yFRgEt5112SgSqde0SL59Ef7Py5QN25WwVQKrMf/eN/aZSWDVjPM7m
bfpeTX3WWqptYv/h+SSCjftpWse6YKbUOfSRfr0keZQaGBHxdVyCuiTmD0kwbZYf
S8Ni9zexReM/v9lPc8iNvtMt+CjOeVitjXMMN17fPvNqIMNuh1/MIoKHWsxqvNQz
RKjYUmC0cfYbIEogP74Vgqm6OG9Hgfgd9sWWZOAJrurmGO2d4vXq5c4ZwJnb7T1s
pupik6OyO/nKdNr9flKLQAy6D38KUk+TebvAN8eTcOVWchRk3L0Fz2Gy6gwn4Rwr
hYq4tmZb9o0nKiQKv79sF7VEppdp74dKMjEzUOJUL9X0UsIxPE8mmt5Rk2JPUL8q
ue2Jj999o0Pl6jXElk6EcaXiL+WBfTGMgGA/5uAqSa9WEudHy0eVUx3epyIcapY+
RX2zmGMSC/cl5mPxnM7i7LGx+q5MSOMf9NDd9ccQoXKJ0/GXr74UHD2z9M0E/0Ie
Q+z5ndDt7iLiwznM+iYoKy+niNVpty2N+LOAZDJIYCJ4wOCtVLar3XeTiQdpfDHY
34xdeSUiNIZ/6xeQmEIg0D0VyiqHyosqSFC4U+SkPjS7/cmE9kLuSuiDaYdybk8t
sYpOPwn11BJ2k7n1BJpIehrQ3iBgPtt2oewgrXjFA/qdZg/8hce93MfspiElr+JD
J1NonsXu4he7/RDgqio9mmnD13yt/VvW1ZrZvVpRZOKmzHvm5vCWdeZiTqvKxKMs
znsuH2fOvLd1RUbfL8mvwQ66QuouIAjTR9Vtagy3oDnGkHhoGw8GbzWSqurTcHxQ
btXe2JNddWp2mTOHfooKdqTNsDIIhPPG7Zt5RwiGrGF9Y+UNkGANCYRYxY6qE/Cm
O2G0CDUWPAbtcbiAd1xzbmVj4SQduR3N8t4jn9HzXGym8Kfq9Xc5UtxI3gVa1gox
r8PQ/AQuAzW4WHYtoKheueWAWxL3f4uK61d6kcm1jc3hJnLDayIHuAq0kUk7zm3f
JTzMXp4RXYumBf6PfhAk9eEAwKqcxYxSyag7WO5mLJIS8ZuTSuq11L+3WGyidSbd
QeGm5a+xCYasWBvL0F8qNnTPfhq8UN4GAT55bWxVnsB49aztBxuUTwJ1dD2nDYaP
ceyeSJnaNcEZ8kO+iyfgZz7pWnEuTQXLViXM3ze9UU/NJR2LF+C9OCdCvIF4kGK1
2TjDAJQ3HRp6RF815ekmniRCh1QdjmtoawJaTH6MpdOIuGak+JjGy7eimBCBLLI+
6dx8pMIw+G2MuhS2RAK1fDbasNgVJuEY4EKqIZWQFYFPOKvOA9KFrj+j6p3qOs0w
iEKuVN93flT0VWfbGD1yxtrTlEYYI92/kMU6/rVupcQkliYUdcv7UG6Rr6Kpda9s
afuThWM3zugxQ0TZvQ+3NhuwLVlsE1TyEZk2Y34fZLOBXx19lumpsZ/JM9QEmAh6
qmJJFcvCEUfNf06JKeVszolYxP2F7zDwNcwP82vNowqZDb3VVHC73HM50UR/spkA
G+l70xM01pdd8792luvzQjcr0sizJLTWgqYbAchMynlOEIQSPjJWke3+I9rxL99o
pOrpgYz9NnnUsFdI4YIF5eT3KIi3EACuwd//AVktSuqrzHgJ9sA8TmeBOvviKRxp
2GuTv5Ya+8ihbrCVJiUPCdJBjnxRY3Zfda1KYj1iiBVROAJATIqIHSETxt1Qhifj
sAROaxJQmALzLmfGWJjQtOlJBWTm5/EJkc1J0pV0BR2j00sCrxTowV+pQdGD7D8a
5MDKv1RpJ8mZq181abivFI2RgQIZH2EfHTV7P3ARNy+2hCtAkDGq2GCf+U86ZBfU
Lp7Hr4Ccx5US218iOJ9PMswEt14svbaGrTb13eZ2AAO/b2rKywH7JK3JZzAAupnu
jIPYTiM+leO2fZd8xftBFVDpBtzbpfi44xLNlVSIR5Y3gxSWmXfVWwTice4ZVSCC
x9etPuWVF8Vpycan5T8qo8AwrGCLV0/QJep0/DEovSx+RqKl4c526gYkKGbWYT2r
bJUZ2GBvSAYCR5KDukowfcJvfD/PsSU90FrP3+tAdvXiHxWfw6KT1FHK+Gzbp4Eq
BF+gF+a06fyapsF6N0eAr0odIkK0VmeEDjypOiFYPiXzL0XZvgB5x/ffZWOm9lHp
LFpGPx1Z0SlFXAfIlHz0cXpohC91giUTOEOJI/K3tdhaiA6hH64yoj5zrqwK2KxE
sVTcFsg1nY6qWgalIGykSuXZhp/LugloO7eDWLokOeJcWLa0WlxJA8i0F+s/ogMb
7izHBX1h5nK/uYHsfflM64RXiPLCOqmRi7r2h24+jtGPcMsqJRJePerppFfzj8bF
G7z9M6b9vmEqyrzIKJve+AO8KyfBAYkzx+aHnDdukwxdXrSMcGsjn7rwor0Y9r3i
9V+Khm+L+p0YdV/Vm7xgY/6NHllCQlvwWuPmLyUwjfktcwqGq0/9pprZh7Ngaa6j
1WpBuHvSB6Rijt2g4J8rmzjuii5knBHr6241lMOqzuiT0Izrq/nMAkqukLTmxOT7
rPJdhZnK1+ixEhWl2CW6fF7W2yjp8hCoXOAyGXbUxywhr4SuCfVeO5avat3qFwvH
FyEgfxcxritYOg5mfnjKEEtX6mOhfl4gn7DOTnFhwKu4w0aX5ebYOeWkd30c8STf
5VZkt5umtqoAsz0cWiN7ptw85tIfg3l9Vods190Dva+xpW60C8QUdoXY7CUkEes4
HqsqHweeSuF7+j9mJA8hlDB68eK0b7UK2Ix5JlGR+gpkMSFXGbBDv7nqm1hTcKLv
PzI/Eewb5qS+T0BLP3jOJap6+WrfR7gAssrN1jdekWc+hkXjfGGKIG1VFqM+DftZ
SJqWx4ltjS6BjvxEenFalre9WjWSGoY9KC6v8n6IsiT2HI06YO6ZUdTbcVwA1TIS
EerMOTWTWNFxuLfIFLZAHE6zoZngflTjNl5PZyR5PjJ0rwf54BBZfprjil8JRIYq
dF/ziGNCdhocrAqOMgR7QkyN3YelXzqUyfU+4onyZIreB2bUQOgrvfeIMtMNA1sV
bzpETiF4Sle2r2uyCy1pfbWtQVBGqtOheXEn52CpJ+66xSlKs4CJVzL3zLdNwuZ9
5XjNTsO6ill2R5vOfe/M8Zbb4K6q4OmqUVSRqgt45oClMjXwrOxHJjYzByFrYmp1
PJcTUX5iOdmbj5AGT6KWbS+RBgmL8cQfqATSIbaphTz9ZDNovdQ/JNmNso3bVrMd
1jlqkMD8rEwbUBmRw0Po6oj6LMjpEq1QuJE90Qp05njXPWVZ9rhMfZMyBze59MH+
PyJfQHHreCRu3lgthWSCUAAAyRX6jz1/DTi/I08z5MQX+ERWFFg9bn8AZRVnKn3e
msk6nERsBAbdj/EYZsV72IQxKxcAiV5f94UZkZ+Pvpan2gzsmJ/f7Uyi6fBGVHOU
f7bf5hhfoeOzwRS7g8IvlD9G7lw5cieg2fWAaMIT5y4opt3xK7suy6NJ28kV2HJP
Vqs3wy2Uiv2pzIuvjHVf/f+EOOX4USD+TQcHL2WprDhnfYQoTkeVIx5G3AMQiRg3
WXzofX190ozdRItFbLdTtmkMi3qWaS8hccfgHTEaNoO7jROjHOuDnvH56UYaiJdS
lMHbqzWEmGssM6qz+pRRPkm2n1UylsA8pHfXD2vCj68kMzjbjxwN+Ulkl8z0lgAp
iuN+bQD2ljfHeN5RFyAVou4D/a2eFcPy39l7tf5P510xbMO0wjRke5TabvRA5wb+
Rw3/9H1s+xaV/tb0uVYEZltea9hM5o7etGZg9dk6XjTNreJFjWeXFiTf+NjyZabl
dJVEaL04uMvcFxLSsKt4BIARTRgWKrtTJmXaYDx3E+CFqoORXmTTlFp/NmeYnZKj
paXm0j3AeqcjjzO9/fewRln4IflfH1w49Rg5YA+M8xAPtJJ5h6HD1i4Voomc0cdz
3IDz5VHcc6rMfS5s5s9DBJnQ0RZJw6GiOf4aelJA3DT/yo7V51aLyka/U42fdIzw
y8rK/xGB1Sr5CJGV2moIjgznrBSluIBVYcX6Xb2mOOs2UtuwzFwsryrI+RH0RVLR
opL0V8N/dsa2KUKIKxctuQ6sERHvMORBuWH9jlcipFc7LgesQAStdsJ9pXHuQOeD
asq7fLLgtQTXfacyKnHADozHkibQRosuLMzv3CsBrUE8YDdh2v9HyYIQs+cd74l5
1uAe/K1quxJBaGLQUYQZ3OPZnRGLEa2xxNHaS1nqKiIii3+OqdpjpVE0nOFyXw5A
16v6+LOBfEXuRqqO/0gnF6sx73VxJOOSbwWG9tFhuKfK3XbBxLb9nFu+I6vM6iNg
31LKD1FXS+LSgm3BTV+qePXcpHKYNOkq4yx31WoXnjnZV1qjXD8iG/JFp8E5w2T/
BlfrdFcV2y7VPG9Jl123/poDFVSqv95fws5H2q8+p2J7Ru8pXfP6mJlFpcKYgxvl
ZAyXgP2g7Fkm2+LrEsu/pxYOCfPCVaOGFhf4tMgGvo0hDaXmW8+QXau8rCxCLPc9
K81e5wj17+8ufi68UaDwZqU4HYayr/dbnaStI1Kx+N/fdJw7vLPDcFDpLcJwKQ5b
mZKvZda8SEw+ujCMEnYLqLI2FqDigKFaiMXBCoPq4oGQrKdFgQIqHZ4fQNZSuovA
S1CSkJ3B8oPdd5PpmEcQohsNb7FsXIpBRV3jtnBBCYwhmGEduvrs47dcyRzjkiPw
tRj7S4BEjlVOD92eEWniBvRiZWTzw4iiGbYWgbkU8jrXQg5mwFDrf5AbgLOaphy2
YKIDPCMRl59uZNjWMPK5G5C8MM709+GevYl6skGzZoEx3BDuGLsQS+GHUhPemGBv
C7/YVZ1yi+ouiURM5c3eidHqve9EMMgkagh26SW9uBlLIrqYH6NV1CwMgwYoweqc
Knxt/eqNxvNxByKH7K0cXMFZ+7qr0/QLq+QTbEFMcFYodMto1plpJZ7cr7UcMx+d
jbu4xHkHOCCrfZWmF3RAk1G7RgzUJRWIv7wXlKegq9941hYkyYXygIL13WjnJd5Q
8BskV4lQAuKeZaJVrk5R+KPidrKe+ZqmEbmd8n6p863G3QRw6gskp4RMrjypeP1/
qD5GPzrdqwmUqgR0y1oss+wYqlyyFhKqMA6XkGAcPZOAhhSaqeqGbbBL9QXxIp9Q
Mxjviv2CaUOqjK9155jiCXVkFuh2O6NbvAo0rVDs9Damr4xxhUHJ8c8CldSgLSt4
Q+obfZh/02hrcFm5FxxJ7SHO5pTyTOXA8CDBCkCMvTqgkLlGu+nX3sY6G26q5oIx
eZLaO1UjfiEM/nIuK8eU06qY5y8Fq2LMb+6H9FmNjBlC/gQU0bdCWP4m5s5KxVNv
caQx2EzVbZAhQm4lFnqHbtUgnESyp5GSLSQML0y+S8aAEi+smD4/q+f8C6p2odxu
u7WuRPqSZpMsfWLEDrIJm/mOGgX/RzatO++G8CRNRZ0RrFEwkG+F3ciDqBIjWi6O
kdXAulZKMUSaNU5L9zeRR059cYCY0sF1glG9uj+ul2kPiaYe30Pz8ZnAYVeTwQ0Q
nUFQXazqN+v8SggGUiJ4QjwgQ/cdHfJW2s5+gPZwJRmOJTCWo8wtzdf4GsGTpSRw
qNeC0YOSQGFdImzU4YvYgL4l9cCi5xM9jL6S2WHUHp5liZJt0NJNedfG6asm6LlV
WFvMkxtygIwEBVRKQm2A35SSbtWVyIFSiCxqFZIEZpSZUanW61l68b2Wag+HSwj6
W06xkyAUW6XHKJBar0F/OsS+CS3SM64M21S0oR58/z0yyD3ihGXMtynL/4/vxeqR
bBfQBQBO1EcBef/CtwyacLsMIL+TTV8eJuMI0qECukZzSx21MKM6O0pP+UwA8Xap
KtkAnJpNHSCQ3W1qsS+zzMGcM/2rl5Sng+ERFMXC7z7Qh6iByIRTmj8FOIBf1+Pu
cX/H1HvI0aPoZP+GkMRpWROJgeFqZiRDWWwSgDcjs/jmSUyvWpol8ez/iL+WcCwB
5R904hppzRDUaOjDW9eWAfoQaUFDxfY2mF5C0PjA1VyAqzN9Bq5jiJwOA5qRNFbl
VgG8EEGsL8UCGBC6U22jvBzJ1L4yarI04PeSrtgkbNHbvP1Wa7YNTvF/tXxO4feS
aNkoV5oSijv5Ao3oHvo1YfZFObjiVTxOXFFpHatbaqSGt5rs/igc7Tu17UgTR2+M
qqic/TvDVe2XuY60sYUfPF3IK5iiteCFkW7FbpgoMVlTik+ZKYZoLmOVN3kKtWgU
70mGsx2pg5G4zp9vAFoz7nE/czaBVCY1hC66nBwcmhSo22HtukmSuvAP1Oj0hlLr
EGyqP28u5gJCfTs5AsV2wULxMZCGHJ+3rU/bRQ/il3HIL/i8KlDficoMhVyDeVqc
PVGViJwJLGSU212r22s+qVky75QaWwAdIEmAV1Fn4rtl1h3jgKXkCX2sgcOfaIwX
L0sZ1X9J8AiMtJCkpq/wNaXaAt2B0kxVxeLLKfDxd2eKwep4ELOBrWMYxPrm95Ma
xgnB8KzzS3IRtdiStv7rs1FQJjzXsocBmh1tKvWSLTfZ27bauTIrt1iF5KlFNVRR
VHgQYz3vc3sOCColkPglg0C5iWyi020of7lPWyXS6LU5XBxTaKBEd2NygwbBpCzN
lg8bfN3TJYkEvbz/mS9A6S5DIhssBy3BqQvsRiK8/29sGm/QtKxODVUJAGH0jZSy
rbRlN3r1zl6HRqalzxmO5F/Z3SVHdGZi517Wqw+DFHf2TJbink7ch+ntmeeTFEJj
ZQ8yEzXnhB4L4LXV7D0PoEi7DEQA5O12Vob/72DtgosMTK3O3z5a6COiZvo5kA24
o+jbGRUSUYgBEII8vOd2sfhtbvLsTdCyHAQVpXUN+GANN5TMtgMwrYlB7WXF5s/T
QFerTCDCHK5xWJlQ2Ir8Od4SvHQ5n5KJThVFnqXPwW1dNBZSkM/leV1TzzwwVvW0
ufwoXZrSQoFC6GsHk4/0LAWDE7Xpo59YsznmCMb33tzKSCAaRuK/yz1DiJXVVIYi
aaYrdgkaKORl96kTzNKCbbfAG1NYIj4nAaFx4oMRvG91aewINzXx128oSK+NZuhf
bHrWhcowhz8QfBoZpkfoQnrVzUqcmgHpFBjIQpqwKw2zA8zQmlfztQpbJRszA8ha
ZcZA6RUb1+uMKcmZLimL7ELlYiF/JWXOed7Ij1Y0X8UAvFPrnbm1Ye8bkwK5CRxG
7uPx3gkfOw5VRZ3sSta89hWfm/kTeRGh0c80cAfcHtQsNcRqgs9EQci9I+DYy3wl
XuhHzgK4b1Uq8OlX+tQgAZ8iLrdlgHutxyxjJ61H4gffXUglVO0Z7sU13LOcBKy7
9YtsAcXJUY/nTrFhImlgJYXRFPBBAX290WiVpj0gST5xM32UEyfUn+m4LzB6o7b5
HUlzoCEdLAPAJAMKRSzUz42xmNLNEPgrcbdmwrXpme19k0r+wcn8o+ajlRy3VR24
y4Fj7zPCP3cBAny7DUiydTdgtJOmcqkndRv6TN5oG7C8SQ4tAsJLc/U8XMZ1Qt4+
gqUdG6GO5Cp4QtE+IFby5bc1GTIh0aZP/IDEqmM/f3keBCgJl792L5iK+ytParKJ
j8H21LfwtC8PfktLZZiquH1qbnz5RCBptlT5mQ73btqhnVfQE85cHiIS9m6Vbiuv
/j9e2oWO7D41DyC1g++sd9jWy83F5vmZAKMVfseWFT0Xn7Mdi1OEzgSYaj+5Gvsa
2UCt8TC3FGXuzR4/x3Rh8X4huHomqOAd5PJhYWO/MP6zm2mfDxILqC5vlKJyZT0d
35a7pVSDMlVzLJuOC796pBWkGLfzLxo7A5n7dc2RU9WBNZWDGIdObgfphmZ+Tvkb
/Ps7jcRHuYxiWi2GMREoGD7LUnirOSjgbh2v+XWv0PxsYsslgx/bI9/w+qxhphLH
oAw+09bRIIB4lbs0KjGkQVwR7rgGtwVy2MZnzejyaZBEbrGCAxakJ/kNVLEPo8z6
gNgJMVL3vL2no6/a5Gj3lnJabokERr/1645iUbnOguK6RB37B7tJYOlpAWRp90O/
oR9vsn4+p/UV4M19BBK6F92qdeiIVj3MURV3H+DSLFg1IlM3un0m2gNkUz03AKqs
G+kMAS9vxxfzHiUtaLGjl9ucmb1g3hwyMucZMKlxvuZ5e7W48E60/pygkfyxZE2M
spdUhJrCTcoFhH848mdPf43UILRUPiD8ZTXkUezYOhqIk0xhH8ra6DPtFNvY4yJO
yXYyasuf4PeA9Ko89fz7gl0Hq1yoiUXl5tVVF+iwMG3Ob5NXjpNp0bMxLl/6jS/P
OwHxqGWZkX+10NK9epXhqimD5Lw7phYRyBIxOAuuwDTjxHyJl6/GmAfLGdgKRmeH
vMUDwuHnKBLH921LCRDT7o3cAWRxdSSJhQ/IgmoDkafRPjqDC0LG4D3GAYl+iwpN
mm5mj/mI91K4m1P0tKgWWe4ldvPwjCmGc2vIarERy/wiqUCcLA3znp+hqmuhkYsW
RE1Rn6qPy/qZTlphryhB+O7Fak/pTL5dIJlRXUC63ZAwXYIksZFcPlh6581SRMlN
qw8LZYquNFFDd1AuxY/iUmyS3JsHihfw7Pfv11U7fw98to64QyCA3jGS+YH6aC3S
8mQvJndsmYK4V0SHug4j4Jf3ii+fzeti0En7fEBmwVnasidWA35/ggOjEIL9pMW8
C8mnBcLgklsTHN2FXEJP4cu7LaYdpZYvqfEL3NaIehL+ojfhkgcYmt3wypE2H84l
LWZZuyYknu5kgMFurnAs/FoKvMvNuw8aWhyPUMIlZ8zLvOpu9May0ktgFopBBl5o
6O5FADwzmHn2LkwwAtyXRi09rtCtfwEaqpHjiu7qBLIDJAlqj5N2O6SO3NYoXvIe
O1bo/ZGefJ/dd94xudaIAKvoAN1VL2ZcQQ+bYm+mlSNqLoumwlfuRYOaJi4a43sq
NaqNC6RRpCN+UxHnq3W885KjPyHdx5HAY0dDycawxBSbAyBmo84DyubFqDXnJWcW
GQ5EdnuDJKt3cr4AKHDDhBgWm4ge8Ry/VoLXC9CDSG1EZoXh6nX1qCih8tgv1u/D
tq6d8OMJD7X289ElRqZb5BciJy0vwQGCzx4xJTw3spPkgyqpG/rs0AobuX2qyXWd
y+du/DcYNiDK8ZIZd4FWWzPj1ccsjpEvzSKpyMJkAj47oht5tWNO7rMhDNCIg8t3
TaE1QZDEpAB+Qk4H8rw0ohwCT+ZLCTnzyx3jKNVUU/5i0vRhPSpXVcJU6CGSpRwQ
9YGtiECHRfjLGX3ntiKPZYIFhwDzLvSnfHlq4ovKdEFUfekRX1b27uDH4L7rkGa0
ONukfS8AbI0OrBAK9Dgo9Of21Wb5bfYqWfxbjd9B5nymQm5XaXYEU2TlWwrNtQL2
xWzOA/f+HhJEzR4bgBbwiJMI95NOTP9i6OSS1pRmPG7T5XJCOrK1PGaW6uBL67jP
xJXK3eroPMddVHXcg5uANOmO2+qZWB2nY88f6nGlIgGkx1wOdgfaGgu+xZXhVNdD
xp9dcKGYlsnpAF5i8wwgegXD8KkmVVNFE2ss68I+1dAs9ABBOGH0DFaOh758xzXd
Cp+eSVBQldchxW6rFKockInQJ9g6Dm64MjZHrpicQ4NIvfGuOrNYjqBorFI1buZP
e6AUdmwianY9lpPIjVEelwjdmN3cvK1a/2UHHRfhC0T41nftMPiR3F7oZ3iLKNNC
BJSD5e6++gJZZps0RIGWgd17zeZF7rzy6JK8TCXGmxrW/dKSTh4fxyGskldb5833
pBDKIRM3WAoa3RDUhKJL1NSYlvRT0fhsuaxYiaV34QlEQigOs/JbsBbk+ZzTOR7t
SJcc4pTrHlq9HOVQiZy8b1dKvrFKUbA//nOV5LSwkIZx+az9qwNiXZXNrqtnkgbL
5Dl+ZOvDnzzwyxSqua1gRTYqIk0/2myDMlVBLGdsTWTYF2cYMPRcsxnBzznGTwPM
/oRzxiw6mt16aA9TfhWKBciJCvZaavxSEPyBkToh3QJSw74cBQJVB94VYT4Sr3Mr
pcYCYRDU6CJQnY3R8nGB/PVJwl4AuuXKDGu16QNLgs/5V7NykuytdrpUR8IQRubc
xlD/WsZiTRkRMn+gefWg5Rc1bEYXbuSw0Xcm8SMHMklR6xzjnoPlE9HGF35q25Ew
kLYNag7BRig7JrLxYzz85cmFKs993A/juKUX4c7ZMFV5LavSCRlfvUpCitMHs2Nh
bkxZ/pleWZZdA+yKLG7uZpYMfDKoDlzJto0uSgFrb8j75nDrjAruotTGSq6n6fr6
Q+a+tvGLbkBxYD9JYrpvs3x+OI08pekCutoS1lCqttpYSGNBTGXJYMkqSpHYTtaB
MT1hvW2UJwFsASIDZ7NhzKdDAKVmGjKjYKOewD495RC/m0lh8U+n0zLyad1/YiI7
jRF9puG8ZEKbIEEvn85BkQTn+TRSCdsgLMdSnt2FZ72CZ7X7o00bUkS1+SFkJHXU
wp4gvBtZXjoqOcakaSSJX+Z8pZDuN1Mrq1o5gpln5AOjtm1ljefqjg7pC0rifXEQ
BSo1KlqnhneBni3oSEK2zbRtKCi6k23p7w4dr1bVY1/xpjLT1+sjxIw3vFfclfGZ
kS2mxa1J1t/l8Nr+Lnj3i+83svyxYf4MavLRt9w1y/RFRM2MpDq5cpzW7wCCrp2I
ditgSTaalW3EtSdOZgo6PG02Yfg6GhVk5wE+egQkO1u3t9aHR9LrkD90icIhqG1C
+J59z+qn7dPJNq5E9a3BQP2kXANHxUZ6N2/GQVqPJH1UkAZqvO2plsH0nu2pZhhh
eYjgoHKuIEc6qYVlve++8sQzIRzDbckoCFq8d/wowRky05AoQPNtNt8UalJclPdd
YOxaQPe5fBlm3TpNSdo6fNbhZ0z4cRWiMGk7ARS53OwqiXOfkmZUznRpOL57T5Z6
d9OBFUl8IpXTxv3GZDlDflbQAcoJCgGJleBQ+39w0W3aFsctw3sycVp9DPnYlnZ4
zY50adZGlrcjNnw81GHHYWhEWNEjo3UYuqGLXPZ6Bgi7mSBGO7++jKh9TxgflHUG
6lSqCcjOX10I7w1DbK/7YD8bm95V/DExfMITzDvJu8/W0kzfoIVuUaOqDERpj2RB
2Ift2kErN5zR280abh8uDvNfrWFdxIjIuQrxy3armWcUU0lYjR+YYmyKTf3ioVJH
+G2mElsJkqERf0qNol5zFafOhws9VwjlMQaYNtUBepTGHDeUM4dpgcCfX52JaSQc
2pEj8JoJbUAOf9+PQWmkNmHX943/jdoFV+FNQgo/H82ZFU/AiPlhlXUr3zHmF0sN
AC32C5KscKMABxqM8vdNuT/yMqX+Si7Ay6r2lIhMh1ms4bxsXAN+q3TfIQ8v43ra
odIxHKEWbzbt4+zfLa23OgGM7Hj9IGiZcS6HocSbdWsShHJoDOMReLjvZzEvHl/B
hA6i2JSicDZt9y1UtaxL4itDSf2AuAiPzUo7eKyij52bhIYhO5VSrIxi3eJFLhfn
4rnone157PrkAKeN8kEAFvOonKdYOu3iK9SWyLeNQSRuafTQveU9irwxQmTAeVH8
sEb8FhqvMjSwXlFZBtlgu0tb7FAS3jGxXQqhw+UUazEmO8WsDHr6FnkxEq+dRJB7
oNtmDb3Ue/0+/1CpKrpJh7+EAm70OKJKZEy8v0Yw6cRuaWyjrJXquKFr956Ws2zB
oenb0TqBWzXYkHsglSCkHDuDl4ZUArvqEqdhu5IjEwc7u9owV7DuhATNzakm8Cjw
k9DyrzYprylD+OTdbZtGb3KK7K8zBcNnARjG9XT59ECbKhPbJKnzctUqx73rsr7+
LmzthODmSdeEodcvNbDG70MORcTABnspsDDaSyhh5opvKCCPSZlC2C02VpLe47A8
k4eniiGdj8GYuJexeIvYaH9DvcaGx06+odu1VMz7xvpvcw7TNpif1uCpqbDetUFi
DXMUqUmlE8+esn/hAwKbQorpQMbpoch3GcEiBhXGp14s58s1DhjnQEivrTzs0hff
HPgQVAELS7FS/iu9yCR0ZJemQwcbzEOKB62H0EeX4K4n8HsMpnyenLAh4PLZS8de
W4uvS7Db/4xWj/NK4UyOotz7ZvXvzgOp6vSMP+zphldVQyC5O+rd/5KdMgNB6F5h
cC7NmVBETEoPBZIjlFq7KmqUcrAndsUD7a0SFoTwoTyBNMVW2wPzr2somuhl14uE
PUtDY+qw/1sZd+TioSsdlFL9HZRZtygDvHYwHU21mq3YDRE6cf5sf4Jmb8S9FwR8
2KNKG+Q+9TWI6Gwc5UvJh7XDJ44ejfw4bVJ5NAmnX0z/AMZ71OanH8ZC1NjWOD28
GBQpDYvNoO6a0V/6gwP3SYJxuXxMLJ4Bw9lMmeFM9IBga2wGH2BQ3zDPXLmZ96RX
mey0i1NOl2rS8p3BruxgES+ad8CaKushE7HJx5JGDRYfV4dQl8VFC1xQg468CB1V
rgL3oj7uc0XkHi8vnTSuXrwSa8uGFj9Y+Juaf4cUgDV/Nak64qnuMRuWDw7/tNw3
LoTBA73l5OAzTFkQaARMHNddx3GWfcTlz6JTgV0IJM7eEJekUqcaK3LAK+/9aXDN
u6wcG0QRjBPdKQeXSDNAiO29Pj7NZ7/h0NFxfRu6LHMtN3x/isewI5iS/86DadfA
Hzc2V65afm/Q7Bn6dUXH3jSgdxH70fqOM0yg1l7DyjYp5Funyrg4MskJ6GXxNmYh
fsHwZ6cXpPZgcwRby+1O4qyd0D1XYdB6N/2Ofl0flcHKdCTgXubZ5TFohD7aEwu8
G2BVbd0UnHPwP8h+0q5mQRYLPcY8FDgpP+QGOxgr0QjNsX+SpMTYX+leaXkdFuta
JivbXZIG8Hllt9yEZBCmBHMuPpRN47Sy1FDKPSR/WkbNpShdwX34mUJ3YOTqU0J2
6BCMaw0Z4at+z853tOfX3rep6BJ0d1lbwPw/wlMPENuQG60MaH8Ty/CzW2berbol
MPUpkHQFtxnO5V/r44YyBvcZwdquSDHjf5KCNiADa1Jd5W/TUYvNBtcWj2f6+zXl
ZrxXbuv/bOGLZ086eA005+c/+LA7MgB4H49y0Nv9VEtculnGW3wAAOLnkkfSrxW7
0l/yf1PFg1jfBnL+fw1RBLJxF0bis3KETrXjgti2jOgJZlw/4JNT5ylkniZkxhDz
IOhB7qVJ8vQHelnmgkeXLFDamgRhmnOzTVk/7bxbgMm9zcsUDoY3W1I72OouOe70
EUUVBNfwGuOqcfRSckul6RKC/dSm9+CiybOLx7mhfxXBeQOiFdwmnWzLqkLBeliZ
zQPuZUZY6+gXgFlamAQnWIsWrXe8aZT6hrJw9jScxkabP0Ktk29Zc9Du9LpsAp+L
f/Bg2QP6a8FikwpJUrCBGSupPwMsKYBjkFAUulhYiuB9lw0+jH6PwN/z2mUsYLU4
FN+7R8siJou97GGazbOmmQKY/80+vryy+4ZEfCUkDiQ8VP1uP4TU9w5U7yIWOF+b
VFFI+CI0FzYxv2Lv3oYuOYTFY/772HetfZcUcjhjmeagOUv64QPHOASEWXAPgBmN
jtXzpi/raNXPuqChucqQHuZxwJ44EJqRwQkGkXv/0d+yu7pQaFcXU/PMg6YZ3NUb
KSVXbCPLjOAnz9EApuewW/BKUimj2veEOw1LCnc9vQYEIGGzrzOa3iyzGhP9fSjw
JAzsB9Bd3mrqvP9eu0FKdO9YVXdcRXwndfTwVFrIgJFfTJd6//N8SxSjQ4uSh37N
aW9tWvOo42aWPrdL73h0D1hNgaWL8ey+GIksooh+14bAc93SwW7t958OBegImu+d
vK6HzPNrz4ZQTsZ9n3rpfJG983pvhdma1Y9FZ0YyhB4kssZpEFJcfZSMS0FbnfCS
9cvIhy4NAg6gQNjUbPDJZrF4kQiLLY0hkCJxP03eK611h5Gp882rVmOIpoym5eRq
U5OG3m9xBW6YF9vsBUB8Y6IbCsXtD71rKxjQ5hrpER/x+Pu+NSxtxy+PGOKJUxiG
GgOiN0QkbgslCcseu297v4BCUKNalwuhmivG45z1WlFO1im+cTRRNXoY1hT4g4aW
qKOFIkVL398enXrfJtuP+U2UVBPQoglGLv79q7WTkEk1/rcO0WcJwbj0xk+OjDUA
iVL+Df7o//fD2Z5qcz7wlutJnXZkZ7VJGamZw/T2mIVi6XjdJLKeij71cmq0bo9h
SQtw9SuJR6xqbqxArKoMRkoay1xuS4VyJ72XYfI1a0oJKwK+Bk95HcWOWyhoHTm8
gvi7JCugUTjHQRBIt+poRQ1fJ9OYjCULwmFHJ+FGDD2yemz5SsNznK9EkR2hXbVx
/PqikWQhtKJd5Z4prsloK+7rNBDzEmqSqpO/vKyH94EaX0+W3wj+i9Iu5fp4um/y
drF1mZQy4CS7TC5okQrR00DN1SbmWzPptc7N0XxejxGNZQS5quRb5LZdlk5YGHUH
spg2vXojACmPoaBWQgZZxJO9KbtcUDcqUO+t8oTfvK021GtD/m1RS36dRNqzMSmS
nZokXXOhqm0FxpQGOlaO+9uSvUPC/BhNc+suTDySe77LqVsA/KY06qAjXwKDemzs
XhhgJ8VQl4QGSnZyHDk5Sj/Z/9jjb+l2893LCPC5k7XWyeAevOYIt/OL8Pl6FGNd
tbm2Szv1iARus/UdA18jQETMhPqACA2rrf2zBg30t2svRAVqNveZB4ZrsLREhzPz
G6X/E0qXjm3AggB5FIjDQX+zAh8BaiOIDAXRUqR7Lx317NzEXeAdSZNjLC1wkadd
8Gbywa3u7qqGE4TVoyAYuWcRlRZku0duYyEog74X0acMpESHXzde/Z/6cdaGSHV0
baGYwnwICm8J3pWISomMNVdZ6rc5zNDMj+nqi1CAkhv4j//9snaeEPpMlZ7iu3FW
GQKQxNRLi3jzbrLUOibv10KQWb51Gq5WyxXqhCsoriTbEc84r8HCM0IoW1lqvuuZ
hiuqp3AwiSLLMiMQ2Mdm831nZaGjv0gAcNyEstLuV3P20VvYva6YTU5wyML6JGiO
+1C5ZiDSxpNhAThoowCPqY3gdDSZwUYu5FyI8zZfbiiTlBwP1qqpECxPrna+4JZF
GwUDl9nJkGvl1wnvyFxtfDPZMdbKbsY4vE1/n7P67X1QfCsr+p12qwNxxe5Ex4BH
RgpAYtytMiGBH8s41orsnxKFDBVW0utCAesZ5zorrDbGMYtB+m3EK6an+LVpAcA/
XnSrD5Y/1Ti+27B34xGyihMYIO7v+kbXD741uswXi5bs+vBl8D0oXJqoDTbZtEP4
P8EGyE5JM8gARVJsvVfcgDJxJlSrclJSaZRzQWEna/XHdrkkN2c4m8VFUW5/gwIg
wlekDClx8VHUwLGyYMn/KHBxhiqjHDhWrq+dSAfrWTGAvAEDsoD6UZ/Di5FduI/B
mHLDNHIa3nnccUPWO3jnI+xut7ce6XdLiCsVOxVPQKx2R1emOLWkGlzk7UeNvmMy
EkB6IM1YsJJxPsDdDd/twBW2T0V3h8aO0XyCiNnbxLGT9g8qow3Ar15Dwlx0EqM5
UasQx+K8d8mIrQmuFf71OOlWZaLgQL/uT70Zt3oLjG5+x62GEQrW01xF+Iwmz+6k
14DmTLMYOeMeqwDi+ObqdWJrqDnSULRo8S9HzfiJRxHonrG46dQfFqYtnq9mbQbL
aDn43DfJZWlWo5y4QlXymOYJZUuVFTEYcrAklee2dBK+Rq/K287coXy6dZ5vpH2Z
xY0mSMZKTaevf/80EvM6zBR6+NzQhDUWG5wYhFZhSMlbqpasbXxcTuy0yqM2SOk0
tGD2eTe2yE3ZAngAsrUTWHqtBu9ZQyJe+FtswA1rcPymHtqeCykg6onGVxuM3QSy
qVQvMLkVrzdW9AQpaUZ1WyQQ2okjPrAd9tIYcSUwu6hgnSFglfN/PyglCCTtKeg+
PNewezqxKTVTNW+6M5aKpgZLwRPAlsYyzgctQEAirSpQUUHafc3Q+pZbsxDdXCre
06774xf4WPNjWCsn9jBYoAHVC52hzSJO9W3LhCIsHKi9iMDgPfpFyTWPlgtdZiwE
qCEo3bAbuRTdC1aE+7Xy+rhXARVJhvqPvVKO7rxqdMjFVUseMOdUv3nArmM3qbfi
YVVhIAbCxCeebYJSDOvicCb7XsiY53KuBg3OcI7YyRiMC7Nuh4NSWHnUJj5/S2k/
HItXv6iIPCDUjmyoFYVnsREyYJ/NrzrSc0CJk0ReFcj0OhUktI07fqrlsFzhogZL
PaTAdPjwS4RnPK0PgnCAvYRTXMcrtepClAdEyoGTYtM9O4vNKCQaeCCWI76Dt9hM
+e9nfTv5Ec5/7PlDf+pYCkU+p2vqG1rlFABeXpASkwHIpEC0kSSDWxvBRHPtNsG4
psxftpvJFBCMn6VfOYHADuRjKF7HYg4+egk8ZrtW70gcguuJLnryY5LT+g0XgdEU
BgE0QBaTzIK1DOjhERenwPOY5GX6JHtgYwhmS6p0J2/dhxZ2zNmcFdp9reK9jZAM
e8L9DXhLjhFrfED+i5ZYnZRwXWVohwPG76ySxM+kjYBFOeBQWzkl8ID9X2JscfYs
fUKQQykMhiBDYVahfc8HNhrWCcHgSw+SyYmsgj58T7h6Wjr46lDhSzWCZFi3mWR0
W+g0g/J7VOyYOHSXUQSZ0ZJH4C+HHalgcaMlG+HJhl8IBSUMvDGZIVxAffU+sEYJ
6iTBfCmoLm9raHgAU8/CHdZmBCBLa9pBlah318ncuK9B85AYt7b74oChkje3oRbE
arQMIyleFF8s88pqrIK1vKd2heWXu+phYxZBv/wQKpUHMJLQxSWIFezX7hHt7oa0
MeCx2bGMz0zvP/ekc8gJg98s6qNX9T+7zWEAN1lox4Uk3QhFJoZzOMoV5TLgj+Vi
l7rK/GnMyWUkQIuIWgzYu0/jldSMfAXkVZ78rwi4hu5b4/At287vYym7a275KGis
cSAwMZ5AhAy8f0n2UDBGH6dcD2X6e3nQbo+MO3Rp8YNfafNHf+GKD/8nRS3eVJii
lQiJl1AX9G5ft8oZ2Y1Wr6p+AUvQPDllvHp5fdtuCNQM0/Pmnc0c6T0KP7XngXuI
hkS/uysxDCFGHnaTbU0Yb+bUiRN0lpvEf+xf/DZH4W4iiIL9ABgS40P1I0olMO1v
XS2edxIAZTcL+9wtSb7ECi8JwFi28F3I6Wu2SUd0OD8AJny7IKS7OVpDIfg01iT7
r6z1HqRPMOkUPZTS+Smgco2DMKAVfdHaquu1pcos2wlkIno5Kz2SBBN05uyrAIeM
I3ESoGTB0Au/CDFvjDgXfChluZEVy98zUKQZzdci9DdZmBlFzwJBtXUUneolD1OL
GM7Osntyn+GraWyCwnu5bEcq32In+gCWwsceiohL93r9H9hznnEnzSP125D7TO8d
OmADov2FxPfRAVBYi9/EoH0c4uAWDjFpKYfZC5kk9XslvoP24wHA/+XVoTdo2zXg
258dzHyQjHaFfvqvQ7X/CgpyY76GoU3O+mr6gJAFbnHCfABjhTr6p+EQbQV2qIet
aEVBMASCcrlB9xe00gRdybyrCU9OvT991AXtyvOKCwA0mjWRl0K1JKe30xug3zTA
I4Z7FjYmEG0I0EnWFFd2w0xJ/FYCbA0kJQjYKh4bHMnBkQGkiytLRmBJoJpAOLIn
RFFdcu3WQ+d+TQJ2WgYLUw4KEoIoAp9u3GmwS9X5X4eg+3yYE4XRVt1VYgtti+1g
/+gbZWB5m8jiqQd0mi5XMo2NnOQ4b+xg1VRbAS6QqGcmwoeccjF9TrdfBLidzzNo
1iRsLUzSNvvI/KtDpgGOtLiltIE41XVItTjg+s9xL2TcW1xp+DK+y6JjzT9SA+qG
n2itgRAOTXi3m6iICSFsKl17hUr/j4kPyv/zgh4W0G5RXQtW8e0eh9/DertGWPeb
Zncv85L6s95oGhmWehhbfonrU3xUsLvURNCUtw5EeO5zFi+3I4x0Wpu+Ljv/V2Fa
BmGvEdLWrPxlilFf4vtJPIEWNLNiBlJ1RE847vq+WISLLrCsRIlRkB/lJa0ZQRrJ
icIjQxevoYNK9ZWRZXorWuzASPFEeDj6J31l+p3EVYzSo5v9QaTbZtl8/DzLBx7J
tgh3QyrE0HS7YrYALMe5AdxmrwMkHysPtAhVjAOWtYGpEP3O890kj4Wntp4nPnxd
65/b5NFVneNErZwjZoIs+AmKcNTabYavdLBVGL5gb1ZUn7s8h7OnreeS/RHGrnuX
XgREaqpcmNg1Wn+qXS624DVvR3Ln6cnnLfTweKVCDTRME4o7YdD4mgDVtAQpaN10
blCJEEJSjAV9apDEZxcj1fc21zvy0XllqM0EU5cr2xc8mmaJRXvV1lwQPm3AFJwY
zlXoGvS0y1wNrm4BhOQ0o96CLI3q0tGQq86eJjZ/TSZA2UmPsxd6UBRqqBIWiy9+
qOG18kq2+bd4P7HKhCpX5mV6IJHU8aZNzwa004o071+Ml7ej5GAEX/4a7QtWaN7G
QdJZUvr0YLhLFAw7rGLVUK4syG2vs/gsqsNBA4xcmUaW9D2QmbK5rWG9sl+oDvr2
LZnP57VP5w78H5zOu1IGkktSqt+/XGWMZrLxqHxF5WPqxlXvBvlCGaWctvhI2uzj
IbTHOkl1VsjvSPlf+nBLppMSKuEXfhMwN5G9W9Cz1iiXNn7Myfesr6Q27nUCVqtD
HRdPyRT61aasLzEpxxoEuTmNOW9k15s9U81srtyvnud4UfvNuePuMZysEcU7CziO
9CrhkBz1Vp7usNyHg5fHHBY3FM4SfnxGDvaMjfve+5VaC/uu16fGv9/Ja68zy2bP
eaZ/4zHFNApJkby/HclglKgbfAN+Cjy/CvmbeDOIdOXhAwRqdVORRWEKa4enGcLw
yVU9RmI7eVjJ7z5s0JKTPpggiHJIC2azOiYPjnhLedJD+/2ormGWYuEgr0rGk1p4
bO67cF/FNvhEm/mj2E+4+UpTGfoMs0UBppWRNBF03rDPwD1z5czMqlGK8EGjAiQS
98hlxKujlS+rx4gqfZJdCFXGRLQWjlnASybOaJip9PtTw5CQ2FuxcVniuFCAPqu5
FE1XxGxYXvMr4BL7o81wZIIPtKEF8ZjvZG/G8IdtjZjVbGdBj8Rvo2KbkggJGeBS
MPw7qz/igaN+dDhyxv/K4ZoAVRljsduZjIY5c+Y/31AuFK/pQwYh7N6ogkal0HMi
2mN61TXj2rHfILPyR3AyghB/oxsIN6E64aZH2oQ3iX4eKPm8pUgRPOi7cjAYFw3F
A1qu3FXIVJQb0y0L0p/6MzvYolybLJzJQxJMwiSUfbcsFa8KPUoRWoN4NTKZNn4D
l9TAnG8AP6ljA88YhJM/kq2/1hrNpb5wO1I3jGMj8GMWP8vzmo/JlG7Kv42LSA35
CHT3IbxAfvO91KSzjlaIxidAZgppDL4b1j3dNFnhaGbCejrsLYtWi9SD3r/MzDgJ
M129+bf88apmRER72JJwCqCQVzeIsnMNgFoETt4gmKj8pqVr5o8LrzyjVmyh6q6l
Y3gXzvt5aknEJjvuTWQPGp8mn8smVYTJhWlcnXkhTyAQ0cRd6PoM9QamGBrsB2p2
xvbT3ei3CYG32oUXq/L6hgJWqxe428rusMjzSjuxXZ8RcDnQKEqODJxI4eAXrZAd
LXyccJICD3OL50hjOiDYa+GysCrSTF1VtadAK3dDjrodkvE4xmwgAn1mwzrBFlaW
iFHM0oZDdXUEbwYEz6clxLoiT4K4Trul049VYLpJU6jM/2TVXT5FT98bDq4fPvcK
XpQQPczxkBG/0Juxo7SlFw4cSdg6PSFeHi82BHgcSX3UsiQe4lvORggRbQmmV3Vy
mcu/yGl8fsTsVE2p/Z5ja9YR20iPwtBk2udMO106TcB3zKvmE++V/PH/qCiykrzA
aunQzmeuPM0aRW9FFYegULskEkXm+C8M0qCJioyK0uMRK2qIf2JcxmwkLFy86kWy
gpzctPqS+HKGP6eQE0LGCpDZXBwUeaDN9ZzY+gu1Z4R2qT3MkGmyb61FQRPTBjLe
oHbQs3HpGtxd1PUqRkqNf/QWenXWfZsgp2Frl1nzdgVDQFc7wJneAW3EMeP25s3D
wtfPC0l44Q9UV+fTmgiONf6wbL34Qd9egmA0oQYMykmT3NPicJRg0W4cUKh0MXwd
XP+sojWfeqCzF24I+jNOCJGJTmu6CvAxcgOkEiEQkqgFPf2nULWxuyWfQZFWPQ8i
Cs3tTzgW/PIAPjmslbHv5ZSiINmhTO2kFsKaQF+C2cP7FrHGW8Go6KGa6X4DURgn
iD3ZWtlI4pdNuYx2yxMa4/pGeeAznH/Y2QSLK/L99yKYwEwyRf4cdtn6cTe4ZdJc
A8KYXB62Yrse5CRZrFIwxNzj8BlOqgQIYtBgJjgoB3zcNhlcCjGjlYM0I+iP5p3d
/bPolchYSEvRgmAdW64qstQV4QRsC6nixbg1tCbDLx75IuWGYqF1ffU9lbMCCJs0
jCaG8dwhsWL1jKDHwxT/ucAAorOYg/zuUNfhPMJdUiSbPlxwWpO7fxZ5yHuDlfy5
7T3ua2oD7Q70ACMvv8qBLg5845LpclDN8idBUT0n7LN8BByVHO2CcNOZE0FvEFzq
s3Wde2/ufWJhtWM7ZYgfe7nG7o2d0hNVDVOhIWxvu/MfLNmgEkNqkZ6NBMJN4shZ
NaI+xFxlHN7+rMoL3GI6We8PrKxtA9XXoR/OXFnAE+7ScJVdRg1ja4hd8zyvNAly
6zTfYPMLKdZ0aOeP3iM+djc7sTWjibYkbOeqcJdItq/5laslSAYcRccsJklGEvE4
d9xEObMkzvzbFVDXNs4DKb99ZPJ23XXxbmach/ZVOMvguqeLO66HrUgGLr05haQ5
duQ/M6PKYFa8z65F1/DlZxhNzbHtDeuE0eLVUBxPd8kQnA8OeUqCbr9WEk2n8fZd
7XVDaXcWvhiakwrX82B/ZWllxrtwsDeIyy9lZa00DLYGLg/OW9gN+jCw0d4ynyTd
nl7skxXI6YQBp+djE6Hg7YTMbeGh7cHk4WabJAHjP+071jZocMo0tv4cM274HjFi
EctNqL4mh3fwZOgrdCokAzrYCVDhmj/Lru4aqxKarttKcRtRe+r8pMOOt/3O7B9a
IXpdWdbI+Z/IrRdfHWoUoxu1W3luEoZiPCRX4DUPj+AqhbDAlC7pCh0zI7bLgGy9
963COgzES3WESzaVZaVeQ/dH7L6cttcDC4I9O6P94az+IGHlzAuQDEul6SJI/wMB
96cuM+iwIKQnexopmgtkoPBAYSX+zJCiMrtxp3xBM/LAXUMv/07CAJ7mYGkC6vma
3w99g8IrfRNU3SRPJmShVOn3BorSmV9abqiy+jpRIF0eqvhzoiyao5sY6HovK77S
KwWAhmEnWT387qHz2x9Y6tzgyIDfqVx4lgXjrY5TOfJgwCPKEGkBLRgcWqUoVOto
ZcTspeolB5Tsi319HI97yS247T9Vg/VwerUDpXNuPJ65iuqAEgK5cBWM/AnHGYDM
buPgS8gXZe9roBByhE6pD+gJ20rugRCecxB5GVqexYboUn/vm9GtN5D7U+5D+avc
/HbHgiYgau1p8OJhals8tP7ACATejoZllZT9uxRnWfx+5cgdPv6+Q/IErlCJhqMm
4XatNhQfeR6WZ4Xpai5qr0ObFPhvFWJOccf3xQnSpHa2pzOBtDPbv3p2ZNwkpHWh
fJgHXA7t9ng91CGVC/8o0YEcObcJHVC0FZ83pTXt2g0RdWUYQib5qc7L4DkfTB/w
BJplYtgL+d6+tQkumfLlXSSg902AfboxQAfTzKKolcDXJ4q2jS1ZXb7HTk/uHSNQ
c1lcW70pnRhwk4mCSD9N6NzS2uaxW1jMbXwB/ya58EXozUSY6MCh9tgcJismlDPO
es6I1g78kGrFWPMgi4SlSFfAAYo5o5qhln9RBZSlkfLl/s6Mzs3/B3KUABxK43GQ
UKF/l2MuyuUl8VHWr8QTmy/CnzhVdXKKt1SzL4Icsl+Tw1I1JLVP1uojDD4Fbhha
4BtTIRLRhBC0L424fVaCbXMQFCiJ1FNX3XQFj8Q/OUpDOuztPd8o94F2JC20jr65
8bdmAkgg0S09ePyH7kJCAPH9qSV9N2NV81eA4Goc6C+kEYOtImm6E7PGkBNUjjT8
D6bkGmWGdKvPHo6C7suUEx2iVw0VKKCMuJ6qPAJo8O0YrVm8HR0ylZLFsjMZAE5o
ldy1pSEuaQpqbb8KCJjWj5SPHJTR51SnWNSH0zHNV6BX2WbZmuOYoOeo/Ydh7+aC
fICQuqSznFQlS/t3x7MATjkVEWItQGstFSXrl9AcP2YJfduqQfrgjCTrqLhl6eu0
qkdpcLBPJyKz80FvJmZaG+Vg7g7EzWPsyffGALGN1Wgt+o2psxM5nVHXAz39Jfh9
ThvpKBBhRjP/m7XS5Gk3HeplULqpncFnDef0eic0iRRq28435NiIRXCP9b9B54oQ
IHf2ONP9HTGysOYkUVuQUXdp3IlRTvpvnOHvmAG6IutKmia8ymQvTbUodEJGkQKr
5IhA8U6FO2WDNSDATo20JsPV5MGV7XAGuc49989GWYo78LKrjwzG7615nGKh5r7v
vIZ2RqovnmJ/1vx8l8jgqKO6XzlGy0LaRkHmhqaaV3X+H+bMc+619ROc0JOdc1J3
8rnv89S6LK9TMfSPbS6qlBwFEq8mRLn39ahKrvU/saWS3rnAYAOumP56OzvRLRrW
cmSG3FGSrwAZemsz/kcTkTsleHZNcKwE43hCOUe+1KyPY498wQRiRREiQMpo8S7I
Jt34N1f1TcxMkcsNQztNLI9F+usSye0PmT9WTmt+UnhlEmyLZNHw4nCDAN44KiXC
enDFm1heO9bbuianXl7qJArjqjFanemUktTW8C4y17DY71r36817bdtIbXzbouRD
/u7EIMm1Cp2pbbDPxTv3hrSyTe2WrpXkBEaDPHYtJW1wyB4PVM4B5ZFLFzkl01T5
9hekdpXiidkJQ3UJnHxFo2/vz7aYwYCHuB7qnk+d1jiuvPAZAOyloP8STTtVeeai
jMkNkIiT7lG8rjD4f7kC890wv/iR/2RxEwEhXto/mMwCFaTnS1vVstmS6IbZucl6
VSykIWTYxlLx9AVI3EXQjLRTIaLuHuHGWzGOsnTgOWu6G6NV7egrVvXiHSFTBJyw
Oo7rOc+1orWj+lxxG+/inpijXhl2PVWEqroZ2cIeHCLd0ikWULstBJ4g+5nAkKB9
o/wAV2TgK4ElDR1wPGwx2eYfMqEck0zuZczwU0pmhn+ijubPjUObzQq7ruV4GDAR
Cm90sQpGD40UCgGRoyHr2wv7ScvLRZlPx9uEOKyNi5L+lLLjEhhMpUq/wi5fPiUV
kC1WsiU1WBAWnlvNyLkuz281F/1EhCf9IvFcSSi89kJSewnrpA3zNsz9TXfT7elV
KrmzDYLYdELaOO1oJxojoYx0zzGxJLPCV2Bc1S8QWML96Tt2UR61yvcrqwjZRdNJ
taSd082nxNkv6Su/ZAD3qX4fTzHdjx2S6A4emjDiqYAmXlqORNvpSYo5SJ405poR
SqQGFsUVZZhzCC1JOSiD0sUG6tIGvrh91z1CiSG3rvzPN+PEfXlFI0+fAsAVu50f
MTNQ/W/1bFnnfkHOw12LuXLBndHbjnUl324288XgW/avfznojL21N30d8Zeqxn0P
iBf6DqA4uS7MJ3r7+HMODBpZdkMj7f3vBV8A7ylGsyao/F+TERBM3TAuUkyv99oL
s3KgV/PZu/agIot5p8uAeARQ4hbPlmF4p8RGqgF5s3Fv34mo9pfXEs/tR/lBSqMC
58afZD0Tu/kPs4XtUh5ZOlonEkJ8JIwVth/I6WAyu/2EME9U7rKj9lOVv0mu3MoG
0Epn/WnbJSbXN6wb3oQTXiezep9Gobo+q3A92w/cZXXihe+hVmKMOqwbqvwuUm2L
js1uXL9NcYsEYrMn4438q5JkL+189PF9uwF2Yh/4LtM1PThYnYs9XeH69gh/Myxl
qAn+XdGqFqs7RmtWLTKkApbSnmcyVz5ySIRocwGDGbPREVrHnWeLIUhoL1ZnrtYy
LIbYLxVPmJSTY+Id3vB0OZ8Ac4qhiezWaKFo7hicXg6Bc86w383N7ug5qcBQutlZ
77p9qxzi6dHqFAeUmEKnU0dkjBKQoOlcaSsEjTnHfBxZHR/W7m2njx4ryYmBbaUV
KjBRaETZspXL74Pc4cafkehp8inf4Nqb5c4RsctnUlPvlQY3NqCPgonHPwLpZGmt
PbFeHCoKEAXeriZXjARoL+NSPPAi2G9JK2XyiVO6Jqk8XnwriFs9aXqawHyUKQ3a
/Zv+IN+b9+b60hLLucRLUquwzFSWFvFcMvCuLpYVb1YDqyjrAyhAiiH/q8vMs0BP
fXHEIYgBm6bReEkHVi5Wc3ok3ljnCQQ3XukUFw6lWtwvVeuZXb/UAaHKMsOTvqBK
E1XGk/S0K335NzqgMU01r/CFSw5xa2JYqEHel3um4ctJ+tB6KQiBKxauACG7JbfG
34TfFRA/uP1iL3+tCM1OelTQKk2vME7Y3hGGOhMrCEOZsOBJfdR4nkl8SoLezXGC
4FfoK6eerSNaXQcqDlJHKk+YRAHfn1iNkccCtVyISl9L2U1OIYJwO1NzIJsI30bn
g75XVx/YAv2tz66HoB10TAdz2ThBC3ZDU8U5vzq6FzS8AcoUIdr7zRQ6b1/xFTOF
M+TMgnSta/5GGwF1/ETUGZ16rhRTrRoogNwLLI9klkudmmlMCsQtISPxgeH4mYF0
r1P9cquhvPZ9wdBwvbRWoYtdfBCByACRRc3Z0IzvKZ19osEP1Up963XSXkAwcV8A
0U1bYd5Qd7xP6b1P+KxtIC8ta9kVDpcdbCKy/H5GP/xlP095oQl8EFB8NZ4Q+ADZ
JWTcoPaYkheG0TiW7/PtoGFsRec0uGFc5KFXlR9FhLCoFVGN35u7fmGU3bDFA3Kv
xIVLKjeKhplxbC/xLQVoXkyZext1z1ivveW5PNxzOnd6V3HM5BImuDehXLn5NGOb
F0hdMVuaPNBS8X/CU6e22ZdEXkFt7kwrxPVzPM2YaMX1hsYk//LmLVuJJj2+dOCo
QOdetX1Fsp1yjh5lMzJd22FA2X+U86Ca77hQ32JQmTvY4eIZrf4HgpMC0WoLrPcW
8sfwPi+Uy+hsD7XS9w5iAJtfWfx3esuQGkxte35995CG//XXozPX2U0zuBUNQPWE
9ebRXrmfYA3VkYPBAfJ5SwsxqrNUOsCwFMAxzxeNTbsQYcDfpNzWXMmB2aTIYxEp
OyOs7M7F+B6iiJn37G83VmBc3MjvkCuqwFEUErFWBj8MQ34KIWWcTGpoJgO2+/D3
SszUBczy1iLum1ZcgLaOLtjIkmdEtTyiq/bCP1lckPiPiWAM2HaVONaaiILe25Xi
OT1p0scBaChDehQmtGt+gVRw7obAGyheszGeCSFcG4D+XSrr7njU6bObMEX1mg92
zdFQfpvAjm4wtF/pSZZDqXi2UzqO8Db5x3X6J/fSCeOz+sLyQtiIweG5vnt4dnZV
FybMzB2FMT+Er40oRT4HDZWLPWFtGDKee2qoV5enezeFv+kyUOQ4p9jYaOnO7qMe
e3kk2+A4N7TQgQRTaPaO6LCnUA6ykjiyFv8yNf/rZHWWZojo5fUyGd+x//e428EY
4jUsvbhKoaha/9J0UdPr6H7XyYjZ3JQ2oPAbjaBDD6dpov4+I/L1a+o3gup3LmPi
+tJLlkgxsT97tTfdQhiYcau60XT7qr/OGh1+3g58mHmxwk35PVAHFuQq75ws8sTD
vgXsvuXmte09qEKb71dr6hSQ59d3Qos+4Bjp7/w3Wfuw6lxxK0td715x5sqfKuEr
xTIFWMQhfML8+c6/xlgXXpJNHrGVmvVdFew495KSy8YJmC9QflDQyAmHX3qItuMp
NIaom9gmUzMVUhdiu6+O+XbPFir9LN1fYl7xNlsUgH0fem8YbJquzyH9IjBKTDHh
JXPnaE9C79mUyBSKYStYwliboVGaBfxlIYePvIFo2qN+uUEsj+bGYTH7h/l02zwX
sH+ry4K6GRdy9PZJXwkWa69UraUWdmr3IAgK7PAQ2POGBHLhHBNXssbbIocrNdLP
+PXPFX9WLtMVHxuRR2AgA5O9hKEkKQNFMLPi17yXrMpmg7bR+ABaALrUleTKtuCo
6MR3rO2/Ty+0d/nXVOzot6PO564pzNIAMDeetkrQu3Vk/lolpABrogUd3fpILjno
bvjmd6xSgNcn2TP8mPunzUe58tsa21BDnLthGKQ7ArPy+Lp8fEpupb5zDfnPKI4k
Vt0xUx7KsGZ4xpcv85KnjjwWq7qLvj+0XYI/u5ZX3ns1F+ClpUHK8sFfBCA4jDc7
LPyuWcONrMLQ9tdnjh+C9ZpNaAupC1UE/T6Dl+RIDYEPHSxwORf+qUABxYuTy9Q8
4eOLBt3JWsYznj1+2yHxav+BtZtlIyfwwX1Z6ZK2jH40DfPEoOnGjP6iV8CzNxn+
QnLERrRUteqy4LT8sazzuCkZVEUiu9XSrSNwHV0AXYxaTGHv44ZcSL3vqLDfRMCe
7aJyfFrdTUmCrvA44qwr1JrqDF/KYRVB8lwDsltyijeohA8T9/6zMy6IlCxco2kP
E2me9J5mlPhe/LPcCuIUCG5qbywyDKNz2nvGAF4YXgpe2y54fOzE6nEAUoX0HaqW
nMTC123oN0A84GdDKzXKfFfZkxnryRRVYWfGCX7V0fpkkbI+YCQQ78i/It36e8rB
iqhDr1MFwgiuEf7PKDvMAR8P/bCTi+W+8V+4FL8kE01T9cDvkJeinJF7U70VBqml
s9/4LsbRm6/YWVKuIeYpZsWlAyu7qEaHnkYipAgtj5MGrOZfARWGu6AvBfQwW3Rx
uLfv1TW7nTuFNKvsFJ6PaSlNe4btf7jHMm81jwl0PilutDoKZZCw+WYg/0i+en/Z
TQQJ+5YER20ChLHlDYaKZlntpi6GLGRenXDwAiYZmiyubJLvugdkhbhYpeIVVpCZ
6k8ZA+PK0JDkfWyk5rdaHkATwkcJuGuAtVQxXRnR/k7AXjUzOo2Fc90vb4ZxPN7C
5djmMr8ybW08P3SEpR6zG5cOO5TpGsccDNtwpA0VIe56DGAVK1/sS6cEZ7nJdzeh
GMk04Rxy39h/ayI87+st8pTfxmurxf5AfUsljWFV5EypA6oSxPevROx8P+fjWhU+
7dZzJeX2Svk1PbSf8fVOhkXONqaz7BEFwAoMM+ZByk5WwRoDKgCANCLbfLTYJQwH
j6ACpxi1A5cfL+Xd6uiB5rifN+OJZpqPSCes9P0nUjfkV1Sjcp3wYqRodCx/y485
J8fvbvRJ5HkKjbuMYnazdL83Nq9rmjKsrwpl/baP69GjgdFVmEMYyIvun1Qyn6oS
TkBPT342mKVq4eSY23yVEG+zAsqsXsOXzP61mSEv/QLueyiPZf1foJXQiZG2YkkI
MtQgNewj2w+VtwrZ0l1CPzSY7dhhQfGO5pbpbcggVru8UsEisHijvFkP8hXUQV8a
XtLGCRSkbBicD6FUpHnetBu1temrxTXSylVq2qICMTW4LM9JoK3awL+mxcVoGZNS
gYbz8VmlDL0odNoabFer1GQgpwe/9nHuQ0IiU8AnWH0dCK/7FfAU+y9X3PrD53uS
sM31PHsi9cyzB36JljpF/PHxn42cYTr869obozNEoiS4X/17WzMmfMR22y9WeqmK
WfTcs68p31KxBArDV0uUuQF9oaerNQNeEIPMDPE1raeJYUKDE8IL4IxqHfrMWZqs
Z8FK2TfCU9zpSaPRYs7kqIT4SC4+AfEPoJzi46iuGOZD93E+46nWqzebsYMyoFys
fmU98kZwcDSd4S+yO2cqlQCrVkpqP7WU/ruA1fILBtEYppe6WmubYJ4e8EBsqJEV
xPKnTKia1CnrwBFIeK8kqIHnfhZ32mLq3Z2pZ9evF9WTIguc5WIfqRwv+vbWzuCs
pYsP+Pn5O4/2sn3USpuniUorUfZlMHeUpLBMmIe8BiPgH/K8IZvB1Vft66TxxXzu
lO6wQtZPrxSs8DHxK0oUz3Y8JMxlqXfO/kbr/4huy/pUUHbnzSEmUe7naPkDvRNl
qNgnE4/FEJRtFOqfGHolBHmGLzUjs8bFpoDHiwqLt1GFDDbArBB5VFiLFkj8rvQH
zJos5PvwV+4iE5ZAzt/Hpr53XU2+2jNQhCglm5WtEGLDEclmXexbVLDm+SBqEde6
Poh7sHxdk39DS0RMl2TTHh0rdx4kMBVIaKyzjAqdsSc9ipOrQLQL068RXBkliVoj
cRBifaWTK1j0DWs0A9kZp5wzjoQg7I7Ifdi/jVlVGb25t5g3KTAvctPNOZbg38qi
S2XG67hy8zILe1bHx9yT4RG1mh5xUk9hPeqbSiecZqo6e1nRrvIYH3PJkqJcf8BG
5MM2FM2oYQp0AvuHD7Vme9CPISgUdhWZRgpTzCaW+AintKR9NZzcEC/MDIs/TvAB
K21r2GMkHP0wU7CC2yWn6fze2c2ShRI6kCvKqfCI30trpD6YLwlupkg0NhFkFX+y
rcplpD6KyFcZx4UNjjsVa7qtmRC0c/gwC98spz2cT2+01WPgusz8fHGmMofMzlcv
BpT2Gvm2cw+ZzqJo1M+DpyLm4TvZxq/qJtHAmj4hTQXJAS0+x54edlDJdL6h5e2j
1fEjcOXIF5e85AZ9nMQRbyjSQXxcVxHGQHEaUYceS9dDeLUNI6MS2tVIN13NeH0c
WTobYRgYZbxb2wnEFQcQDqEaKLpqrmZtaeHagFh282C/kNf7X3QHSKbIeMH+CaB/
aRQeQTmoPqigmrMGVUum7SN7A+sZNrkCQTnaTFc7aE+hObwer6hBuXrbJF62M5xP
7jgJ94XAfedLcOof5gPcJhh94FKo6+lngSSRMpn20lSmEsJ+p79BXDRD/PsV8/FE
yXlTld1vki1+scy973C2SM7wt8yjQ2hDO6hr6ip/yvJC8zeX5zGilUGPE7ynEJ6K
JKlOUnV1rGq15kCDLShOshN2YIHFe+pvXyIGQnE22WDjekrsiDAspqKa5tBHgIge
Ov9Cb4ct35DP611LfJWF3uKGHca/dlhHxT0l1zSXxLhCDX2LUoiWAB3+cx6+3Q/P
5hLWRWqRbBaKqUrBO3ai2N6jKmp737wR4P3kAiqQDfWAqWJyxYyxgkhEoQL7ajTz
wAHKPVJyj54qjOIyW0Ss2fpYPdJFC9NcNXmaNm3UViCAsvgxzQGHXLT0GmyyCiFv
Kb58SK9tGHP2FRntgWLWstNmkLqfNam4M6ifVnqrBpVwCih5kI6tNRZTldUQkEwm
UNjjIVOeKS6PlwAtttrLsl9RS1fWu4YxvXu6pQL3gCeBXYhyEobJU20dEN+sQ/Mt
vn3IMd7iMYDUyP3NV3FtYTztzyQJKvJOotMtCmoZJYhJhwAdSrJLVoenlxzWHPmz
lmVAh12p1D3ehOLJgsaSQtVxRhxX0iOxO6iSAN5fIuREb+BwRHJL7uQmzPwovLvs
CbK8gn4iEk/AE88s4n0g5rww4ULeGaLjc84rPEW07hsCySO9WeqCDcDRjBnCVZa7
tExcZM4ZZ5CZQ8QhRaxW/M8ErxbsstqIHoBl1755sFJLPjQfVKZb/p64M3DGdckQ
owDzatb0a6pFRpcVkPJl1CkabtoGltdyAa1o22Nrba9zV4ArSY6a0Vnq5PzjAPxr
86MYs1kg0Jxl0CCpKstU0kAflFO90S1bRPf5XKnyHXyvxpnPGB5PPfH90LHX+X4E
8H00IO2ZW7OXXnnxud31b7HJRYcNI3UdiZbtMKH0v9f5N7pE3x4zhlot43G8mJwO
qPZhI+6bP6+PiKRAKKiKVNbxJE9hnfkrdleO3O4/XAgzSSoAaUQlFkjnSYIJAuHS
6E27E5UDTakEN0HLSdXPHP0PX7+VW7V6bLeUqV7UKAEoS30nAcIWJFMRiup09Z7Q
p8D3ljRkikANfjsV/izuZIOB5o++lKCjWeECzdp5DDqTleKkezo+vhciVbltVqvx
CkoF9mWU3X748/RReBtBoWIF5wCRH6dVk9r6VlBny1hMsU1qfYXFLvZsQob4rNF/
V512tay2yLXKiDUSP2HcBgW7rwrJZSjrDjNcopdMVFubF5ln7odpHK7F2SKN9FAH
wQkfiUdAKYwQMKKkQ8+flUH83F2LJsSTjBfTMRnhPsG3y6osG6YGP+WAaZbEghYn
HHIvWHMKkr765CZBGriyMhlRtlT5EebVtwYB1EWTgm/6A2Kwg1DxLURsR0jEurUo
dO8HL67tCMyecd0oFu+wYtgVGYFvWyGbCArI2OukCdK1nP7swgSJ4gknjw9yQd+E
v/FUeAez4x0U9gYSRW7BmDmw5mlEDiSpa4dRzUqbeyhbXfmSKsJvUmlY2O6Xrd8v
IxVSy24BIVFlhnVc26LBUzMUcI/FtA56J13636QBzAzl/YUotWTI5iKL/HQh7qWP
mTDUbodSEJNVTelxKhDabftxb8hXV/igqb3b82oTh4P0qowZ4tPBpMv5M+qg9idL
ABDdCAc8EZuK/QIg4gjH4bAFZ60n0JAMjlr22siXWjaZqcuXDZ4wQ+5uJyKpoQXO
oDF8vK0SrMnuITNCpnoU6GlksBQ/2eeGILEQwwI27ZIPvD3aerGZedP0U7q2lNEy
Yg0rIvGS6xgitThB6joMZimBz+PzCsUgCQ60Tfafx59md7TA1kB8DWjqJz+9Zswq
vDDdb4Xc7YxuoaukIR60stZz7JvK9g7MU1T53LGscYSNE0HIO77X17+JvLR6PeWN
xmg7gXNigS641WFKP/IekEptwAqk+2nJpP7Dgcf2hz6vL3c7A4QQxDrA6xMjcXYy
ac7/db0m2a01T1Ql9nS9Dw2SWcoxiXGRbJZkAdb9bQqp8hs/92pP6/LqZhYXoX+T
HjzAi0VArGU4PgqrU9zH/y9R0a0NyyqczS290+0u67kcZSVdazle6pzgqigWZ+ib
6k11VkHKvxcqHfFaryA0oOLVWkA+AM9CGzIdg7DU2JuaPMMcCps+AIK/SimuWurT
XkQY5awfrvcw9xV8ihzN36ywspeB6GcNkXN7rHs8IAKj9Ai/q/I2mrIByehHhJxu
wEAitpsFAppip87T+ob1wGRmll7ZksI0Sd440tRlVUpG4oKSlTwU3YoDzAJ8Xq//
iqaXsSm4aerOfulW3QMxTRavYJG0G08+8H60U1uE8Cbog1qRljkx8WCACIjKVBkD
DTOx5+JOB0aN/o5oN+0tFW2QhFRT6tkTm20cHUSvFXdgBfeQCze5rkZ+KfgSzEIu
yrnYa95zatbKmA1+RRrNUDLX9xZXchWmWxTxB5pAgwCDnx4yLxITTfE62l5c2s1b
pIlDo/zVh4WCjJlD7THApN3G9/8IZ6GVtZWhelO6bQT3kJ5S2k1yRSJQ1Pserblf
GzwqtLPwZSlLT34M1LY9jSXO28J7uc1e+Tt/yNaoT00l0BdnQ6HvAC7RbuFRIHvq
QdX4LCGay8EzoBHp0vLyq8D/7AcuP7IakL74sbXHPXQ3wQBEabp4BMgWvOIAbJcc
HRsSWqi7LOd4BSuyEq/ZS/4Q+w9ux6kf4DncyDSv9KCdwfnLvhGOEjFDHiWElY/D
8cORPPa/8h7vtnvOvtGRiXLuwh93TAsR1cWFnlgxtCxCqQyRTq4WSMdJo2HQPtZm
OSEA5y92QdqdQGDrT6hwOji2BGOP/2HZ8ytCwpL3ObrkwRHSSrRDE8TLYKsptL2j
jhjFUZmhm/J3zUbNzMEjnaLLcFCBAxp3vtWEQJ9u6KIk+GVCJk4iZ834FH/ayos1
w+jArsuOuEfRmY8eTN2jQqJdnfbRpAl7Oqo2vzTzMiL1NRJppKeiOibPXepd2i0H
i+hVm5sfq4N+4nQVcgVEToCW9G8HFMEpPfNxu/0esRGXemo2O8JygoIg7GWkE8Qf
Li6RRSWIwTVhVX0y4rOc+YdoIzVlHZfVUOt3eVts+y4o/lJoW6XflywGb4rLHUvn
eLPh2FaTph3RCY+mNM/G+974uZ3EyocBPRLRkpvsxcSqPxwKKg996awLi1Re/fWw
7JKVv8n45fP6v59DKuVmumTYaxbASIljCoSsFbJ81E/tkBb+WqZDsA4RXL4XJEGi
OBhu0ZHp0o53JBDk6pJk2EnS1Jw5n9YFu2COWsqkVS2QkW3u19B3ECrDdeBCGlAM
Ne9ZzASRd1DILyJ5sCBynEmoA92tW5jnIRgckDA1mS/rNjXeurc/MIh6Z7FbksEk
CPdjAYJLRJrHkAAB+8qkKJ3HQUqg1h/AgGhpsnJ7Ar5PzRrTHE76de+bkY8Ebcbm
VKZkc2Uys09aVpnpDEnNGnIR35XFTwAWErswJo84jk+3nI1n4nWQDcfr8rvu6GDr
oWIWJaNlem51PAvym+GFksRWA1VodB1pSWjOlXdpO50DrLIzFsI8l+DVh+fTvXhb
b4DrKJEB8wcBXx1z+DW/5PT/GIvuNWkjZjDyF/VJIZ4+R5bFfqLXdmtk3QEfgsRA
vbOyhTorrU8Jidxh6q9L0D7cr0ytaF+fWsSy6+KIHnSjftvHMl1PSzVUHqZKwMWp
k8y+ht2hLZmTsCqaLaYApxZG5VLXrgBa66qUSYa9Fk4S4qq5bP3fOxP58UK2E0f2
8MIH1sO9viWgn9vMO0tf/HKlxs6/lnwMSCvpj0m1jRKdMiu8iXQnbdclTLw2rrUI
SaVjS/6WLjWhN+EFO3CWBRWsWjlqDdDdJE1HSn5DMHtaCOI+bBkQn4yXtqC1XxcL
vnksvgNIWgEfZDDdSPSrLDQ/BKLofCeenHzJe4OiNrcHnHl40NyyTp13GLH6RAxl
RA7X5XJuSQo0AQwLbHu/jnnX4paBR3Zzw+nsaQlv4bJohVHj8RyFJdjyR4qkcSPH
5sk+98guWfcuGX4djZPTRNrmYok++nbeSNPUNarYk//NZYQj3dkZbGh2Mkf8Grf4
vIKrqSCowpcNy7y8W3SgmTYPYjsdrSVJpRdqyovfo1uFVYY+icslMF/YFyxU9Ojh
NBFqi6ydF1Vt7iTr9K9L5Qk+v3Bljo2YgOidNpZjSeteYXRsiKsjSp3X4mxBFUah
YWrBY4rqrFpyxNV+uXTaTIaXolN9L/XJ/9cVEbSnXfVTtDjxgocDjM/i3HWJwb4Z
dBhdEopAU7jAqtCdlaUXlt6JYKw4AzotSTN2VsQVK9G0QY6RKrZADTkHPn6Jrt07
bkmsJIqcXZbdqoN8dGtOfIZBFRbO/10RsDTX7zyTDV6BRcLB/fYxvi6uIUPjLgLA
Kw3S6ycMXNlNmbd9Q/0s1cgL/MAxEWiyb3b/mQ+RUmhWxDNzA6eS3Bl5sW/4zqZd
PMkTHa7AWAgS5IiUD5Os+H3bsoOr2+u7UTqZs3694adtO++kd0dMflOJx5D3UsaO
N+hDrtwAblUFMcUj+BAFXwB2OeRGTIHAR/by2KAZCpXbiMAINFKcsN6qfIe1MWyP
IbloPGzmbUmeMhKRN4XItE4tn2bBAJ3Q24yCoXczcKY6IV7OSj9zrd3taGTyxKa6
lqXwYRxSnT80AggH8Oc/ohvKNMOJlA0E4QNJs2hoI2EnmKL2tN+OhjJRre23C9YS
yk4A9eOq8F1fsTtG8gznBDvsOcyLzirb5/553ozBYOwx7n8jduKP9c2RLx7M6z4i
UZme/70Ah/GdkCKsVW0+LBKcNlZk3+eifmh8cx+N4iZQqUEswBoQzAfUs+sdPrBZ
QLFzBn3xUNvp2QeUj47561rJ6csUBQAX5Z8JPH3ReZ9gtf3B416Z9vyD3O5ey/Ht
pDM/BwNdNcIuGaLjUEJIZAQaFLVBg4kfeLbzn//g/LdFBT2UHL3ytcUECuJfGXT9
CR/W1Vr9h82i09CsA+vQiHJFh6tl6icBSDl/CvBuPdC++1TVzCnEHlP2TPu3VMyA
ej0skgtJhpAn+syW8jYnXt4xgxGCT98CZMhQ1vhAKkk7UQss5+fZLCAD1ARdYL59
6TzHnl4s+502qaUYI+G2Tm/evkixtCU1wgbKAzAkoGu3aPenbVW78XPG7zlxI5jl
8Vziu9PGqW7eN6yWdJR0dz45rCh3mkNovF2QGn7ydaFBmtQHH5T7mFsOf8eP5I8M
jxWPBUWnABvHMjO3iTTs/uC0NR9OtrPfeAiUSu2IHf1nBGlWTKR1qLUyFt+hkMYU
CqsmdjNGmvP8xtu/7JqUdRwDBzFOLkqCfuz7647R6+1J6JqjHooppY9DpM6jYV9x
DGMTmpxYAABj2MhOXhRiN4YPfHJYcZQKg9b+OzrqQxDGTDwbMHszHlBevpjT/+GL
9N5unsXUpmXO3oqRGTmqCGVV8VpTU8136PcdD9oUaxTK/A9RyETldP/MVqiQNEpY
Qv91x38RgI/QQ+Qn2ob6rpQLIIdrqfM1KQ/xhww2S1RRZTjy8yUaDtOCLoZdIHjy
ELxgYFB13Q3xKzBzUdhuwZplTnvS32KOuFaAwUXfIEyD8F87UicNtW4/ODNzqEqg
v8HtcOAiNetMG9lIhgBCtH2G3p3o7JYFemLGkrCyqtqQJQES0R/TuQOb8o3v7Kiq
jQu4Ce1bSxhGEmrcfjozgWfWO/ANy0EETQn7fwcVMj6YmNS3vrxMmXGIWjq7PCe/
UNSwuY3IuO6jYbC9b7T4qtNxRQLeGtzG/ggiVbuVGsjR00EToVT5HPGLScQ3xA5A
HiT/GCke5NObUa+3FFd7MOMxv+rgsVutdTzw5vczGR+RuvXBvtqGU615d/Tz76IM
6plIQuO4981lyE0gQClAPKbfN0K4JFymNyLRZSI6nhdFIjSFRVMqmn7V2kvFP3CW
BedteiU7aGpLLR2RG5uqHab8Ln88WUK0DnAm/Y9hycpabdBhuuo3J6+NC+B94END
7r1KhMDoIzci8wp+Fo/m3CuC+BpHbCmYSGwlSNSeq5ofQED8isGIOL3b9GsCgerk
ccw0N/NO8EQSdYIy0/20wNMR24HH0iuP1uZH6IdaReIayXzSVucL/lkoCtQiQ1U5
SDobiR2p6m2YRI4VRGnO16Xje/o19Snt4nSbcLFAS39ugzxbBczcTvwtUEP4u7H7
YJSN3oE6KrMvlJ78aoMD/3WiYhuPyUlPXYdYBBIOD6jJASkm4ulWok+xADjy/5lu
/EnlNcOHVAuy9FYm9rlgo/TsgCbzDw+fhlkLTV3N1FERlBpfW+m2CwZ6zLdQYdj5
OWBMdAtfNspcckg7G7yzzRsDhUkYfJUwXjK22l/fn5bKlze8ijqe2T9Yz4SCF9+d
Wnaw5vOyojRj6iCVi+gEIivGZ6a5xcYsi+NqcaimSN8ce1hBPLtR5B9l4dgdWud4
ZT/r1D3nHomB3nvq4OeDaY03ovBixTSqEkF47JHXsVf6Am+Wde04WIh+9L4sLA1P
x1UyL2VB5GKvYIWfiL5D2PJ9Z+zFVL4FvjPQdb3qXtQDLFYR89d+ucEjbVVaLDV7
8/4grNS2SMPn2pys8epypTpqBndVf5TQX17sfYtZmYIvGrdQQ6KY3FOwPdSwLDDq
El8/C0qNxc5UTp+WqWbUwYnocEi9o7KZoCWwcP8kPFEPNK+fd7cVIY8SSgjaprAK
GxlPl7X3uFjt/U5mcOnWnDrqeQEcqLe5YVkO8HmLTs1ZwPPIEXhOAVrlJ/LSDuI/
mvWTtL5LOEkk/pK70Py8f0LtHFdFHTnFfOLQ/jWtxpNsul9rxaNt90hf4aCno+UQ
UY5NLF/iugWPrNjLyl9dicN+EgtkwhdASjBvZTPlKLMPbkcm+5uCb7FttLFG5+58
7NfAuJsc2dFpSSIJVIyfNPZMxHCRSA2zB+e3ozibHie2AezAG16fPXPO7R8nFsRi
1KepzEWGwQxnVjNEW0ukDVkGmaxN43sHz456v7sHTfv5gaVpLTbgCeZW/2aPKwD1
zlNR+U5rjGNE9X7VnqoFdEd6qMwXc+/5kg22wVrvQdcNmVK0Jqb1I2fZsiB5WJBG
kqwNU3jS0iZpHoX2K6aYSsDnAiz7wh7Gq/09uJxafhV7R5XnG6em4FHBL2mrYrK8
A38jak/T87k0C8F3xSf/Hm9b/wwoahanUtJl/AgYuJ2h3LWn2H0YqL5WwXYs4VTI
TD0pImjYuihOMapDNnT5K1+FlO4q8h8OInE+IbYpVqJFYqbAtQySXHgYSQv2Hjfl
rqWl+1MCiuzPkVixUn5Pc3otK+COLAFnGHucwyGvUtrBmObdQ/GlUPZGU2G6oIsx
KjPvUioKDnhiTj2IXQ5KXalqO38zcDWhGQD5WddmiMSPm+w4/Yoh8wl8D7NR+tC7
mAyS5yWoIPQhUkBi2lEO9U+I78IlQCbQrf0LWFGS1/XWXByrkNLyjgFIa4ck2P4m
XtOof2gvAU2Ym4v6jKEOIpEtG+6i+878SHPzWGwMRTeIPjLOGEElUH7OoXn4pZAp
/UNAodCtnILIT6KlNAFQPNCiFu5yd0p4tZHELyP/T36jqMerPhDTkgj2Dxttq10G
C6oMLHeRwRrcZw+RT5KscAflBUK31CDzADtaSDyLlYnaxpO7jBLioHjncpxSfjX6
m3PM2k+ZQTXepEXn4J+xlKAajH1Tin/Lm0ZZz1zm6I9P9Y3pZ/cg0zY0Jz/9hYxK
XMSPB/+ZYzNV+XpfCIVr9KG551sfw2HkTodcwa4f/3bm59YG+45cMePsyRFYlOPM
pfS5O0UahRgbILX1y05nRHNmhN6CZNeFtPk6+1sgDnQf6mnzqywaGQdAB7QX6+li
xsVrPvVAGTDUQLVc23As9HjG0Wv3kjuv2ZqNP/dL/suTnrikgMrdHoVPUPR/YytD
sr8ZgzYFkOic4FtaEEdO0eLao7wp5gj7loQEx3zVceImFCERHQRVsQUB1prTUNGx
ktLZNYkB0Ip/ESVO74CPW4m2nkjJzSK89yFHfKQCqVyQMTtty2eZcFtdqtNS9oaK
IKmnfdJiWNf/dNpfxaAONFkA1MKfQ6ZlqtqQ7vui0jXH3DkeFZTov+S3ZODtYI3L
bOyvAk45w58ZSEv0HoqZQOT8Gy90iRhZVp0RcmHMex25d7JrS57egNTCIfJf4Ius
K0+DN1eVByFSxVNJYhNOw3bb9On6bE3POQOldyc+0bOUXLyZ7rjRXm03TynWRsPU
H6XK5DZ49vOzZSNFtEXpLnOI5NFwxRXos7lN+c+8SmUIiuTlLYNRH/VcQPIaPWZD
DtP+3QbK0jp59yx9x5/6gtHsThmacKJHGq7CpcvtMaleX1ktheunejSUxAiAMtea
3KC/6d/nOI6C/+RDwffMXSiOBcWtMByDyjcA6HiJQa69GcfTdTRqO/AhlTty+1C6
E5HoBkeQMtnGYLgecrQnFbKHb1vYE3EV4xGj5dDnLsiv0ad5gBtCRCifVyac4H8i
Que6xGr5jlIIFK8LJ1K/aE4yo0VFPPjPoDoBwDKJAoBmNmg2UhWqLWHhSSYRvcUD
LuJxNjsyLwcKE+LYpbNu0zDdb9KzW89ey+4CuAJg+U5jy3L72lkHmiSFOP6rJa//
7+re7mhimUqalBM/vpypOT9gsRzVGUcVWBaWy6/jrj1LrU62A84NleK3vMg/HBRz
Gtw3desnLq1Ll2IhiUyVUy+uft9YTjkp4+7aqAAkuiw3G6njS95UEuJrz27BjbWO
Pk5ygW38Ld7v0QzGnujZNWlN43d2COfXzbfCKzdfhU+YApkpYpezAM3k/KbNpQrS
kLUfMsUfacAw7L22wem4E3FzzoUC+otP5pI263TzZ2NI0uzUVIHuREpOLM80HO70
Oa1g1xqwwRH6H7xEtoT8lP7RowcIel5qIzc8yzXIfKE+2fFRQNLmsb5RqhsUHhUp
tz6QI/jqWlONUafRphTdR77O6455Surdt9qT/EuZ7W6gaI7HfO5+4pmte3R1H6/0
AZf0HGiQYdi7+NRnV96xrnEvJ+BoHaDCFP7T4HuXBnCeP1DkOet76sh4rGkxFVpZ
GkMCog2yLzqnN3wgyPpSRh2LnAPikc7R//PXS683FSQRFo6+nPXBxuFPJG6myku2
2Qw8NCiwUjdoj6/b1ZfD6zuIGMl2UAghavyzrweoJ50UhgBnZfdfUTSW3Z4pSyYY
j2ObLzPPwBmPQmBijXic/Hu4YgOs+fvN64Cs32e4UgVJEs0aijadKtD6Pe9+ENFO
Eu/J0SgQHg2+OcEYwCB6YC8iMh1SLkLul0vWsxA558Qx7PGZq59j3KDHLqE33Oeg
UxZGvh9kXZ7CV4GKsdff1EMMtvuxS7ytWpmyYBfMJ9rCyU8RiPqSCSSSINCBH7BQ
DK/wrgJL7p7jAXv+q578hQ8ryj9HCW1GLb2pZcuFBE0RCpkO8887UUbNuUDWr259
zSUn9hSssWP4TaClY7neVD/zYqEUKKSY2dYhGRegl4AEGwvpMbzw1d5WfHjOqioX
zGDJugGv+NZfWzkLaTPj8fK/UQjwkrNvbk1lbxlOBZEfkUgCracFogtqjYQi6Z7Z
RjCMV2cUAaKHkTQ6TUTKNYksyAZ1aSy15YTczLCm7Lh8Qu7xYkfTDBFBiP4uMtwQ
Wk3owKxTylY4s6ZkC8J7K+xa94wfxXBr5d8e+peI3aSakIQCqwA2rSi7wu8TRvoA
wlbFPZAjdOqxiX71jaHmw0xiopPw8U55CNZsrAGisleHAjKK4Y2Eu75a7XqXbfMB
RW28RUz7Zh0TBYweRMCKEku35A994pMtl0pEUx9M981hoV/U/DrLC/qy4hJqHZDk
7ZTbZde1gzZPp33duyylp35a4/IHefbfNHCQKxQr21oCa1mOLIDVRnJXeTtfgZkF
BAda7+jZT4bC/r9JPClnFne+BXUd0dp6L8hjxfBr/Duwmtoku0vqcws4LfQCF3Rs
1epASyhZd3qVFLzE/kyLjApMrLEmn8TMX65Xo+FdARxsjP5pQs+tW92kAi5Jwhqw
516OktYQiv+geaM1tDLMGVh9H7QZMKxKCbk1wg8EUfOouvaabgv+BIV8wnWPII0T
kpcUhlSiwE31Iw9epcXsarbZzgLnjtYLlLGDL7ZMZHhFsj0XcbntlPLs9DSTH8ez
eKIp1V2gjQ6BQk5scX1/kI9SCIGBYWO9RxLv8tZpmJfkN5OCVTJ8yOyDD9IleJjC
7NlKF1t1aqB9GtaPxDGWNmDPHjAAXipXcmuMtMw6qOBSVk6JYe62cjaTL2lrkRBR
al4uI77rwI3izhfri//4ziHpjRD/ztkj4IAlIQSD5je0FoUEfDO9Jn+huUiifMbC
Jgjp/d0CpsxweRxl+vb/+91Sq0wLhBNeg0WlxNa23VzVI6XtKYFqIWrT+I5/1yNG
wMrmEM+sCguJMsQ5wPvefdxOLmHCBk2lnDypac1RBwtyjlJBj1QMCPtvcC/qnS8L
dMkpAmgMitQ30qjzfYWGUW4aR1J5zGV1l0IPZ9iSAodK/Qltf3MbKS/hXqgiVvAu
WCOu7Q5Uca07ImqSDEOQA0NIMmN4FY6qeS1Nviby0Sh37gMD7oaAnYUg1l9sXP4C
5q8Mhqxh9EAvCohYGkccWTvqxctz/mMw7gqOVud0DEIs+at3L2PjSyqkzPZf1ElX
GYs3QRaoerNZxNamuMXwIMV78TMEqC9JhwhdIrjZj4o2Qtn74rQiDPfjIHkGjOOC
fK303UsjfGAoR1WxgkqoYm+b9OG0PEgdx89DnFUfVXH2KLOwCJJnTfhDcRrOF9tY
1t4Nvi6dVc86LbQJAnABTr746pKfx4F856aeJcVSV+IyGcc09Tbtq8hx6wtiCvM1
/US2fZAomK6q2kct4fk5hLnB7lKoFtZncReVcG9VbDvT8pkerhd6EqTS0vNviJ/N
PeOH9YcETi2z2y2B77WIaQ4gDazV1bghrYm8U3ah/Vq2Fwx1kKSiSeKRJUr3N/GM
dGJsdyK0sG4tfLD5oWWnG6wCqisjleU2hKHyShOSfligOHnNCNiXoRv6qyxB8ORa
Dqz0Yjp50Px/0tYXkWjvCzaGxgIEwX6P3+XyLNYA57Nl9/DzBt7ytVpQKVZY+nvR
lqQVMsndbhaXQputUjO3YQV1eAh/n8jr+u/VLpat9c0fT/wP350Dq1a/7KAF9Fn0
NjtDhRZBcb5ePH6L+o1OU59/+wbXt+BAfAoT6S5rWd8fvh54DVyd3sYKnHGZko8V
azf1PDfhHTCVSepV+6clG3/sxwV4fpWQWrzhf03GzYVBA9ptzdk7qWq0aZAmIBpO
5Aq/mDE17UMzojUz8xHjLA20biGt3HhD4d0hFO2KuBgKKy1bggVmp+wtpo/FWuGH
AZqSSeeRsLV8WmVVXNGXn5mgKv2BWfAS2QM/bXvXL1c0nDapUxz5fhZVbvsYMI/e
StKO+fKRivvypBV/bfhQn7a3scerfom5h7slC9W5B8BTzE0xnjcs21eLuTCa1jIL
dLFM9VTjcrTNGc7VXbzZjkKfWT/WxZHLwK7mEjCjf4pVSVqRbcr1mk849aPbx9+5
Yg6FjHvz1MdnwHhicKdopXS+m3UbJd9F4mE18mnI+XAfU5fbDH6fjxvt24tqM2uw
LgGgmzc5wxZoIJV5R0h2u4NpRqodul99gy6l+Xx6HTu7CMlSp/rjyG/ajW/sm/Y7
jWnJfqFxHgo9vjmxhmfX+0TsM+37ffeWNXnqTQrIBsGQgbve6fGlkyABBPVgZJ4K
B2vl1Jg5epes89lQWXcwRCbF9mbi2nP54WBC2uNMfEe9qPjilhE0Wub6SEYviXId
LNXg81dIeU/ynKT/9EZCcaFvF9KxjtTqLL6IbwXYDTn9JWgqEUJatrqoOLTsHjaX
ICHLfMDGkre6vy0Q49qSE2rcZwZqh1DX/bTbshKc6uu8EcOaNnYN22Z1Z6TDdbkl
GE6r5vwYiVkwgOCKT7nqyj5Rd8CsOKkCghkSr2OBnkLt9hTSx4TPvK1BEcswb2GZ
gYssD0uDgZ6ziS3J6FCLzU5W0EMsumynczVnivuF0EURvIQ6KbFKNZcE/otPygjA
Ehg2rJqn3d+rjJyFxXlOd/vIBsu1YaexGJkkC9zGxxeC/Ff+VFrGvdOd3VQ3DXdq
zz3dQI3sFMS5nq5XiIuykZxKWan/UOlfvQ5mvsjKzc2ypy0vNe2Rle1LAWZetzNF
W/PlOCK0olWHwjSW1+3IM8B5b9rQzs1H9eikLcTvvwUZy8qaLzSzIZ5I2UTwgt/n
9TyNg9uR5sJimQiu0SzCR3yeqDqUs3s9BYavMfMrAGdZ3VHRcSKAogNeHuiEZkpX
8oP4ZjNDDXkXKFhf7jV15yy+JfGSL0vZlXcp3F7xS4v2Je31MkxIQjxFy0o6KVp/
FDWbwSMXT8RNR3ozCh+Gu2IqQZvukHmWTSNPIt6Va7lk8Qrj6siV3Kv0OS5qxeHf
bcIabb+DOp5l+HoJckf96ZRMGO93L3kolt1V4xD+BtngHwzHMNax94FgEAaOJsBy
/EdNGKKuvwSsfE2+IKEurGaz2r8O1AQusvb5lYOjpT7KG35lciE2a0BDTVF1fNuj
T4Iik1+hQ55uIwE74VmaqfaePV11/cqUy0lyYUggNs1W12p7uJ6ZMTTXSljvQM8F
yw9/EWo5J8dqdQ0LbN/lG/iwlU8IJ71EofBN4TZV7N0IGb5FbHl0bzzXtsFMlpwW
TEom2aOqMeJs+/PHcTxot/Q8cBKQ2e3YQiaYhaF062m8uW1ZchmRiwGpbimyKAzK
IimeRIFC/52lg/17kVz7/BFLvlTgVWxwf4ccFlxKcK7zEYgS1eL23oV2BE09/ZN5
y351p1EIJa0++I0A8/iMNcYUSncJgXWSSQQiNrbq952zmU0BOreMohwrlu7bjujG
/SuDhXyDiy4ISZ9tA+zv9hYIhOCcm2L11z7euE7shKgra6+LapbNhYKzohr5Grex
zcSTgirc6CRgAJNZbWKoW1r9fJIcPZao5b9wsyXk8So7QWSmjNdUEUjfF9O4z6pO
m9VxQRwJRDyefFSsTMS8xVw7Le0fMIaG83Tf1f6HuNfrLDbcx73XOdGvBsBu4DKr
0wU9GQ9tzzf1LU+zEWG20nc/ZxCF50SutYplKsFXZgUeQGXt6xfKXcZ/NZTZdtet
xUkICAI+bVQ7FTEz1cHHe0NVCnRqUl2yaEAUrObY5JDw+nd+N10mD2E8ZQZLowGd
KSK9YNlwNKDU0CEkCjvxHEYzmAauTXNoBgfT/JEODFK3sAcQ4SuDXAhdOAAPs/me
l3oWAZBNAZBIquJkYjnPS4ZuEAGerj9wt2eMshD5ls7qO6/VV0CbMTq/0WEKkdls
GHK+4j8gG1X4ju4QpHLRbGuJ8px5Z2CD/NbSbTwtqxoySiNIRSu3MsDNoPJ6Uv63
e/Sii5pqm9B8v5AVx2+e/y3km9JaW3ufZXlHfqWoaexFaG+4w+RsnAk0GL7lS0r6
Pez+Ntb2H31h4mkSK2HuAZn8IF0ydHqLWepO7TaCJnpII7T43ta1wRHV24UCt1A7
F34PCzjl3irboJ/ZpLeRj1+RLfpSgax+pMXF0onM5vpZRwQZyDMXptr43XSdgWDx
L/KUcMcHngDwS80bu/OKGo/vufCNQDjNnu1I6CM+ZcNys2q5b+aNZ9OVmxwcggp7
tyRWYWfjTagYgo2RH4uVVMcaPGakd7XbZWlMTPwHqO+q0FbHBWSN8rBOigMeHeG4
JYmU37aCXL6ZlF9TQBoH/1A3xE8WO2ripAoEarSZ/CTeHWC4u8hskEOjLNdnTzdr
rhEr+ulJr1vj4CcE+k05mRM6z/d5ohIVetuWIf1pe8p2j0mh6Vl/r4bt/3S8Z1LR
vnqKQ49BcVBryQIm9EGDgvgc0dnyhTG7h8lryTiS7bHWtRca9cAkzGBSZo15IVbO
HW/yAXrcXvr/NcD+FzZ7/gtTCmtPOEPoVhrnmXKWZabdsmaMLOYrdmLgSWHW/w5S
H5wUXW642QPUzPV0bJFz8nX0eRHrPICi0G6/kDX2iqdlYb89OQ4MTaMf70DihE54
qLyc+217Z9YKUP+pn3e/ydv2E8DgstEGZ9jjWfCErMJVXPHqsp6Zs2xnpZ5rA9IO
u5AULfnarTybVvKhoUTll+I4KC2E1OD+Faz244FmeE/V6BhZmtNnhLB276wjLGbw
J3kFuHtsTB3rUAS5MwXQ4AYlkzbDUPLUbRailZFCYtmnXHdaAgoUi4ZO7nZofKgw
aXDegMdUaFyyki5xUrqn4M45wUtEKt17ZhwWdP311rkXKWgAeusuvqTX6eNQTiaP
B6ML+oABI+Rwzg/at4fgj8DNGAuPb5taS449E87LR8QsymgmHMIR9uof4KojiqNf
frKSAlZ1ezxCBR88sR0WWjXe9TEJ5Af6J4k9ivsYkwFSOIOQoXfv5D7K7eG152xC
HafX0wfvx0X7MjJbpb+6tVxYzkMKOkqRs7cFo1PaaJOq2xYWYPQmB41S5vhe9me9
b6KxeCRuf8JZucPgj1HeRSPNk4m383V4rbeEHSDJSB11UDg0mOrRfAs88g4O5dVu
mWOnAC1SB2jxbO5MKOPiLk04HbclRhcy+hj3kr9LqF929cEE1jHgcnY/3MFTxiBy
aDSCgH/GmMj/MqcUibIS/pnnkDR+eNP9zGhDKfV7elfxFu28R61LtdlZ1Csfnu8G
A739Xptu7nSkKGPcEkPO85cPfdQYDsGeTBiMElgwMLk55H/Yb2x5Kmg9uYiwufOl
aY5r7XqyBazWGuwN+hJGI2RbanGQ6zdDygty2AS/icrtEZKFxGmgFylbc9QK2RKv
/Cpeb1p+vFHMeCSYIxEoIi5pPb1OkLQhxqzO5Y/aHopb1oTD5pwJtdxJRniAkVdB
dRlocP83u8ctYzwVtYqvOdu3BIN7+KsOH5FzgURh0zBnG/U8fNP9xrxaaJ61abw8
Ynjwp/x0kPXEgBGN1nZ0kctMMW6LdfJ2NtaGXSg+UMHZw51tf0zjARHoxr5hOVPQ
3ZwBNNgxj1oMFAdoD9nQqqI21lgg2zv7w/bpkJiZNYLf5RJpj+NRY0IRr23KWV1c
0B445lqSx9z+OUgYTGB6xnNmSucbiv0I+9cxUUT6ih6JOQCnUvxDU5W5KhBY5h9/
YgGmXYKjJ1Z0Phks7lg9jcQiXIdB6DBGn/k8UvCYYYTFV8WqXrtsmQa/6XJPe09L
f9nX27v9g+0BRFmFmK+lp8+YDvxy2fjDZKbCQxDURuOAH6m+CK9PWTUIj8PzFjEs
xnWuhswSatLZWPPiQc9tFnsLvgR5fEWa4/qg9X41ZL6USZsZI4ZLWneR7EYWXifG
3dbVCHloG1Uh0xLtoM2hGDdxAHoRIZR79HBiyHBXcXoGUkpb+JHjW1Rwpc6TYXKB
FAdlA7ndAOz0h70BX1KdaeXbWy67ME9LW3aezKdPFHlkpdyU2RJ4nvdlclE/6DZA
j9dHwQGR1hZ/msEh05VVlacD/f96IhWrnaMJXojq9kiT6P5ANmg31AsOOA391BwP
lZjd8mL0bvlN5oQa5zzO6LXT4zDy6JNXIsj2LS36CxfRf9vOmXB78p+B94ZR2Io5
4gXYjRZIchBEbueBAn7c1/CJGA6+vGKFlSg1YWV2bGOVbEnTM55wSpFmm+83wxkm
5Uak/7IbMPOrs8TQuT9ykjFkZ3MJlpEOUd3US8m3IUoYKYF70WDpMRti1r4/e8vR
ba8vT5kzCuXVSmyfVExrC+S8Mrz0oDPXxCQ1l8J30DVfHrcfkzNdpi3WkhvJm4uk
IXR3N0YAll3Fo0PYTnRMVPxCukQFa65D7fYpFMJB3PSPUgoNBsNEmQtGbBRXLUZH
3h/k8D+wOWMGCYV1ck5qwhSF5JIHV+7W5bAawcWsumih05RzOfGOCykMeWdPA4y1
1Z8lA16Uglv6uPFOqvNSZtu7qz7itMztXHY/L8x+265nvyCJ53HwvWS29DvEdPLL
AYEV4yB5zfIkmPU12XRc9w1vtJlCHFZUlRAoFrXjLOhxspb17Gci3xFT/Un31gDN
EetSDJc63iN72EmCHtmh2c6GAWCcTOjE91/U4yVLhJlVtNXSRhqPSbElbzHQahCG
qzfCUaz3XhJQdX+Jwjg4EspfWO8YVNOo781mpc/7bAPIgGuszQ7k1/GL6DV23xbB
5L4nqnTW8oWDIRzNRYCJgGiMZW2xrzr27OfZ61gvTEMVt8PbDcnqTcmzqx32EEBQ
U/qjPGBGsb+iTM+ucMaAHBK3GkUux3T2cTH/Da2ZyzMu8P8Q/R8Ylexe/1tpWWjF
2ynhCRcoQWtG/yym+bfh1sMLdnGWcPu6RT2MFUFG90Wwrt0bv1fWGTHfIdJACz+k
0Sncc9u3eqfugEafGu+49CXyAXnx/wd3wphoYRQK4eG61Ueo7X8ypRU9mmPBMMtt
AZKhyubQAe5RdphxnbuXrBk/U1kgpxXTRriAyOpj0apei5w691JUoausZd65x9WX
eLuG5aq3aWA+ItHJgrI2omCc33jWzNQa3qHhwO2Lk9zRzvlKgjx9SxkxI+GMaX97
y6ZS1yG6gK/G+0oGzuLGx9lNAIgeSU4ebT4kK+Kd8P8Vn+HctLd9srExGFwX3hN3
PkJw+92YAcjyfpbaglen5y8yfQt+RT3pcTt8ScOAiNFyt124rSgp5Wt7ccP/tfrl
cgmGpEsJxlb+TPah8e5Br3YhDiCy3Du6Pl9LiLhLTDQkN0mvNAJo4KCfX9KXvWfi
HfTNL37KZes8JvVKlsh1F2Dw0i4DWdDHj08VyIU25h50C/hBGOJJUmj+UaAP3ZRL
wCWnq9TxuOdGhauKz6CuHyIdJEAr5GDSxE/DvCnCz8LXd9eUPGHYZZL/34bZBqMm
YXPeUcynJiDKOAulhL4QZUk6PIP8F8qhTuQbdSy/EMEnG+31hOIHuP6gKzJccD9D
lyJ9H5JROs5BWBkJ7K+J+ofwp+MgTzTBnNywyc9f+/zlYmJZ488n3gHU7u/Td+OY
NzicLVot+5Cua1IA7cbQQMTkV88SC8IXJc7/uLQsfdaMGz16Av0tUW155TDzqhoD
EibWTEtFOEuyefbmJUIN/lYFpt/6n9vJaGIPQ6SnrasBglI7n+Az5t8SKkiLleFq
mOscL14HcDme0UcB2EW5Owt+3SJovIf4P3YeuBPplrDjtTzQoMVyqrS1pWazDuW8
hJgDlT2dypJVJfOLEwSKicbWGRYGG1Hn9DNxIAadLkrhm7Owl2tqkDbomiL4MLiD
UYJIjxhrbRHFI4D+rSyvvmCrujKDX0yZ2R1yTpz5TwFF0CHSkW91GlRKhhovehBs
UXpILb0gydmKuNYeaYETrNNEuslgid7mCq3su3XWD2wc4wkMgHM3iNWmxBnxkW+9
+tGz6RlmJFqzVLWse8S2VEhZidOpd2xnBAvYWsncY8i9X82ufgUlZmryNfIehcUP
E7VaN24F2DcveNs8pi3oKFUm78PiRP+wYNcfOQmqJp8CKinYsiLZOAyZ/y7IKqVN
z0rSUMmxvYO3LGla2bnPAcXqf8lekPFtine6SkBDU5Gk+YpMsE8r0VLkAYHS6sKb
Uk//z8nuafqtVUplmUzcs/eutvQkRJy4Q23GP5YNHqSKnnfSg6rsn4fnhvAf90z0
UAfG1K3+4AsN+VopaKmq2/2CxEWhpq8MUTOPbGN57ZbVXuBr2YY34C1nDIuUSChv
WhPSM2ZuraAvr+unikxxwGhtXyivBsb4PKbVdpZo2rOyZCmSyeDAbvZrbNzp1k5n
qiYWH1pypmMMtwIESrumYXd7TlRxQBAQjMH8cDKLib+spAv1tWJhpDkj/VSGavFD
kNjgarLxkoiGCb+K7iZaTElzTekp2gKmnpG8czE8J4xop17+e5X861TYO3IkLUS5
8Jd5G3xaini5/fF3F0FlTr7gasKX87DGBR6IuJ8C3W4ckXMwsVEQnHiXTNL2M+NB
LW4h7FKo0OYLOjQc2BqRywYRE6saXQsAUMl52i3YtpB8Ny+ODgN1DW4R5PLFTqQQ
Ms95zqAQOEuDOhL4WqpmSvkygZGzfoRj9LPYGr7tAecXqolGYULM6C4GLVs8AQYK
tbrmL+gv8Aiwa2hXNrmjBSVX5v7zJzgqJxtNoA/voMEYKATKQnjVSa4gwiPBn/Dx
+n0QTlW+xHMDnzMGlnlOsv0ui2p0Ktufg/C5oe9g48ClffLQCJy7sFgBSLIIMOKS
DjQ/X+5oqJpxdaHm9V7t/j93D04J+ofa8EfyBTICBZXdoOEKJUcBFmrFCIK2R2DQ
acgZbeCLjjrnDBW27LaTaEkSbaKR44yLnUhJ48cVILIx5vhbpbVx6K5v42NIxPeQ
rivxX0TTlDh+5+e0yRtnfS6XxneUyQ7Oe4vgldHeK4wucqpo23dHuW8mG38n+U7S
0kVK8VZ9lNgvOe7NIRmM2TseNswt5C1vk6tl7i9HIZuBWxcxfQNgc8sVCO8ohHy5
ass2IzqQP0qEPGALFoMbkPDSM7Z146hojoaEXSu9s7HPSZC0uCj46frsw7D5hLaJ
d/c+vZko1riMV00is4q+pgfQfjL8odQTd401dX/B3sM+ufaixMp+RHwGIatMwajq
pZUlpL60kuMiCQW2RjE7dBd+sZde5Qu8qV3x1qqWMYubxpAqWpd23k6rVW8Bioc6
1k74uW0VFQ1pPnJ2rbM/ilAcF3f2njzZZLLrB3N7pFRYd8jBLWydtLSf/a2qYsaN
YCGHUF8ya/ywDnGuFfb7uh5uYPQJ1kjCKiosvbfZ+t0rA0y95gm2jAL9huK/4y1A
hOj3/ig+5pptXwZxzsknMurEvtGJYKEJCbnakyTVtuPjkqnKIWBQPbnJMMMJEbT2
8bMZRaiMsqJGBoEd4Z/ip/3K0Wt6aB/y4fpWexQdAzUy4yNxF4c1oGqHszF8WCDB
vxw8Yesgvx5mtoGpQSto9BUm9ibdCQPij81EvJ7vx5qt8HC8pnwKYvO+KDbQwv0T
u3lFIcL9L7KdFf8vqB6ptTkWJ3ro9B6i54Hd5N3WweFvl0yumF4Eatn95EmMNwBK
VVlQ0mi9WkuICGPxxWTdu0d4AgzjHAy0dJ8ls2FVltda0R4O+7tzwxMZ0gm/9V9M
jTbcnUYUIfgbJMAxqTBmsMNTGtPNkkVnbvinhOwSLjQ7EfbzKt3V8HPN38g8QAhg
PO4eOmAKLTU6czeZ0zExVME1yUzElO2bqvSzJNLkQQBwXaGZdncptL1hgKKQ0XF9
XwcUyuMUuTihe9XVxgggZ/5UHj3f4Md7SZgeeCnTf43lFk5/eQ9IxGZNjFvr+4ml
ynHfJ8dD3ezf5qRa7kOA4Et4h/zCwEi8hX2886w8Vouo1+gQNlsM5n5RGBNcSwFH
E/EG8ni47NNKiEUkswkKw4CfsofoAUUpyFCWjmRW89p6ougDn1bDenPXvQI0Jyzf
OziZXbmZPKBUgGXKWzKZyZFbZrMC93Eo19sp1VhBaImEWvrkS50M8ID/N5rqXISw
nZhiCbxe4QLbN2Z2sGt+WJluEMtW2fWmnZy5YVBOWIeB0HiL/Wh/DIGSjwTbOCeT
4rmD9WLdQ9+pC4Fwzvf4jAYDJYkhmakcmbzVWdPV9/NkyqhCPcur6CWNQQdBtW2s
Ih9axnO4pkzVBn48OVVXsb+ftgQnX2LLPdZzaUrWQQhdMszETqIH6JlcvWlB+DQp
DtiYf/lPUqRjqt71Ik6K3huB7QIsCyQftUbuaKFiHJVIHzqPH4pLyS8Bldx1XTRA
9zikRuw++4jH/uow9a7Al++mhbdf+X3811W5pKdYKhXpjq6gH65M3iN9+D2mmvTC
DsDh4yCx9S6//6gOLVpDVx9/U3LGgqT8b7llvvLSHtgiu+9HZSzmXaz1b/VXvklE
odjXgcXaoKNENCUUpFbR2gnJxlnnY+/BtD6B+PcCXL5O6PcsboIs7Udo3Wh8Ywn2
OY/4lGB7lFhdeqtXjjI3NP5J4U91l/4QviupYzusDXlo9xjkYjLP9LymkpDrzb3r
POrHy4PaJqD6+4s+cwyy+ZFxGJepZHa7cpi+Oinok5YnBp+xa4Hb5DNCfDZEu3y5
xtIh3+Mq77U7KfgUEsnCvDL3AHGra0MOgp5Ger/kvdShyl8I/P9bRTujztPgRGxG
j8dofLvDYceKEqbOlFFve+pMGiIi0vy35HT10pp3ZypKjLZjeRAZsf+V8wsd4cJk
HUYJUEkBJ8lk2RT60NIu1FI+7AeY5P4FHpqyCS8c+otEZU3zz69N3rf9lF/jT9vd
qJXWKkIvl0TSzOsFnWd4FQNl13FB90ltzlaNYRdWC13zEEv0kWuhIYyi4zifddc+
n3wgS+AaaaMUdZd7spmvOTDMd+iJ9kkwnsFbnNWABCX83QLB6rrl7Ij00wauMXxg
CTTOPmmwUaRfyWdfSj0cb5GxLVCkJKKB2P7tGwIfjbscotiKKRXJs8X2RaQcIXtr
rWqJEqAZar4mF6BxVCzarLC6wSaKmkoU8d8SKuyrfhhcA/i2nLEmkdAiqIiAKa7n
H+Z3ezOz2DckrwEqORUK5fayUVd2FOoAVyxUUZcubuPtu83Lhar+h4hiAt5X3c5f
ZUiOmJEwSWlqPTe9GfaQtEmiKmHsQvt9ANNEnGisyoSqPhwNPwgDWTML+bSVEawh
jiuyTAlCF6+AvhV/ZrQjkiZcFSE3h7Y7hE5izBvhAa9qjEPBAFPUzgKdTvomFMo2
5+I/qIkJAlExyn+kXIta7677STZLLMLDOL7p4UqzE4y6AF8/LLXNla2vx9+PT9qH
EJWIEOxEIvOhYMeU6pqW8dkpmfwXnh4a/3QF08Tc2dOTtbm7rSF0ahfm6vtxn5za
JjxXJdFLINfVqBuvlEXmc3Hi2Oss4+VsYfGUnemH/ieH7d72L5+NKgU1+OaePpQA
BVk4u65oXnD8dnI7jrLCgxsabB8GmMwV5dJmCNw+ihMdBBeSwx7F/t9uWQ1tr3YU
0csqIPr2IUZpO24pSqTaPZKjfz4dGibey/7rGb7SYi/VBuo0htmQ563tFvXjiSEH
Que9GIjGttu3qCPwub5ioY3UKzYWKrfEWQKBH6ryyuzKgCb13e18L4fm9MODhxbN
xFZ4BAnkSrgtVeLoH0skbVDZeIp4TNiuZ0fztL+zipFCBcipLDQZDJ4G+gTwNew2
rKkoaGrjEFlcyTVFXynLOYqi4Py12rMh8kZ4Ztlu5KrAQFGbiAp9hjw8GVlxu+QW
e4oJqwjX5nFW5IJE0tSbQU2iOx4U1Tx5/nmfLuEaUb3mfq8o1+wcChfDZ+3vEBoB
rwcFm3gC+yQHMWf42v1BnuycW8tvqKaOb+NeTIZ7Z2k8apv9XvPvXv8w43hM3vwv
DbKa4s9BnNJ/w0SBSWbjjQkadix3u+xv4P1lBQJcqxMhPnX0FD6Uit+nqUDmMCQe
jgTErzDvu1gS+rBxc9DzGXt6HHYwGDNVqudzEOQQRes5IGcxWKujQGQQd2hkU92V
gC4bKYENX/kV1vNqkkMuE/D/7Jiqgj1LY18M3j2ynwiTqc1UUhNQYyfWaA/JlP9B
6wbxzmQSENU+pmESqK/sCATW8ONhF9aeCie/A99uZYA8oIzXtlr/IdJX/rJf1Ygc
xAHJyt2tNo7ex0PdhW9TtRLe+y2Pte2Jv1qwK2YN4u8DT/PYBnbYp/HBLFeZifqo
cFIp0fT3THyH95oM18eE1S7mzH+2mgxyP18obN6xZiqYachLPfzziDNW5IWPFxoH
qDTB8kYvchksP6ybhvIByG1ENPlnRIDNJMG+jyZ3dnt8xN4r7xj40sxJCr/jq0NJ
wLXt3mUlpx2k9mX+WbtOFhVrhSrrDNqK1frGh2a0/Sj5SL3ZjRaJEcRSukFwr5tu
3+MBXkPYFVXTvzUa+9AkkLx+t9Mb2o9/k+2Zea51jHRgkkgFUSnP8U4+J7+CJfWe
PBxkMXTxgw5uPdXw7qPdMs2ftB9vDg28j0sGYnrDWmOpLek8YUQdWzPrRTCY06cG
hnHoJwqkQFZj/KdacZ63Kf55yy9KCy+munOEYG9m6la4AghVNFll5StsZWwyH8QP
/585/Td3aTzLLCtE8cnzlXyG0771ibN93FGwec2y8+Q65+ISvRrgdtXgveaAEEES
b5huRa7KvQb+uM96BMH691tMpG/F3U4QatCB2QmPMw3gba+B9LLT58gLK6DTC1lc
vw6QlpgwrD7br2igrbNCqlOP6zDNIN1gyJsoyFhpHuWxpl2vwkSODmMSXYNJDBKF
XEle/2mdvrsQVcjjmKJKiqI3pf6FKjKb/ieFv9gVSsqmH2STedq1Kk35vmdrdmAG
Tf1roC25SdYWaUEpvtPvtstRhbQdfcirF9Pm5nk/u9bd1K0d5vxhco9QZRWCJXfb
G+lsRiGE+oSk2zLsl1ygO4Y3PY29MYoStEjv04oBJ8HKTSIOyL3djZQ1QSVHgaB3
LuHwlKAEPfvnvvXyD5txWm5/UJBVcVGEbpRR+cydlIqinZihKzfmdnOnt54OZjdV
Q7ADkndmVzPMjsvjFKtgllFCbREkKiptK6PZeLsd6Wc9xkf/W9Q8ejWnheFnpLzR
EZ5Nnp/1FH48svSgGXrYdWSlpjkvqyxQlX95/1A/1R6GDzleBRpmbzNsfG5Mtb/0
mi6Hd21X7pg5OU88CLCN57C9WF0lV53d1ATIv/TjQvuMG5oQGEQRdttkxll9TPsy
iRsDEjq0IHjec1DbBBYOtDXIPjXsMTLlCA41yd5Tr3YPmnYmJAIAS9GHmKMhnrpH
YP851Fg4MT/7EgC/HyKtclpDvdW60bUVnw6DJCB0c1XSJAW7t8Bl8HJO8FFJkU2f
V1lA4i9gBcw6EEmHUbcFP+VPeq3yCebaiGoGKKjwjYixnNAJXPMZ14vYxHGj/TKG
/2O91KZYNhRW9xpgnsHiOMRArej8BuZYtBKYdKcMFk7LSHjK99sn2YYS7wDloLw0
aB2vrKByxXD6YCnqRMzK1cUB+CASUKY+BzD/HzEFn/1VAJhnnDvXSU2Pi+4bBdDN
QLU/9p0Ghek+MeZ3Z157LYFDPaid4Dh5OXY/2jcYPxr8k8JxpUWY/Vo6/pl4kzkR
rLDIGXr56FOadHGIiBdkRAmsYH6E+RKBcZObJFSTlBlk+r5Hbe9o0RdJSLIvWZiK
OJoSkSvPGEkqM/7dmdCxGkzVzdRaQrH08mGJHIvy3A/MN7fRZY21c9eVcO8i+N9A
A+eYyNqbWGZbB0ip+ctGJDiHdh5b/19PwPc2VTtfJowRjNYk3DTpahrkBcmo463R
mwi1XENwvqrz6NdM+glMyVsM+/cRxucon1UhkfPJJFrv1hZgGvDAka6vqhIiYzeq
q1ohFkpAlYyF7ciEKqn2ERyN4lNNMBWz+TEED/2md65a9Ab7FiStYkbHm5qiGQqo
lTG4gT5xkDHc7A4FB2QxFOPJxLzOFXmJj/d1WItURc8yY822ZlCcAJfqcSirZEMA
f8dSWkieMEDYBeWqIGOhAaLaswKxku8XVl1tWIT0HeSaX8Hr+VzW+T7ieYTcVo44
AwW1aMC9gv/gAOlKA69b5WOmevP4YMly/uZ2+LLZsfRI3Bo7Pre5LiqmEXNSIaGK
p6DRGglsCka6+moRZkRUgXun0ph7BI9q41OXVAuVeBDNYbOWtYO/U4uFBgioIbgC
VbuJ80ghkTuLy+tDiWsElgS4C9Ap2jI7nQ/09wd7MntUf0j8m6B23gg5Daed+52O
PBxf+tOZpAzZ2+nyBOSEOmRTMI+r6vnKGqRdrF2KGkTvQtDHAKGzWktkFbuK7eBO
SR7a0iHYngYXN2tmDMalVTzmJ7hKT+6SIrZq29baw0nnRQZW+FYr+VjS1r0zGbWW
SKMfQI56Qj/LdsxtnLDS/KuHN/fF5CYrKlNcsZKUnFjilbXxNtegjzSNejivceHh
rRUga6BByWof1XFU7ybpN8cjB36STeJmdqufyKItK2+hE5qYhDGodhaoEyMokMVW
MWaHwa5LXhk+G1gQ72QdxNxJY/dQJFH+0/dKZcGhg5BOlScTTNUunxtCa6sDHxmx
3BIrOIyC9lSnLv8xfY030FDF7jzweioHtC+7H3fsd81PbDRlm0laXtZVYYfgMZE8
4tlQYnqGbo5BtnI8fJOLxToeypdcNZeHdAYDarUJAIzSdVKXBTfECkOsg3cHybGb
mLddAYZ5RZ55kF5p7rHBQjNStCi+RSEp0K3VY6URvmaLlZdKmEChzN6JGIaiQKfT
hAKiWVqz0oFcjRiSRPA9qe1FThjflrCNaaz2FGIyl1leRDOhZkX6vGC/pUWfspXa
GMcGrHQPcd3xcqFTuhj8cEGHr3rXQx18yeTSOLUDS4638lA+wtQmW+PPkfupEmMJ
WpJdlz5ky/zEQDi/LQAMjV83kfxDFCaF1xKb1leV7Tk2HiJj3gyuq72rc7F3eaKI
JGRp9leyz8sh12GLi4QoVnp474bTVAf7ArlXBAhfshAUmTG8XKM4/eWjvMOzt8E5
6YQAUKb0xgNI++RVcXQPXa5J0GLVECRvNnjXAB4jqE+b/ZdnxSZVvY6uVFqB5Oyy
zSNLJ7Yr2gHS0ZxLwdxIPLBMurc2iaJgaIx0u6ndjXHAXlb18oMl7f/vsMqnic+P
ga7wwrsOZrr6wjGgkZYieZ/AB2gmk3WiI/UhPfKxbM/Z+wHshQHDJ86nClX7xrtS
kOAwSfEwHLAAzFWjzw/yiNFssFQblNhFATt2nzEin1UxBsHOaDnyoWYPBMcUkZvT
6utHhc2q5/YbmX214mFTsb7zoyai51iPVsRUj8b0ppCSgzu9EHKMLk+olk8EY+Eb
cInJVPRQbqLDZGt+H/cJEJDsWrd9JGa0Z8Hiy8CN40nuiDZlDuKGw+rAv0AtNmx0
/HUHCyd668FbXSyAErbGGDTnfcPli44e2iB3Pm2Szwh1juxhl9qHhOPXkhhYw6iG
2KPYVNJwv6qZJrJF1ddB8MCmkVqqOjpk92ldniHj+l+UrxV7NIhDe30VDadU/pu2
2F3lUQaN2cDrqNRaNLTEZcVm1kw7FAtdpJ+rJK2LyD8pDWVvRHEaQntpFY+yvesc
UUReKgpzoANOGToRpCK5kSqDpZpMGfXVjQNd5E4PMcICAs1SbYiTL74QNXTPSrS8
f0j32zzzZv6+6NNBudzvTKHWxC84xHb8FJhBgtqYCGnGUCrmjeAvFnAe0ATBn79y
oeVyS9qZRe8OQto57UFYEdJ9CjOlG8oQffUB6ATIeHyEuIn4jp4LjlAtAB8eCWhE
DAgkeTUaAobNhW7rTm6x7ZF4+IftXKAqSjfco7FVYbjsLVfJ7rFOrNiTL8U0x2xO
dxBifr2ruWSNRs7V8APQ8+MCH8SOBAuFHW/zg5MBZOCo2zjH+IaSX2hDU0eiW0MZ
3joi4HjkagQAgHqBDan3V9gP6XFIhsly3VemiO1XBsBD/sXv3Fokj7i0ya+f4dP/
MownDqoiIK//Js8foJyysQxjv7e6ibEndI7yElK5gQEiXCv8txhxnj+X49qMD4DD
Vg4Doij9TfvrMWYUtmxh2BxMFkn6l7CNQkVoX9ZtAl8URpaGU7shQAqfDHvQpkK5
j8fr7e3RG/RlAv7DuPPxKkz17lxsDCSfHL9U0Rqhi291VdEHfg7u3lMDju9vHMJ0
RxxzL0f0kV2DeWaLWU6oMChkDuQW/o7t9B74zPVEOapDv1xmj5PtpfWc4x7OpUz0
mqkUawfQpwFERWuRbT/DRe3zIn78E4gJ2jtCfTPNXk0PcsjEdX/2OQyQLYhhLLyg
qduFztMf8PNpmEngQBBK6ACw08hyX2IzMuoBpbsRRtA8p+e6YYt2QQmTqcW5W1Uy
P4e9cXHPZXk1hudS1v/HDrBReOKrZxufTXfh4KMf8VI3FH0DDs6Dph9iVyTuU6SR
zlys4onHFFrr2SqPi/Cvr20ebHyvx52VvsU/jpneM2Wj1k+AwIvSFmXBDc61qPHy
e1kT9V6OZdgRRElrgWrJwY8uGMVduXZOceqpFGv6LS+I4N+arDWwDoIb8g8ItUuZ
Flw6tb78FIDhdjmI1/xq70NGy76OL9j68bFqN0vJVPiuUCuJOZVBQzJufhkV/kS1
+BuYArf5JoatYE7+sVvbxSQj5y+Wr4PbiGceLKScwLRq83FPSNgfz0a/VWvcSHst
KisvRhd/1oa8YWZFwW5KUgDc2qBALxN8D0ugi9nFy0UxuFEVcxlTBRRQmH+PhomW
J3i1wbfuRYxYJbqJe38V72Kh64gkdg0eetWS0jaIPrVjYkdn+OvvzDZlTTDiSDV7
Xm4NRbgziFoka+A9CEr6pUKTcCzG87nrE3q29cOG2RMK6eYNoHu72MpZ2BJzvRH+
qOjMablL1kZHNd27Uq+Jd6ckY7fHp/cXz927njJIjrxC5cmv5PbNEvpeC2E9g2wK
3qgYE641FVtNNtdF6men6ktLBv9PWFngQ6TpcTYi5m/Sd0ueuoEnXziR+MvXSZlE
NQsWinQrLVCwAr3Tevq7CiKixkRfn4xlqVn3Vregn7AXGflhCWFKjvhQPca5MbH5
4/zvPIbUrsD3Q8MQpEUAZM+Ee/KYRKKC++g/oRnXAuxyuAZisEENtCiB+6zA774C
OeBZ+XYUYB3bleLJeU5JdqzFqNFpaIPNOdyDc9yuiZXiBflXB3drymOE+UXcm+M1
fhs+HFf4edHx5zBbXr2Gj9MAF8/8zIAbvMkR3yMLhAO6bde/EbFEOIokXPGHBO59
S6GzmhRCP4eva9mYIV+GOzZXp1drD2u63XRu7XablgWHHQngbSp4anvP0/94OYV3
ZXx0pKHOcqYpzJ7jTP9rqn8gA0u+MLYspbWf+NQltcaHhVj0ntelYawOk3RNM1GG
9h/Wssy9aKv3SMxSz730blqIVaLHGlZNMyWdj4VzOqmUpELXhDvJYCUeE5AW3QpM
C9L9zp/jsdhCwvtSuwtSpdOnGGyulCq4NS3dQnqSBAXcighfJH7Tn7az6IQVEtFM
caq2ukovYTLNjY5jFRuY9+PmQPKdUkYwh//Enu7OGj24WLLS8eFGH+RRzcZK1xlO
U6LLqg9Jo/yLhvJNzZv2WQrNgW6KV9GJfOBEiHIg4Oj+pYlJhJZs3SmT19icc4kn
gSEtQ1aoFUh+JBcTV5Id2/kbxKifwN9KxPt8m3oq5lZWovswiK83vZOGPCRJ1e2t
JEp73Ch1tQ6P0Aq4p/1Hb02EvnlUiXSWtja9muNSJE26gjFUQZCVFHIyg8kWI7iU
DJBn8GQQLqfp+0YgeGlvRie6PrBNyYtexAnK5TUPDp/cmfoiARhGJMKGeZBzU1sz
yBOKMjOO37FzLp3xHSN3kWjm0HJ4l+nfO7hIp7/l9xrSr1Pnay7ad2/dA2gZFH0Y
6HFiavQEhXB7GkGd9GQVf6luRE2WtPYV3qpeZGIVsH2FAu779QdHA2b/oWaPL9Pe
YgE5vXfvCOIPT7hiZ3Z1Wpyxdx1pj8RQsHUT5bw9UtcBSmd2rfDsfUInRn1dLPV2
KzZfzkAOe39OTYJ6susWPhj/QNt/a4zhxw+HoVtZA1Q3jdWs0ltzRZoaoctSSyHn
cW8Y9d2iuwOtojxgILVLHTB1TbeWbHbuGOXvBMIp2bnMqFF9f6JiNMC44fRUCFv+
Is7BgWh5HKpiQSqGutVoSLExYqZYLMWNrgjPBrNDfvdMtY60RS2uSBrrgWyZHyDi
lEvkGOIe7JAYeQ+rhUJO/SGmACBHgQ2M9/ZWZFujWmU3341rlO+PxMa9eoItAn3E
QIm3eArF5mnQ6i04/yoCXyCPHAl8q7wmEpthab1lPeCiQzsewZtbhBTMboZeBGNO
pishy9yPcVEo2bOde6dpAQv70LxVpXWnM+/kch8mSrSwSj078PmrlSt/XqymWVQA
hLicoQ9SXiGX9GN20p0gJdLY+aFPYPfNg+ratio3sHjjRJCn5jUsnJTui4vaB/uf
ln+Vth3h9YWchJ/YUklUQyoFlybn943Wm5n8ofi5r1ri/QFdos4THZzVTdx/cOOm
Z5hoMu1QzMMKTSWC3aeGhgwJqhrZWZr+PNRB41l7lh6EkGCPs+2VYJD5lMCQeUJq
HtSv5CQzOOucfxchbWn0Bgk+ErXG0OTYFSHk8wolX5FJStWRp/lE7VqJILQPcnVq
kCTQMVgYU2BqQouZVZwBB+rewCvHBmg3635JBGZSVj9aWyCdFJxwdrPMK+gVdoo7
YFPIiRRPnrqEC5LzylHVxTRlCTnC7I2yODntCXIQLeVdkfVV6CQC3HX7AlZL2E31
U/rgx15QCk0FozXQTwfuIXdqvvfv6NpBAJU58mi0rPAmzM9uEUL3lJzYuBSbuhDM
ywBJkGEBTWiX/0T3tdjIa+Z/3lhybvCNKYIdEvtcMrofTie8C4fIsVL11qAPFE29
R447FtM81Qk/kn0EcaJFiXxmT6bDbaszeIs1bFtibrfgw8MlXxoPwNTvght4ri02
R25p+dGEUvwfaVWCDTYBq/9VwaNgm2T/uOomQ9run1FLNW25IA2LcwCTu6JfrhtU
SUz03GN2pD92ASB87wgUcqQ+bk2IhodE9esQIEVkcWJcIzrGFNqimDNaRk3gjwts
AJfW7N6QaNwsubUVOh1sozIiCGWfBeV1hbJnRZbw9qCpZGQb+8ObwQaxmdnW60vH
s4aGn45E0OeiwalscCMDJ0qNK1a/ijACONNF8g0C+r8h5yeQkYMZl7TIT89DsxGF
jTfNM5XW11FBBWZrCPFW12VcMQuBcVmqNZbOViuor+2u5Klg1LVcF/dM4LNjiDS2
izKG8n7L9ppWflzsCheMAmha0f4rBh5EdJkMOGFgqmJqbJLFBuU7TAQL12ZxhEOQ
JpgQMkgW9krRf4OtO54LdLOcTRJ2Xna7y68zB00fkKCjqkK03oYXcuhAbWymai93
P5TQ1vkDCj7U9P4G2ksCobSaxVLpYmS749YZFcrN/GuaaBqBV0eAYsMkz5ARVzyd
XroXe4TcKEbbmaQa16urtmS96+0krxvEHWbpdFfvKIQCkhH+uFOY9jr7gw21aLoT
bt6s9LdxYFe++VijaOu2I21/foExinee+AAdOu3+JWc6XuI0Wb08AhIkVGZIK2Ra
YitTgBOryhM5u7ej/ok7zfo2CEXg22nlP0QrRJfo/Ny5EuIOIqPQG2CfZHSEkhD2
JiguZIxDizpK+I9UT3RRigZ/uOiz3y5MbTSMnWPkWYTBlh0FkXLjMzfZLBLIVjmA
vVaHaSbDU23ZKz5PqwHZGaICaRe0jwQE7yY2wwsBW1ld824SiMUcO5zQG7qWgVy9
dkYRC2vKkubzf8oWK8PXT9nCdYwdO3E2s2RsIsGkvRreB7SgGVi3QZgNwrgOLIT+
VOVmaRlVID6ahnN0zHibCmrFRc2RM8grWJCRwioAMVuNc0vyK+8CjKlrt5vsCyzC
zb6Q7EzWjSPegS3lXEtIzmjkfi+HHOm/DSoyoUvbqv0UmNaf6AcuunJXP77dhNkE
if/zQM76UnZ0RIGk+d/u1fzb/by3XkUEcdoGpa97DDh8+WMZS3w56IqS3tnsPjpU
UXO+yoBkp/mW0ydHaeixRjkBz5DuO9yhoRX4p0wvW5JUVrPWBIjSPV6G+KzWGBJN
tFPZeDY6ySlORqD4P0r8q+uJnlvm0exlJ+deccupMw50GrD7mRpGwQZ1V5P4jrHa
Hl6IiYDnEBuabrGQkY6NUzqlx2IdS/nzyiPzfuH1Jyop8SJvzr2Z4WFNF0Qo0zGt
1wtJcLqlrBEnISsChSG0p/Jm8+sb4P2Oekur3XRUxfVdlNAd7zfSW30QV2rN598S
UWz5ENosmvBP0IMHzi+tp8XpdzudrwxWrUAQMNewvKffONY60tNB4pUqkH61tA+n
+Ui391w6WSqA7QPzoXF0wUPYJ0JUSoeXkd1lBJQG0lEiEghziUS7jy2kGyFlJW3/
6QXL4LX8P+sMXNui0m03vUgSkUdC76GW5F390N3yagUUtagzW75mqcUjvTXDxECw
eM52QY/0udiAHTBsoW76O/lF6Lkot3yarekuy24ZskP/9IBHKLjRKJdaRhG/5xJC
GLIuvdNaeVrDhhoXT4A5gKcd09UxFv/AhoXM+7Bdwc+MfxMhC8Cl0u8lS3+l1MER
Qnh2UEcIz4ZGYC42eZ6j9y1UtN39IVOD3+MXf8roLkOcNNtw7GFjcjoCzWfOiliF
UinKXK0rillsYjILiofHeVIUEe3GL7Mc6rUG2CjMx2kRFNqixptD1MdOmDbxZVD2
sdLf24Txy9FcV6BzAVxZRrzGPHIAi44i3AhOiiWGzcw0QO0tBZ4UN0USmzkm4cT9
1Ex96a4vxxfSEAipZKF13WHC3vzXgA5/YQ1g55DcM0aD31o67OcUrtr9hU5eJzhA
KL/Jq2BPD/JQj88Y2xbReElsFtBtKO0UO7z7S4gvrfWLFV/Dm0JzMlbW440FUXlu
R2DjoLnrp6d1GsgyOR7SCqoF/1LDhkx3xolIj2lKj2kc/nTQ6TOZbRPSRk0BEbLa
PPC1g9LIDEfrZ+UcEwQk30Bhn6SY6IoiMco2vHwycqP7VWoDPnlJXKUQRgoaMOte
G+Uosm2j9vwtAyDAcl7BeBkOwb2w0jXHnEgFHSSkLVqKDP9xNESBC/fEEfZkOTF1
/d8/rIkJxfDFYqfa47BrVapmJnrEObdVtrWpQHqHwic0FP7vYvAggAX5A8dCi89c
giqMkOSE8kwtUV8fS4x7cjGCnsqQ+tnf0LL6vJAUTpl1ZOnZDlRm7qgbJmi65C2g
/yWbcs2cCwwiyxrZ4yKMc4pZZwW53rJuia6BE1puQs6IM/jn5Kh7GNjA5kjGendn
AQd1qh7VBs0/67iDVi57RsGZjnujBilih2Mc6sPpJcuQIx+L3ci1jmduHJAbW/Wf
vODmuV/hS4FWVJBrGqb+WYsZvApjKVZ1X4xLPsgXBVK8iyucx6Y4bAx5e6nxLfyS
lDtEB7zeqP3gFOCDwwabx4F11ceK2h1Rbf4r1KS2gmIUdUD6XjpY0Nwmqi5nbRhc
Xc32ulyDd8XhEqzwAeEtXmg+KHkYFAsZpnwPguo58RqAPsRWIQcVf9iCbgcpX2lX
qiaDTcm3QwSlHNQ87OUmYV7d7xPc0/T0vyohHRTfgZubyL5ZKZozoW1AQLrEU8j0
zSQL08/UcxVBmfqO4oij6S1KjU0Wnu9/czoOaph5eTX0xb25OKCmqj6I7VMiddmG
2OSeG7XXSTLaYrJwUKX3NjcT7gHZCUUhM24TBbpsjowvy8NLkImZNNpTtswb7aGV
GEQ0WGV+waaVAKKcVDBR6UG/OP0QHCURYUt1ymXFjB+0kuntTJVGsAvUkmp1tHIh
IDZVIg8ZzAWgGQTW0Sqyg50lgSp28NhxejYz0K489P9RaKeWkzMwhuwLU44Dotl/
uixwim3L2xXizmlYJ07sO7uqQNGJgjF0DgD97R0R2xETWYeyGPYYL4l/G9tbZ7dD
+TwblFNfZgrFgpPJOrTFgrABQSgSXVDpqXmsgazK/2J7nao46ckhV2falvqrZoZ2
I+sBf1vU6WiyEFrqROspZHs+BVQFdfRlsMOTAaNGC/pWX4fb/ivWquTL/yVH7vAs
VAf13QuEnKDX09X9grVBm17BQwO1CKaNwjQILYPoVkw8OUv//D+ZlQ4C4FbRHe71
60rcZf18BDTnjjcUhy4K4G8NRWYma3uMi/ykDzIQhpB5tn5q+VSa7WCpiqC4bm//
IL65lHcyRNwKVUa9k3IfpzRWQjQ7v23fCKDmsiRF6UpJ/Lt6EaqmBTgi3RZ1wIo2
/jMxpooRMY23M++4FM7HXqnbLI/X8reexjtZjEXARwUCpY3ovXFoT6tqSzjj8Hdz
qOmaE2RnEd5jkmvIVbCN/2Wdf6ydBGrnILY31l7z+GbP8NkpcjgKQsR+x0g6jlHf
p5fgPoNvjdRvzfg6FE2p5h8VLSmRnLQKVvTCMMWt9u0WglRJMwesG7BtiWn3SSdu
IA/v4M4SIAtsZ/1oAfhIWx5gux/PXFW79cfgKEcssEv2FLsDLIbLcoovGMFpl6FD
imiYbU4mLqR0HYCZxSRQF9r1Gi3T2s2RxkmpCGn7DH5FFuQWm2fNJ3iISbdUcy0U
u2fNzJLbFjezDsTHSr0zSFasYEbq+sg092r8yANhVVjTYcl0PNKhSO2VlFRETe2W
jn7jyXbNhoCl4vGxDU64zIWidC8NtZ/LmScEVHBy8ZeOcoSVGwN17prJNSYR6zM3
c0NPAH7q2ElfSTwqYVseGgzb+8tsidbkSO0muKISYTPvbJwaKov+G1S9MbjXwAih
+JHRk/ISvxYAfytLFbLcFkIsfgQSw/TZ0LAAuCRWnv+FF7bIt0JAtmiB8b9ESx12
DJLcWSmefuCUt9Cmlbj8htJyEgpKFTQ/MtGKnBL8M/ig9kDthQ83pQEiKPBtKumO
SDBSlUsF59jInCpAVFCa5zPhNXanyH+KgIjKSTd6+wKUlH3YPmP56K//LImc4Hjc
vhxrWgffTfneV+/hVaAPiQ4GrDvrY2YZ9oB2P3+NYwVYJCujFMP16cC/xZEaiCPp
2gempHvw56IWxqH9dYrbUnA6zF01baximhwfz+uhcHeSpZZz5SY1Wu/6bmvEXARg
w/wA5Rn7UWsvWG+9MFpKFvrE5vq3h5Flc1U2V6CPN5GzdddKpDhxQ7CQdWsr/Rzu
Q4ROoctKkE4CeNILMvtQltYPRABNgBKPmRGZdr82GBokdrpv/qkYyjvrkRRP/l1z
E0jWB4NzvVx8zBCSpBv7/nOTjfEVGyn62tDujjHy1d7TKZIvFpCW1LEGdLTKInHX
93KMRtxt8f145zE/TYWqt85/rEI3FnamwJ3E/6KbzfHMjnFgzWjwqTZIjJzKvKSg
n0nMus1CPtC1XYLobqBHHGa75ZhSqlsB6x4d5D+IBmAioEVMhHSEY+nl+CdKZLAv
nNg7VzXjCTNQf8HllxjMeCwn0OfcCxGBDXfAqUNN6Yp4aDFEZhRYbFLuAvqvvThh
HoAHELRIKzij0b57+HAGPYALiZiUQmz6tonr3zaSWpFBNGKn4mxws3w4vkyETAIR
K/4Na4zDM2Ur1Ev7gYNikPbzrMGPTA+NYTs3tu3RFGQnGpo7eDmVoUcmiO6KvQjl
St6o2ktlN1+nxPSn59DNL6mUVoASUaCSlV3t/x2ZcdWx6PmxgIrS8qyzP7GtdI4U
yoWIH0jR2rnSo/PoZimy6MC3KYu7Q+w6VZycEjnF0UcrPtOZLDX1mADasmGT0t5D
Uxlmunrc4ZtGFtGdToV556WoxfYmo0Mpy9A35n0tuSwX9goz52iN3ADfr3nroVpX
3miHoVFvaQqTnG8oaYceRsuXqQV/qggWPMjLfaRAkSuZdmBQe0EpxBqZBCK4jri2
lC/My0I2AP8s86QNZ2E0hMGu4+uc/hKneUkvSubPCBpnjcuazCySggG+LrpOKqbp
uDT4h7630aVqYTivF8A439U+LEwTdqEJkUqOZa8FbyXZEzqLQLolM1SJtiPXZaN3
tP+Wo2306i4PpvBL5fktydC6NlYrq2x/t2PvKh58MuI7Vmt3YXlhnMEiidxwpB6r
TDZdCFJiERgbJ0w+vz7vSZRhG3zFbLI5nbr1xIr+N/AC1D88pAmr8MLoOJZgat9C
SUTDXmfNfyijjOzlKTWztW11pOULDg3sQLl1L4RFbb8JKONFelXCXRFS/64h27/i
QRkldSiGGM6DoyVG3Kj7QBAHrkV0w/xtKlfJNbY7TTjBwR77tPNcq7A+tLIK4k1Q
yRY9O9kffzwn5Q6ATWC58ZOXEyZbySqgaJcVDzNE479oXtKWF9bg9pY21Dc4uvxt
7TwNkFe9SyP/OTlktc2Rn82VsLex+LRjmsYvsG6BYePuFalTgIRDgwPa/b96BLeo
mGRUBnWjVgZpiJwA327cGigFBWCh9lQIN/ZcghcxtWEL0cLdTEWC+bFF0nunbynq
ru6Xr2CHFcCxmPcyCxDgGeWJr0PxQdf5u677EYeTX1IWbt0WfMIuX8D+Z80ZJ+55
mCKgu12/nWqWdgOHDX2Hg//X4+GsXqAyTnc6dm/dj/zRenoLO36anY0allQUtlaL
lf/skSQ7MamV4pOBnMkJ0mqXa6UgNdY6prW6vEScdGdr3Ct0SDFzdiQM2WrMIMWo
Z9330I3sB3WXv6jiRwjuh57iRlc60vokHu4vRDEBqYrYaztRssYb2KTLwq1WeGgw
ignKS1yvdW0yWj4xg65Pq3ycAdmbKcH5sbDcoAbifa7bXXf0lTnpJPTkNpqVkkbN
UApEY5ZCcN+dtEsRTzj0Hw45PecsQLfKPGeIKgtqt1TgL5RKediK8f39LuO2RVtC
1kMdKwYR9kFWqWm+nOe4Cwj3qDuQl0pDEsHFHCLpAM3AiGkmb9CCHISokkEmBDON
0fu48dcdiZzou63YxlvaZKrihMnnkvy0BDKcVB9gUo1vZMbGImWt+Dkk+ZsOfB/o
TjKcnFUsyrio8oGUU9w5VKiivHQkWwuJhI4fAPHN2SbY+QgKQsaRcgdBEUDzuyFg
7jilvuD5HeLQ9vDag2mAIvyXuzoV+altgL4xdH9eCrxcdMcOng+vKehxKR/DWoHA
weAaJexwq5XncTficRQm+o4jhCznmwOGzBl5HXLNBOH0zUsXyKkuTol4rRnwKUJu
VK9RSrdp7MmTlQjmF8a7zRPvNksZgiS/SWowd8K65icIW5Ro7ge4/MchmNn3P3vh
K/kS5eJ8yvAtxh0oAjf01cP0QbjSbPppEDkVpkQpmJC6n/7MDUxzkOvg40/QAzbK
vK6drHTOt0LAgw2cFBSd7epdnVftQRGQs+wPdy3l+uNXVlI4sPLfadn8Cb56tlyJ
HxS13DooXZLHhK9ICzeH6RaJpn9hiGWUn+XPk8/tY0tRWWGfThSlkNVDhH0NtVb+
+SBU0UUMhDuIt9qhqI419YA02FD/LlSkF2Shympnu/LkKqJBrElBd2AJ5YrnwsnQ
ccMqkUkDLonlzEHocDM58PjLM8/Lh1Hmtd1B2lwNp6Fz2ctwFnTII3ip9+fnTAuf
G1q11/VH2GQiSLh9S0Gt/H0yNbUhIglbH507pMepXfzYxgDNo8DADiGePhsYxlW7
ZRss4m5StOOswYWLCaCnZ8SShiFgC1k25h+FoO0EWu7szXSR4MdK8squomLWHAnC
AQHTd5zLwE0QEapptRMaNEzOmkr1BiG6YQkUDyqnnh9lFvGEJmACSU+/Dga93WGV
Lcf3gskixgNBdGQo6qjgFH6EwvFFvRJralP4p4GKOjNV5xVSeQh5pmBGLxfNIyMr
zx57MaOVh58c7IgY7XbTNUGHFikg5/U8moK7bevoVmqcfeT6annfZzXzW1WV8c37
zfKf/TmgvxJSlV/dAp/WbGUEEQNBi+AoHzoE/eQ95BUOdgEH2tU020PehZlxX6Ve
5XVXwisYIMp0i23p9WjKd9H4BmTPtHJwSPoXqojRTjRvYR5XsGnkss6QWGvR7sea
iUg35xUXv2QurfKOTBRGhTsaB+fVmyHCoA5Onc8y3WluEf99TByuKeukVz35IFGz
4Z+bFuL8jJ5rAqTXBMgeDHHEwUAjZv6e2xomRuLDw9X/Or9P6J123Oqn0h/UX1lQ
ogjToD0o3Cf/4RUSLj4BA0fIIUqVTJQtf6HDX5jKDVCR3cRQJdJPwN2XDxM3bJUK
mGbM+3s5AqygYYFZEgUaGRQD7WjMpse4dYsWlairQusJFRoPfQ5F42RN0GFNb0WX
dJtonKVRDnAS6u1GbujcPX87mk4viNJyW5u7HXYQIfoFYMIWwRRL6CZGBSJ7/I9U
nDAga26mH48sBcBffGA0tpwN7LX/WU/AdSEpLX5UXkVxEaJRTH+zTTC+ypto6fyu
REANICRENrjJQeLKPLNOnv5UnQQeiRLOeWMJY2yX0Oytmq+nvri498AtnCEMoxBp
MD9UQ6MnegMyYLmDmrbZAwrkp5eAPAzDM1L/U6zBRmoSUpT+f5ALwVU7ni6Mq/2F
KkY2/MRK38103O8WxX+fthQJK+oVtk8jrLy+V4saVPSrTf7D+MBVJJZAKf0XHOaY
MvEsNWGh5CkLuY8xz9Nyxw+NR5FKgjPhP8Iz4alZztLt9VXsjgtIJiJhRq6iO3Gp
4Zs75n8GPOvEE30MjpndFIYiY/fGR5KEQse4xtcIz4saoYbEnUAJaAMaIWe3akYM
xDoIMM+dRTBlIm+9023yhzjFna6pRNAygDdmZNOl0/J43vH6wXd1uXcoK8RX3306
El28fR7Lb7+4tl5kjS1RcDVOhcI4yOSELeUR4EGykEohTWgdc5jgdKpWE2pL6WoR
tLbggbj58ezDL4i4c4M16T+yZh5/fga/fKO+MRkkEZv9n3ZNHfnuQgHZtSZrm5Kh
cHfX08r6zU8HZupK7dCuC+/lNRRrfVpZpxOY7aGwalAkQffoWMN9esdMKafSjfre
O8hP6pnXyiSfvx+YNTxLo7o74ogCpafEhxhqAm1wJcZC84ULvhGlSYJL2CRQ5YNs
r11nhiLMfk+zcUY6vdawAua8EWkO5o9CzhzlwfXIziLdR3D6EqrO8ESusUD6mkSy
ZjymAhJzp+deN+seEaC5RJA8CvOgBzcUwsJI6N7Rt+WDNBMwx5PWlZ2P+wFEg+X9
8BDLGG05q80nnqCcgYwS6Na+dgcinA3qQZ8rswlH1XziyQkP/nkrgm7lgjcgsy/r
tgjAPpq1LaMkWhCLsRjR+cRxBdFR73Snyc5f/eW++2jL1Ddxbj6q2pbXBBbULOrS
0oPOvUzA7QmElR1VBFDL4fAAOzYIJ0xE4Z3cDG/CioFOSfNPknx3zyLyMwTKF3to
OcdBsBejIFhr4JWdX5TMa5H+CUOhdgB/Bigjm3txcjlHffn7/uD3gPTNaAV7rbUr
EEXRXZi99jsGMoWdVgESmYrGyAEmZ/LYFPVLVY+EfF9wC9m36Lgbma5pbCerXFYx
ShDK2E9UKRhzPYtwYKZ8s4tpkizcipT9ion1URbo+nKrkisw/v/fVDqmSFlcTjbe
c8ZW4exr4fQdxb1ADHRaVZIIBmB2eIyi5PBc1PVWwamkdeMpz2BDp/qPhZzCGZCI
o6WPl6i8CArqroeaJ+BmYcV8tzgvIrlzfqn019cAzGByZWNJKkkUzmZhMhuLbKHc
mxfnt/jNE3DIFIKHS0HO9ZahUjBtCdhC52q52urN+2wOpSmOSu+Mq5+58snEUgWb
FxKUxLDCFpB4roOSI3yazK/lt+FGBfc9N0pc9YDs5OZKeE1y2EfZJNqoiIZY/MiB
uBIOh+v4JSEQDvhzVxYe/TgsZlTPSRJC4174/x87UaTS36nmx6uSaqYYvEElDMK7
TH165lnhDN2uLXp4HAlhEP0a8IAP+ZnU0rup8lS1JVy5vhMlySXaepspI/iP17Jl
3XRgCg3G1YdI7AkH7L5fokvvpBANvnMrQHArliVf4uz9EdGfB0dpmr5to3ZzIeZp
BEAKX7/J9+yfEQ1st5FO59c7asgaosDJzlQtvUk2X49C/iKe1CAZNFG6gDYCLDku
v9Osl6+AlPxiUJDXrcTdCvj2+wYcsslTjPxKj48D7z6wEm8JQBXyZK1eVq/x3/Jt
DXNoyKAdbIqw2O/aEYSjzfJ9oT0CnFmsgFoWP73gaqvVgO3+Z8airIYC4H76l08X
OiO1RxPOUNlAfaOokJC3NM1IIataHXQ4OWuVeHpeR4WmZC8nwXbMqjrkqijr4CZ8
UI2qmBzC+Drd4FvUOQKQyQoHYbCTONAboJpe7d6wgp3uX2XJ0rmk1QW1ZNYEI1xA
RSLpAJ6WHyBKVGuLlvlfm5XFa58/nuSQXU8tib7U/D/dp1nq2eG0yvERda8vZ63D
jEQKOOvtqml+7krCPCMVED7A/yxN0p6tlqRAS8bFjl/ATyUUzxBJPjYeN4LKOah4
s6/M1HGnm29fDI3KbJoLHJB3QGLxITVoRHXWjHgjnEs7Jo50mno3VP7t4QG5Lbk+
270G1pLOLD/rH56WDKwb2UC+XZJC6/FUXB7CUEH/yltIlW8rEat1dYKQl+51OTn5
2nUd5X7KHKvS53dfa9MWau9DtjfBihS+IrT0Jokv4k+6KU00oLRyb5jQKmag7VkQ
GAckg6xYyMQJ/iSPTkNYPKosNDhLAABslsVERef7P4noH2pPium7FGdvfOTCKjPb
M1pVRHEzucNrNZo6UfGBO/7SOCi/eK68nKVC89T9dDBxK8rvAviAU4KvWQI8QYZg
EGNnzxOAGsZ2ky503sqxB+rVJhB8gDYkKq5Asn5DMMcQFycPVubo7KmHQHwXcGIw
76CUofY8Qte08vepcCfZ9icEUSbN5tlBhK+xoOH6fGpeZFb2Chmlz3twuTA6CPj7
X7uiBSo9MWdZCPkleorSwddXPmRbFbQ2XzLYBC6k0c7Sh6Zkspip7lqyaAgLCdUW
hMpnX9GNZ6g7vY6CcVStfySdgItAg1T7NQYKee1NpW+ASrX6MOEzkex29448GBTC
gR17f0pFPqCZ90vhtcyaZKyVXEG1fdnOox0U2MXXnSxMRoce++KdaTyhFaeBqOEA
w9hlt5FnNz/r4jv9omf/Kh+7nbmKPTLppOChWMun+83gDkVRiiQOzDA7l0ZY+Jb+
OD5ngQbmHAgpngIDFlct1eqSUO7g3hsG054FXe8H1E2T9w/LL/mmKw6AcGlnCg+a
ZqtX2drguOdVaitju6l+V71pP7D+eGur3kS0cbj7j58vjfDEJKV3Q4ViYUtKFRTp
Z+VpjOJwgO/PJRuP74N1aonXTTb/K+3bI8r2YUtj8Hdgh0XlHFCC5mEMk7UgUXS6
4aga4ytRML75r/dq9Jih9J2j+IKCSpq7qDAnIc4t/I/TIexKNnH0sKcwfywt2z7z
F2mNYw0X6XRxCF3T+y+IkBJ1+GwWTYm1TaHWc5dysMcL4GH8BBnVS01nSG9syitO
vS99tlWDc6sGhM+zMLYbMCnIBhAVbr8Tzj4BCJGjyXiA5CIwWnPxPOnFDueldCjY
/llQbnvNyWJcBONOhxIUMK7jEFw4/EfWS6sZxTFs8aIERzXoI/1Ddl21Eb5WWWlj
bunafgOjvHbc11WEqwgY220/Dyl1QhYIUdO9N0h95vutLpV0xso8l/T1DjpQdTtP
CbcBsajVgHX1GK375ga+S7EaK0yeaSzFys8kCU/88UrCoUwFXr3ppZrmG75rjIsD
74/ZPdbdhODfaB4cH/QMLIDvj3BfnLOu+IaSHejQKn12upo2jOQv9NoiQTjidll6
vcwlKBJlS+chMFX+R7rMNmlVLLj5I0ec+g7SrLHBWlFz5re7PX073UK0iH6k50qJ
wTpzXD7XWXJF1ScryM9N6vpShsD3I3mrfigPdMWvI2qzshpQGSJDfF1u1DHzEqcF
lFnYeMrTCvgRNrc+e4JgO17fOtOSGAZBN4BD0BDt37jxfvoLljZoyo6arNy7pAZZ
dSpxKejibYJoWRxsnXD1hS7HogCuF3EXixK8BDEwwYokoTkn/wd0iMijX/387sS9
pOcsA9dN1Hjz1tDrm9o0HcLkyDBp4afV8uMJp8AQNNpZMxIKcjWqMyi2YZ74Zkon
qEzZxYDE2q2D+52qKRlJynRwKtYelIrvUuu2HH/w4rYgIKeKzhZt/xBEMQLW19mX
2Moknez14gToUG01AG2lAciY4m5FnT/84wwgFfdkGsjLhmi5LWwZMKb5M9y91Vzx
q36WFQ84rFio1OY60TyUbr5cnVLXbqI0xZRaHZ9U24DXzmyevPXlg/jSlCnfZGxd
3PdHabTZGrniOL0bxZr8SMadD5CG4yL8KM82AqJqx8h+snl7B0ziXFYSirSRcQtR
g+2SqIC3oxmkwT+JrqaMaR8jS+UCpHotkswAuTUDhD26oDm4k+x6DyeaO33VGqJP
MpYzqJLZMQuKH23c00iqiT+b0/d9+3HR2gumWPr9XX4QT0SceYpO/QmoZQM3FKsg
eFKuHxxJr+ghGgVEt+nITt6iQYdE77hkkOcRbrJZbjtzRZbL8/0rnFelnjm5g/At
OJbXP9uyY/8qMacljH8TGTZ8TdRoAhrqav2rbTKKBj21RsSLxZnH+7d7yNT3K7AN
wsvg7WyhFeLGLwIaT6mcIs1RtstQqSL3B/gaSlU7wVs/geZAu6ANNaRAjlPXzzm/
Jh2bQrhFPGLhksdkHyP2PmPsLpmGrZY6gAgOfBay0AtCj+Slp87JoigTG7kOfPZt
loF2E+9kEkjuJG7y8cRX7349G00NnRUAUyC246iMiftlq6XEPEZda7e6J22tkt0g
bi9Z08Ig330viehTvPkphzXCVTsn1zni/7QpMYf35OKsc6V/3VEQVCbGQML7pjmH
hDkopmx3vrtdE7+qbfFHqslBT2h1SfZfhETYOa+1I9p6sml0A52KQlGuTz8whsDY
8xgGxVcV200W6yVy8HnCPj50XiWxSOQocUhfPVoflz4tPk3DwqWqao2a/SPqaYcW
X1pyB4ZnclHeo21FM6ClCGfRsn7GABS/d5P31jlLjA9BOknDRQxASYckWaWl+M7M
Vh/T1eopPDIzWaJp0tYSUEvhhmI0BgXNLXAp3F0CiRRZ15KMZDpSPMD4BLuCzhqT
g84+ScthcozEgfHP8EEa96svteX3zQBzLBlwgQjl+6/XGQHTCwsuzn108lA2VKWJ
ea+4gK5i2RjjgfSQbuei9z2sq23lQ/YGU+ykWj+UICP38SHM9SV6xVnOcaBY1bl1
eAHc4UxCe7tPTqEJfz0FA2wXx42cWlL2Zf7iU20s0CPl1K9tE7P7WqnGQpjzUfJ7
iDkIkT4vMGZfKq+pddWuxoBf1emRfT+1Z89imT8rVIrrqHBGf9mWJLhi3grouA88
HSyGsTwVUn5L9nolLc+W8zES+leSXURnRPUkQ3YbXUOBhwNpwXvVKc87IaIUEYUy
uJTUQS74vNJ/h6JpKSe4vfFWIWzqHGfTkfb5lx346fSRdoVdQ6nHb3ZMsQpr9viC
Dj6oQL9pNe9qD+g+BZ35sFmwTrXkNkByx7LhzT5CcNtz7IaHEVJm043CbeZxorSe
n14b7iKObN2+ns6Kd6hWSNlrm7i4Aj6Bbc67DKtMJ/sQtyA5pJdHycy1T4wIACDV
5AWkmoI8T7zQVMoOxQY1AbpX3JidSozbMDW1RLs1x/1Cu1Hng2SlTBNaqYfl1c4E
8xEdm9LwkQyoJDMUxdmtP89ENRWggOJaLbH2nIAAzCznn2H3+kgmmOJdJPiCf575
ZsS9DgiFxRBkPPuhk6sk7s7Tr3OhTnwo9Io8UYJaNc66HtVffgbawzXTGH8lkORm
cDiKx1JozNcLcXJS3YeI16aojT1fTfnPhy4OjtPbaaIBh+xGLYll4y+I0Kf7ul6e
5BaEfBeC+6SdctuAXm/zXgVvva6GbR/EsnuAUsy/qePnjjCTOS/ML9yeeivWX/Xu
G/gn/b2IJNnS5ucpC2jdNk8ngOZYTaGdH4j0sDHdca5iFtaSz67ItZxhlZzKCbzd
+mFmvaw8ELSQLPjabaib4jFANhQjoPCTreJ1g2EdvexutWPIcMycL4ojIHHAXwS/
z8j+JnBWcCDLnvIVZ9YEo0K09EYo/X1BIsr/El7TsmEzisnqamy9DREgrktwvfUy
vfh6wxSTPUpcsM0oJ09el/jn2F5RmvsOpdbm29l87p4csoW8vlRqNSEDSkXxS338
gf0yE2WTh/3V0FCOVu4+PBkeQekWDEpSoZcaj3lWruYqLvnTiW0tx323t9LinqSI
eillSn/IbJXG5yQhoun9YSEXI16w0jHVCdVFfLrtG/g/jURDwZkA5TCwBHvQnTdm
86MbX44bIT9lYg/y3yiFrGiFENfuJj0hpJ3OoRRo1qwJ4U/bIFIW3LxiTny3Lg2+
PBGW23VRs91EFCujFAm3omlKdPhczFBloFS2Rwv5BSSeGdtrlZ/P3xFekj4mnQYK
qYi0be7+K3No6Letuv9NlUzSxvgTNa38M6xDUm/j1KIVxk30tFJt45uFgmoakA2c
PcBwbUNJH0Kb5kyDa2PX0CdcwP09EuqokBAwc/fbQ29gPTHnVPo6t1WhtXN69cFb
7yMhcCjzR0dsVDrEbK6MuIj4oT+6LbjmsvOTS4h0BJNizwCIjyn5+ea0s+uPQxyU
ZXEnrybxei5PJiCuc0CDSyn3iuQnU3zn4PUtvBax0JmEz3Ev6mEBgfJ7ihtnPKIp
zogjL0PNb8NQfc9hz78c/hfAfQGev+JOkDBWWUMZIYB3b2g8HVj4efRzfYRNPzun
eapznqPW/f9vBIPxiv8qGLchnl4e7lywcjHhoF8/H9GGfHEtm1U8eYcF+0uJOeyz
dsXJdeokte1SKPr8LyUXPhr9Xu53sJFeoOhf7rLnjI4rNsLeYKVQloQSWx7g1cdD
xiXJyfIUxWzAkrBKPrQBd/Pxuuhb9+qMXESpHHDJPQCM4AerHFT2uUKf27T5Uk/i
zR22+Nvl2wU7Pt05l402tS36JEut6hEp7nZZX83XPOJqXxrHDiK5ZDuirDOX4gpE
HiGbZLc/9bar3OY4nPQWQbA22o3FSdRYG+AjD8y83DqnxRAYwoCAt2/4Cbybhkdd
7EgLR0m7OIkFRqGYcsL6ynwOQ5+6tuLgiDc29W+c8SuiTDsBjIsAyxqgktf9Dg8f
c9Z2rwgSjXg3+BYBHMWVYU+LpTgN0BSPGU5Nbng7Rk61SXK0o++he2QCRXqAGFTu
bd2uMicaYTquXJNJeid+VIBoma1+8vi5SXCMCfhfaJmzwwyKq3GTF2+GMLh2sF8K
yG7oUWelArmjBfM2r+ETd+aA2oTbljhppTtZEhg6YYgj1qBsnIkgcGg01L/l1Z90
515fg8/D9c2gjdCIrlkV+hQPY2d5AZRxJ5nCy6/P38RIrs6laMlnEqFd5gnnotDT
gQQ28ZI5jr+H3oW8BVFwHNisWnh/UtaRI+l9FQmtJkSJz17NmS7NaMQaevWGLJBd
SLghlTbVJNr2GC+R3f+0whNRMrBA1QXvctNnXz1muxaovwFftHmhcHi2vOSP9WeD
1lRH15EZ5TeinlpV0oMlp+hZBMKzdL4MAMC4oiZCu/hmw3HFBv3m8aiOJxnaOreH
a2gZW8j8fbmF1EuZB9r8rcuuNo1Dvt4yMNtYOBKuf/eE6urkPN340fmo0nhAj4fc
o+FqmahEhtTIbBKhSVXc3bAMY/9EByyRs7xDd2LZYoOssauURhfdelcZuvEd4Ewr
FNgoU7389A/s/6KPTNWq0ylJ4nn5l9h0HFRjn45URe1UGnmeBGC3tJ9PC/Bfvvgy
bBci5FN+XGRuhhVfh68U5r0zqjL5gKDl4q3UL1L0BR0A3oiarHdHMizSvljUPZCQ
rXDN2zyKkNKQdVrx+edn22kpBQxjfpqG4ydXZkl1agDXjVfKMq9OWxEfBu+ZhODG
K+GeXirZwIEuD4nY2gJuy8z/Yn/LoZNxO8OmJFmSl38rSGz3bKwpouV+1WqQBWwZ
petQuVD4YnE7RXlwZZY3KDEcdUg4Ot1DJG90Db6ZnehXvN4sKPKnq6o3hJU2DvuD
dRWXOyUSSJPtDm6sOOGtGhd6d7Ks8SN5k04HIlLqKiyW3at+hKaw00laHo4C2rhP
lC0tF4fRW6uTo2mlaqYSlDeJKhlOJVIf2ui/sYrEqB/q0V+AZAQavi3rGquiDYN5
YUHYuanZazulci+XNTwYLgtFAy6TLMEaZH0iKuYh11D8aRZHlB1whzQgWKLaSZTt
SPGdGm5scKUQG4RTr/1/PI2ZTU61mv6PDojzddPl/M/+3YMekDWIRuEr46v2dKFL
LYz2iWc/rZbhCfzfIb6uCNvrIIdqydDEZ5jU/XfGq4AxFHRBfLhAJ+9b+Qw7wZVM
enpmN6lBadinuAnrRBaOLnfKyArygODdbDQG/9Q6vCDln5cAMWPTTz3T8j1LRH5A
HKE6EvrySz+Slib5FpY+Vj+J9UJnW88HiYJ8AYkTnTXLDEM+e/nsK9+NDLbiBIpp
AHPHWV+9xNm7N3YTJKKxDn2be/JvqmGCX0rE2ywR2Jt9fwFtQOrbIG0vWBuAmEjS
fuUW0qlog6TWk9SGcnWtGlmhDryb60NSPDiiWwp2vqZAFX6rSAsShuSjjf6jDzP4
LT/w6D4nNrkM8ciukqE8LjIbCVqCyGa6ij69hiZXff01+AvRt5djuxiTBA00l8zz
ijDn69bEj/EUHzmLdNoRvjD1ChZujWNDXJxX5y+u2K1KaGGRSKPO5T/pk699FBoI
OMeJwpDqNuAxKAYqUv9nPYPylIxnuSfl0DXNwrAZjJ4yDbBGknUH7p3ioYWNerRx
V7afDlT5mFccv48L6fPAcQvpRU3y/9K0d6ro30n2bG6vRdcr0u+oIoAV2wB4i2+i
qMbgX8K/b35U5W4p/WI/5D6wAoNlgCDhCiSHWuD+N3mG2EqQfkA/0HkBIJt3eOPb
M6BEiKpPHLoTAXs2ShKOzHDfD1fxeqldmmhfk6TAhTh3QWZ1ZNrdBWcwmyuwCLs0
iG/RPODy86aR604+TPwGbhSncUur4M/51QwNpZ3r59aQ9zwnfGUScz5+SkEoQitx
+vv9L3Ix54xQneU9jT5J6e0D+EWpk2pTtMrnX456SwLykEvgvq7rFNVBg8kHnbW9
DP7s4Si3z7xm00AvjZYWVENKk+lq8tirXfsgoZd3mKu2tkHRiBuHKbdKLreqUShO
q/aCrmPUiszml3H/+OKElbns+pRxOOYxe4zpSFc0pGlJ2SFtmk7qF3oMPqeGerMc
Ekw3ODLrYZFz62DjvgXXScFv2QQxlGPihD6T7ryG3BwSfbeUWtMiol46xf0Gj3ib
YoBDSfzDPKaofITt6tPegKdZbFs3CfVJNQG0TV2fUY6Ufw0ZN4mpR4hQF5qdADDw
j+AjzUm23dHYTBxC3THYkVSYwuJ9n9En+z36zFDqCzpdK+IoxXAN2lNkt4+3N6Zu
fXOvzVMsaFMEvYSp2AxuvEj6H9MwRkI2D+lLu8ZRkMrbzphmfoVwGQJSjJYlmmxn
jRxx/lIP0c/Kfv2l9y8t3AbBTSlXYYcYl8hG6gWcVmZfffWw/sbcQ/KRkal+Gcpj
ExrnCuc1bgQoLDagxE9iDX0DQK4Fgcu7tn7GYgJNW/LfZlz3IIVUpw8BEioR0UeT
z7ijOVblAcAOYUu4OS0DFZZQVADLta32icFNIACtF/EbiZomAXUaIuKBYl4721GS
ZxAebeQGsX08iVWh9KUMet67WpFwNJrN/kLiKgwrIg/7CskbC27l0mEENqrWm7hx
9nV3nFI0QLbPiWnXZrgeT+cn4v8tN9OSrQPsvWABc4S5o1MTQNWz6gISPons36e0
fXKN+v5IHaQVYoo0M5VsLInkzWhmuY6ZEB2x0yx6yAuWLUPiqXk0Gd0WwXyBHwTR
mv6Xg7UnV7Jz5mFllrGFsCRKhUrFJPQhgJLxYK2jE6UaAOgoCfB+IunEbXHncm1D
OjkYV03zweqfCD6n2lCcc7/SCr0UveNzi0W2CTE1qoiGTIvDOVk3dyqoecOK174Q
CPv5XaS9wHjqRev9aGO+9JR0bjtnNE54pWdUbPSHdf8tndPtLQiQCXfs7IdMsGLk
2y/rFg6wEZ+uKtQDQUAMAS96Bnhzlv+ciQDQC6PxI25//UC/q+tZZXlVcewTlZ/0
ZAH1t5UCACC5RlGXMYPjGwL0CkfOI6dMzlpdmNVd89IDM+Oux+9746R2jU6jIV2v
HK0M7HVQ4L1GVy1IyoJ9NJ/f8Ewx6LJpgKEaz7SmiyPlA+5SaIjq6M33HGxxPZVU
z9YFAu2EYv4lggKte90IE3an46rfNZPEa+EGr/BZZYMMevvtPIkRsGuZUHa3tNLM
p+byjvXJdXEXml8Rs6+/rV+C6hZ78arJZxGaL6tb5jnCNTPLPP9aUYo02kMyyZrX
w8GIeNszsbeu8d0kCtLXjPjl1pxfPt8XAYYQ5Q1nJtuE5fXTXl73hJEqyeuurWEz
Y8qmxU4R1tDP+8unaaCWCrQztSbbZKOUmD54lcufD4nZ/mr+9Ol0hCKec4pllGo6
ifsLUWkCIq7Upvr/96zn3J+sW4h1tU3nB5Nz+DgQej3rFzXVtxuggvQ6xgha+4pQ
zQ+xh+YTVH1jvsQ7Hjo1ZfRR0RMUwcIpo/cJniE/iG2T7x8rZrQaCEgaFuVr/QxG
02/SONj21UHmOAdmRCOmyn5q663LY23xv4teQu7JMOeT6BJufbEfuHkRmGAzU/nR
1yvHxTc5bGl1NJu381NcPGlqFvhQFcpcMnRIO7NpUFI5BmZ59z7cHOI7cAKD/X1U
3/JChuENvkQ7OLF+lJxNdGbacef7/P9aEnenpg4AgIx84XApMAY7kZ7vxXKFkKmx
XF9BUDudnu/gjf+TMBVcRD9JzxUhICld44Eo+bNcjuqId67upoO8I3nXKu4kcWGI
RCZG4vYaow7s0WoJs8aEnQVKNAkdCwo+ZO1y0A0UzxlYkgh/P1GGoDL1s0qGL1v3
fN3UHnReur1Ep33oZtSqyEjgoUwzJ+e9Fn44leroBFcfuZRyKI97/TlmDInzRrOK
f3O3FgdZlBNJgvh6BHla3FpmH4MLaFY/eu4n6V4xgppzWX4yObp1HT3icZujZLZ6
vwTClm1a/3nMOF6aFl1n1Xt4JPWrFCL2KUQSNbkmNzKrSdj+sum2/ioaqc7kSEwm
ZZhGxC2gt2RfU63cDgajdvE+QZw2yqZZGj442ekcvTplvXso+d+iRpA4Cx+O0rWg
MLwzruwb71e7eqZCMwHeRx8Zdt4xnvxQvnw/7YD9wLMAr9QgFl7/aAGsfsp2Hlo9
LvnsgMW5YOf6GuIAX9OAWPk/pr7EXEjnwYUrKdoLC6RKlDxGeJCN5ylPFatGJ/jM
hVMkO/1fHzUg6W96OUojjlwTINChTfoYQ5CbownYt5p0TUzzYfLUEItxD/9AGjX8
XY+45UqQMcEeljIhA2m600OWDhMORr9+hN8K8aEIiHhQzLZVg9dkrxLWqi3G2gXr
zChfX/OhILbqrxI/nXJ7d/q4iEz1nf0GYn9//XwXeVWUOQfJy5K6IaVRlGotusYm
JUt2t13f+I7aFPUM+zc4F+JqDqlAuUgsM8V6pubBiSNZudKuS9OqKczAQ4bsi7QS
8ZB43mVTZGMqu5wc3Zdrt/ZcapR++ETiCnyNanqj7tDscZBBEaWWT9EHVzL6KRAH
KpIgNOtwWwNIpX1xmBfsGTrg656ZfyGg9mNsV/NsGb+hK6lHEwTcnPfnuVoaSpkC
O3UESTlHlI7qjnVvQJKt9icZheNUprnTejTSDLA4hzFFoTIeuJLCqt+n9HCjrL9x
FAFAz4Hper0i9D1Xck10CZ5E3kzGEviSpYXSfgKyE73TOtqiQt0G/ocARwFNc7xO
kXFA38Il7JWhwtyMEkF16P9esDiPehGRJksmbSOBYnOXng1WmdSeXS6TmaDybiZj
FU8kYEK0VmFTHpTlcUCmuyHtQi6trVv/Giqoo14mYUWRyAMFr3gIaMID71+ruR6R
zeT2AYn5ZkL/HyEpmddtrFmr7UyJYKEuToPtFqpnPdlUdKQjAcgvTnanA+me4t/g
+uaC0tqX5DzCVlsqya2xrRC8cjV1QaRMAskMUCgPn9IFI403VlbP0spHj5Rau2yZ
Ztn7bvsE2z534Ul7OdeyF571S5lqPqrNPueRn1JH8KoD2UDVCXVHatqiMNPSLKoo
Mj+Uif5QQAgH+cOUKYUbPTf5Hrfl46ZBv0j2cILhGCHo4RkmVQW8bmPBeA3Wg4K7
1Qt4PXKGpLaLTjfeHjkU5SwNdbRvmFvFyKCeJMExcIeDR95kL6OstGxVHj7nz78H
AdgOgvUXEV0aTvKKPuBAfhdRAiQ0Q9MUFmm0ihRhuHiXqKmVEo1xV0p5kqyWF78V
Hme93iOd3gajY4ovNCrwPrSNT+waNCgfmeweikGjx8pjD0BLyorfTLYCSVxWTQEZ
/XavTPdZOhuEMGIrqOM4BYnyoi62xcTxeAxKKbdDHEdbhP3ziM1uzYEzt1LbigrT
RA6F9kqNY3NpraLL8O4kYU09tE94Isa3KLzkjTzo1hbWG4yrJne3vw6uH49aCDld
gR9LFKCDecWHLIMmUqh5J+dbzHj9cT4/h58OXFaK24/ViANU2qCe743dwHYSFify
gEsywWQA2Jhp8ya2svDkizPzyjzImuHdY4th/shmLMAJ3T2X85qr5OUxLu9jti48
Xr4voXud6k+GCtC92r1o7HjgVA7xXQsywo+BgC7xHwReec47NdTXgJsluhOfLjOp
Hz2PSTU2VjHJMTkQEpCq1SMpGKJ3RzRKHXqQtOv0ChTwKd0DHOH4C0jpFFPL6P42
PtUkOq4eSvfq3s60bmHxs+SkWuf8y6/SVoCkWQBgTF7Gt24SVwpymBWVAgTVEazD
H+RW7mwbXVtzZGLjb6f5E1ZcBLb3IGi/IQUr91vth/OXYkClqVTkeHaOE27x/SxV
jERHDIZSZu+yaZrmtxdbGwU9Tm0bAfzN/vRD2p9njBj/CI5KD8NrPAwGbx9pQvvF
trkimLiyZMK01HRe79ZdShfSLRa2iuSqg3uUDA0ybPc66SEZEqvAZYb0cp+sE9/s
sweb5yZvy8615IpChSL/xzsYkyAVE9jJb8gRLjAf9BDGpT1hCBz5CQ3LcHz1EYwn
KI+xC7I4zgThH128I5r1fdEkWRKBPHtTSS3Li00yUIKS8JKhVvQOIOVypGCVi7FX
ZXj+MM4xVUOYrwkJ3TQ0ooAG4Pt6HRjviyJSG3tzs4XCCOxbWDv+62/2BND5ns9n
LtIaj70XRF2AnHvN7fP90Na79pEbBhRGvb1orTvI7y5JzULH/bVoCcTq4Uq6kW8z
duC6KYv7Pyyuro+7vi36DnxNU4Aoy2WuG44/9TCQb0MieUBWWv4Eqg36yPnGzRbp
Pd3mPrvn2Tk4HKW3K5+/UylRa82bgax4nUO7ERgw2Y5Tn31h1E0Si+IDpGqq+80g
lA+ZT0CYbk76w7tNMFCdj9E7E6+jxCaCljbj6SVYViWp/e55YHeC9Z/yYFnQZfOR
dPiUjDIxpJ/sb1LeZT5Xq3MHh/x2GqvlM8LqGn9hjVFogL4BZ5NtKkReDLtKRUxe
/rvVLWeMQT0vdDypJag5ubg9dVR1OnPLxbBpCWLNn+AWkfLeGujE/3chK7/5J0BI
Nb2GZzRSefaepcfRs3tgvzfmwQrnH3Ra9A2fVsjDOpvtQhjN4+//aFBiGlhAc4OV
DGsgeWA4ZzKn05m/IVBDd/aVygh4529zuow3B4h+dvAyQDJiibnmqAofgIr5UWEE
Ux+bU2+f2TX9Ss+DgSHEYx0v2zNSGUmIKrQl2LWJUW/NHImT4w7NbYjBnYOcRA8M
i0gATU8XE8lUCEZWMAUwr0IQ/H2pqI7jS9iJTQVPlJeb7awWH0Uxq7LuKxlKGNs7
6DLSNh6LhiOTPWP2fNWu6anrwueuYQyMIANourjJgWbSooVYVPm42TIEtBdr7cNK
yfzT0kd2Dr6PlvUuPfIirhKAcevsTxz9vTa9iTYN2o1gdjxAs9CSffQ9Ys68icju
HZwdwmRFrOdSXg+DpT7kNaPE+ibZQBHFWXRjdGBqrQFpzMRLThrllWGi0nAv4pIl
eEmcLSWYVwBKNdoYD1DJar1O2GrF3oRviRd/VJpLXtu+BWZ90Mws5rl5IdVdm9U3
D+o2duQfQpeqEok03flFXt8beBWMBabtSOnhzTvGclpcF+64RWni9V2xe8x3SVRB
lbe3erq6PsNZgaeTvfnbFrhB/idPjHgoaP9bnVzzXlztb9t+WrjnJTcmiboxAbBm
bghg4EP3/+Ktjd3S4+jb273wCJ/YRaT+Tj6ITA7F70NtDIxDWlkyTM0TAq5JBn4V
aqF2Mo4zSWSf/7Oxpg+k06cH4RNxLnIH0aN3loY/Xhh1WsGCaMVAcQN99ZLFC7X6
KSGWXo3ZyhOmkw3nvrBtdXFfxzmB9lZZaFKU8gOR9Fo7FKNCA2YfbQoNrl0VHc7n
KF8VyVVPjGnHt/An1qAa2+7TwLOter4m9tTfCZBGpsxwGm0/9Gky5KiwCCLkmCOq
b+8vTQiBmjLOGZK9PNGweVOPWqPqX1mws1ufNX0x8vHaaikExDXCOXmxRcuAz7Sl
Jb4oLHDNJqKWpqUnzzmQQqOyD0+Nl+ov309RSolvPUbpAJ/5u2QrP6kY4Kbi/yVB
vQtMU7kUUxY1+AWQmSkVDU3hnsLKV2jIrDhjNgQRxIT2SQiJIqVOfwyRNJmBs3yM
6S8nVk641cZHkoULP9AOt3+kQxq205sCGq3i8ULTljjvbOIgugtBq/CCoF/SMvg/
hNFKBwdaHZrtz146ixE3i4ITTLJ2gVq8xwSlE0gY2eoChlJauzxQe1DDuws2jUMR
gAZWGiR3OdLkSx47RRggmfhtMfT5VD9zaac0yMMVxmoyZPvMD5v2XQ3ClQDJd8bc
GDZ6lt0N++irlJCRPVTaQ3E+S/IgSoiuEdvfMO91584l+TxNct1ubS28FG6tC//u
5xhrOpbTBb/90e2kdkheQBhWEO6s27TUP861GujFTCKibhBT4AiBos1zbxLemZ0C
QCsoMAXLhOBJySKWAu4z82VLotF10R47RNJMQ25mqWSpfOH4DZYKbG4KmpB63YSe
HJkLjf47aboQcETUeX/Zm0Z9ay/c+TAiuYq9x6qJtAWwFz4v7lyqCRIlTxnzrXNW
krVkcxOFI3Sif8l01eHTJTo74T7Lsk/WmGIKt2BhNNSVvwLUx05i7C9d1zrcZT1B
GxOBtu7Gugp0buJbIA2Q48qWH6LlcN34FW0u+iYGgYNByVSOPzqpoyWi5Vbh/GC8
Rl8q6qXYmbRqeixavUevEhhx1wWGsZYJdLXOnHV0bRQ42g37xHBmN8ZcKAfXJjlh
gstmV4jOnc0O4ZgpXUSHSjjW0mO8qPQQUgnXdYJLn4eRYo6q6g3jxlm4eSmlrpLA
j45Rb3oFUCdQqAVCkV1pj7RvHhE8YWWF3btW8Cr5njb2VmrPDTMhZnGxdNJ0F9oS
TSN5AQgz+DCNVn1iSrTt2wziKb1SmHyZw09OnIkgA++zzmrKJB9Xh2KujqJcXl04
GxyD0O/dmTJpRcpIFIV6t1hUMeTQPJvU0rkPZ6erzBXyILSKYRk9Kf5rXnppdc6f
OQ/YFNt3AuSrL3GZCcI7LovBx6PPpw76RbdHRwZh1lQ4JvAEKyyAjOtuVjlto2Gz
rgEM9i5Q665FjUg5oWEQ28xveILGrWFGlQJIS/4QC4RQ2Tk1nO0W1vOlmSAWzZRl
xfENeUpTc5902qfk+ckFeXkyDPXpYMMgu9VxuG7BnBGkhddpzQOEc4QieSnvLnQR
fAruPYSbB7v6PMtZoomPDoNvTx0Otg++gqhe2y19oL3JhfyQjil93sT86x2f01s5
RrbUuIXN1q9mHxKM4sR3L0heovBip9eHCDYf8QHDHkq9hVuqG4lm1gYMfawH3qd+
Cj8QFVRX7bwYrkysuAdwHpkdWwNHPoV36T/+NAIVt+25ZYhW9/rQZle0oR+jT9uN
m0bHgj0S+OIzAvx/WYlCShHaYkcm8IJ4sJmIeRsNrbB7p5Kb3FBhY3fYzq6J8UzM
YOIYZFDkjbgVl4aYaws1xQm2s5Vb+KmUlOmNSOavAeDfAvRpmX0zIapuH1FC3NAh
2M2KmEaeP/0WqgwayE24LZKTKUS+KBxjgskGGWIC8coespbED21AAoNmw9gaENZq
dBf4l9boU3MxFTjSgt5Xonk/Wfty4ckU9qVGsG5Y/phepOkWYgA6YJE5hTmJKFus
hOJluCRNuNlV3Oq6r4K77UicBYtEbhgN4YqTMt6y4gFMDlC2SYyUaByJ/PS4O1gH
VEYYirL9HQFOjBhxnJg2wiflh3swKKu4NTBb7+lCEUOAS+QpBmDG13x/+kMTCt6b
iNw3P+x+RluZrC3n9Xs+SMGSzgrNUF0A+OcR6SXGy2yAkPocDsgO6YMShK1BK5AB
QPouh8CrtLUCG4WOTVbIbsS3kxhtxogxd+aSoTzk5QXjea3xmVqssv4dXSYoFTwR
Svm0shKeFG8anUREhR5Lz9ea8/FaAJNI3chY5j4aX83YqtXq3tD5Y2c5LndJRIcF
4SKDEeGx6CPbVMUKNKZ2ZfMtHIFkjY2ogb4fYcJ50fK+qKQOr/KTANTgmXOnZBjc
zahQgqE2KvidrLQYJNBCli/QkEfhivx9uJcFUerhgzeyRqwliDJtgW2GiNsB/tZs
m4/QEVDitkDb5K8kciwjDJf5JOMf2M6guZdhc8g8viHL5xdj+xdcDmiAc0nt9d9p
Ro9sgJWxxTKZU5c4qT5sJviG48hO22SdMWOLsxqP54zqGTbpIZeg33+HwM2kC4GQ
xl3G+MC2NyPB37kdTIo4j9IZhD/bg+TmYpr7pfGS7GKPv156cRQ7Ry6vdiCaEUHC
+I6xTzMTXWU/vbLHx3Jq6/3qtF9NoiChNpLWygM7/piYF0vYIB6mGZrpcPDfA0oT
BG7cWvopU0w/1JUywZTCxjKQwwcd7WdUXY72wrHb1HDoBhhMInOzchzqTRqA3SW1
6DCUJRUhRtlMsQYdWhTGfidriJUe4US8xSZ1Vid5MiCYQODrAX1q7cauiM7cTvgS
BvNflKU3foBapaWP36Yv5rq5fXT7bdptpPKTAONsWjRU0+9dKBkW+MoHir9Z2OBw
pbsDshcHVSqQ/HPlHt82I7AjHtuEgw/jeAFFtHqtH1xYywEPdZP+mxoN57oduqd3
hFPtTGArPQXmZP7mlZmoFXrIkPFNWgIDlsdY7OIRzi9L3M/j6yL17K/vpVP50Of+
HkOB6kYGtlA/PBqKea8TRfb05OwzZ5O5VVM58naZrQTEZAY361kTMH2ktKwh4uln
MpW93A8jXlFAGdNSE/jETwDJOQIqjBf8VdI2TSEre4PIrFnM+AyoXrAwLmneUnTF
Mtiy1Fj7wErXaWY8qEsbC6e0di8ID2K4B8Gy/h7Or2aM1Qpn5ukg4Xr2cix8T23K
/tEx/56UNIzvt4hF5lh4/SS0pVFw2u8thTUxZsENhoMOj+hp0Q/eTKqjQYJpeSbx
twXAFyuw4CTqf4wfV6/0Nmbb5jbCncdL6Mkf4GKq8L9i2sKTHtegf/0A16CHSCgf
UDQYdnslj2retIKXKXWazMDVq16RE6/OjyeC82RoDyOPTkGwJTiz6Pfu12zWCphz
trYTe/p1PTDHv6VsIEBDVlAx4IPHCbHB3ncgEpsoYPU3N8F+jBrdxyPCedoT5GQ8
ji3nvhZ3Ilr2Kov20T6aRPJE5DMiZrC2u2Wy0qGRLmJqipkMjmgdWpUqlGO+z82t
lwWIJpfkcO2lPR1lypx4D0mlYiALhoxK1z3NFtv9Sqncc9kuAoF/2clSMc5WScbl
yBC9TLZbgTmtAkCGH3AOCF+30BWc0SA1fhQlkA3Blb8Rukz36G8KojyNK/Gfad5V
JgS5Ei6e2Oa53KzrLLKHn0jPdFFz1uQqypQNLZtTTUGHuS6YDiXHjFdUI8dr72iW
aByZM8ryOg5oKuynwV663Rwjq0pn4A7fowXIxnVYoX4AAj90hnY6NFbhFjETiFjg
V0ipTvHMgCSBKP+XV7ImiD1whvrMNdZal9LKxLFDLBBIcFSkBoXBK9fUq5Sv7y8x
06g2JVECiHdCRfthRUZHwYLE4NYzHHa9A3XVl8VilVyXw6B+/ILbTuLEmGuwXWIC
wztw0P4r/Pl+zXzbbecG5/S1z+uKT6yX/SnR/4N8Xf0ktO2+3u82Y1KQykMu6b9w
pGsHSKzuKTSIhI4AC9o6rjDm4f2yDH4+Jxmia4Doa9NXA6n9Uy/fLsZpXFAy6o+W
hVwRJCvKZ1S5iIp27QeA0EbOWs27M8zt8zicmm+4KpHX3zki5ZZhkEXOb+tK6M0F
/3+38IUPgGFm1pdxBdCsX+u5lqqN4iUKMNkGLnVjXRC+EVHair36DMPmiXKP7oMB
8hBcRdOGmh2PtxkjcFO7vZW86lLlg9f7C7HeHeptPCAbA3V5dUPa4ye2OGeugCt6
4aa7pKPamHFeA3rz0aXQAwD0s1nuDHzAli7dvPGvjuRp2v1AU7P3MR7HUgwcaHMx
mRaee7sZEG4Zh9lij7Gb1WAwcNGU/SxIDCfwuN9pgDrb/CTV+73T5tC4s/WYrwXs
ZIjgcBujMnyIyLJTblGhXwS7QNTEjXQT//HL3/LjzhHIwFMU42F/k83Db+29Oz2q
mIu6j3tE5k690X2lQPnD3gSwGzRXhtuXoFx4YlDgOa8YUEKaELEsyLg/P1HprzCB
uZVcGbtwynCuzqvJqsDH7Klp1cqkwWCRnxrPa1XjkTO6xYIajnheqUBuh3+ryYMu
+wtYpT0ZgTxxHoneVBrjwcqVCg9ONkHGfTbUpdbcMh95nGKnQ9NZIadTanbdGN59
+N8lL7KkNvJdY+OwUDE3ANT/3wROIbaPhs/ZmTfC2laflXKANn+KBIEQMTaGOXJp
8vOJZJspiR3nZIMaPzN7c1T2HPGyNSN0OA1AqRh/rOelgl+bO5k3Qqc5zbfhkruf
7GZ/S/TWwWeEuvuLmobIWcUEFlnOtg/yt9xEQ7Ub6wBeGA07n0CdUX8+HmqdpOeJ
nPmczL1OzhpH7nukNNWFWUYSK9GH1bqkd7RxZC0zvxXBilQ6adnU/3rZZ3nmWG9w
bURvtzlB8RckLOuYrEX74PT1SWh1OQUko0szJpj1MrIF9FdtB8aZtIZUyriSkoxe
ckrxJtkWcL+IU9DXVKarguGnywGjrTw/smLFp6UfsFAisHoVVGb+fKeKHuqyh7w9
766ECxkHNalr+FdRcNq2/sq1C+AJnUqDGN49Izn/iua1NmTjbAZDSbHSb0BakIGi
cvF4A6oppOWLyf1YpHUrDh6a7leKougOcQTlqh0Y9QmBx858lLCuWo9x/vEO6p3B
Uogq0i7m2lwm58b2ae8ehs5wuk9EUlon+WCYDEy+Avc5GQmgCb2iK0r9nz8/RyVo
RaCqOm0KT0bhxm1oi8UH53loOc9iiHShkP4pjN4QrO16KeUpedJe4oIy3wKy605K
XoCw/zjEFUQyc6Qntfh/hVtGMx+vm2erse4RdbMnEN3xaWwzuGRlCIN1PF1g5NSB
IqK8Quj7vfU206aw0vKJ+iUDecZ+Yij6vy/PHlHrcxIH/U+lX9o9maK/q9fM2EDl
F7e5oRYGioi2K25tG6Jebwh2/4zUCzq83pvDxXEeca68+R2RxMkxekwhsKeYaaLM
n4XWdd1VaYSjaHjdWcNfUegqvXDk99EL0YP/ohTtX8JwzQK2m5Cu4kxc2OMrQ6cF
J7upGmVQBlUO955h/zDAfCaHlgoBwQjyDXszzYYAE3jJzXWYL9m+XIX8YlN26LrW
uLQ/fV8D8Zcd1X7dt3cX9GbxbgjuEOwcHnZXSQ5POdnpx/hUsoDpoaZ2MhLBlVl8
eQG8SjySFsZgYm249WwAbhNEzmlR750QaksAuHBbbeKjkexLHxjqw+I5o3MO63Sp
Nxro0LQ/oL7LEviEH5Bthm4U+sbKvB+z1jZNKlzVvXusnB5lKA0mqDff/nTLsrOe
4UrVxtjF18eWwkeGV2zDqGDjS7GlUpaXDKjODCTUYVyGnBK4wPejcraGrCbys2au
IgVpP2alNVMupJ8JkwQiFH6I6tWPU1UTkbKIOYIQ9qjRmjQjvv19xzK0/o+wCZWS
W4qbqW3PA+7xEHuDjj61Bf3YP3+75rr0/BrkK7+hrxTcoGvcttMLIpKYPikp0SyR
EXmjKvbe3I+IiAFqlnE352qfbXePgfszupWpAhFF9UDFb6muwgHJ48QzE/9hFIiF
Ydckroq0LGzoncpJBXIBtTP8TujCXymR+nfJZXve3zx7lBCIq8i2bQftrSirVvgY
jG0PPiOZ3k2xiM0lamRTgZaRt1eVkQ8KMyKXJjNFcGKKPNI3AXdTpgLu48PDZfKI
RFRRMr5AFui1GYKoCtbzRWwW2W8EbEAR3cOBdkF6ZuOChcHTYpiG3naxUTYKojOQ
iFUtTJT1A16ilFeNSYd6pFmRgyUz2adUSZQj4e/rngURQW3G7BOXDQDmcFuFQ7zN
gKU9P0mdsKkqLCMsFLcO0aID/b0vUqXXZC2Ee6bhuXBN5Ly11bekCJMALPN7iA5O
aE5Z+JFaG1wPAR2JLaTCCd9qGO43yWaVVTK60WzA2zO5J8G5YP3qacVzQq0xPiBK
Ca9HgIp3jmZXkOAz77uQItL48oKb4QTcVlaCRJ4CBCItnErVy12Jm5f0KGixoc0+
PrI2E0zc5TfY9eS68PUlr7Tbd1YAZJVqN8uG/WQo/1/tCUbPGOPZNHzMAKLGqqTr
jE/P2+heKjY7kVc+XYIz6E8UV7ZXgdR+haiopW6LHZs9bR++EKWsWmIRCyFEXg9g
sqKC2Rfi4G+VTc+Q6hoEeqdNpCTH/sWyPCOzjAK6Dz6KmY8+T6072twY/Nj/i/A4
Fl820X8M3goj+cKoHHjf7V3pPEg0wxHUtHDwnQOcM9oODHQkcaFzpujwU6gpjIuL
WQaEX2MPg38p9yygdZUp0R+Hduv91Z+Yv+ACXMG2PotJbLSU9oWW7qdeZMnBBANZ
GK+O4smjaVNC4URsI3cvVhTX1FFLsNvXqeUoWT9StKfgUoLpkL/nedMrXio4omug
JYlSCwj+07AFL7R2JfsAQjrfdpx0Y92r5PCMCnjMNgawUsC9AouQEghxm6ipxrnI
+fx4LDcdKWIBH6EVnaXQKsnq7CVINfH1FwddLjzmXf2qrjlhlMO6EBkm8UzKGX2T
NKWh2ZfOIeGFRy5IEetcDwkSimZGqX8RMSvsgFbr4vr5cX4ML7Af1HLsSAHM115y
wtOEZLFz/D0/HfFmYE6ZvJ+bje11kECyi6SLN4T8+VMFBJFvpEDd4RemteeGylMN
0pnSbhQ08t6C68ZTN1dwRasb2LjGi3L3An2413i1vN8o81CGYn6XVeW9Tl5/jzwE
hI/vDbOR/en5yfaCXdhvXazuWI10xBISDBpoEoyGsvCzrGKRNhtUmDqpGO8NvUT2
mWIif5fqRlgSFesENi0tDPVq6u5yGiMF8+M0El1V8THKmj/StFvfRa+KFScKneca
kunQnAhnP21QVjFGJrTTF02c66kTE7VXVuiVEMtspsV0QpuQUmcAVi1TKXrQGL+h
ZSkojil/S5PARWGM2rLb27LvxuW/RV/dtkxNO26lMxnkWftJKz1125MOjekM+2n0
1o+8HxX3hR9EEXH7iq2mN3DGSzh1Fs8jzWDLfvJn4KfK8UPaUnLdtPKgRdWtEunL
rxb0B5zkmTGeYGQCqZwnvdX68wytswvttEGt1XjzeiMXLwyeWvo3/yklaVKoMDc3
pw0toEAWXltk35RMNiy6b3WNn4sdTZFhjcwVYqHMb8peSuaAsVbY0d7EjRm3JPAT
kG+RNjEzPXbhJiy55i7QsxurtoM/+1sKouto/xMNIxvkeeB9rimwTHZKNqmh4+hd
0BNMKEXCfgO1akMxUtboGXLp/3mi99G8OV2EYPq5rsKadG8W+k9UUdxhP9j2DzQP
uj5XcxdYC2of045226IOZWf1SD/Kvp6JbUUvSriCXetHo5m4yor6vr+/JKOY4XDX
EquOcKdewgOUUBluL/sjRsgChLCrciMI7S3CgU1sOk0xic+2TB+v+usASLT2uin8
zQWO4vPy6ji11GmZj+r31H4w+hxpT9CVhzZO1toGAfpBrn2mwkS5XX2+L/URqNTx
WadnlmrEiFONVCSRcDgX6gZCf+R9bitIdsPrkVhtkMcv1AB/ozpc2e7ogmlXofOb
NQFEuQ5LGrb8F0QqiQ28vzER57R2Nx8fv4M+ivVezB1jYMoo494fbs5gHTvMBj6m
+zHzzw1ezBdmXCqk1DR1VJBO+zIdyckMKclaAZdzqcR6yT2Ic/jB4j3L6ZNvDsJn
pQhxMv0jZ0Axve1ZTEt8ZkM/7NMJoln+MAT0uJpYOUjxb5Ixe75XFlJbrfE+olbr
mim6uEhMNy0zSovlSonRcf7d9FQuRLlfb2BiIMghIzWbiBwHGxldfhZPDHJpK2RL
EyQXQ6h8uCfElCN/2hQW7Lm0zZCowqUMYveNFQWC/qRAM/ulfiO+ydEfWw0wUaDQ
qKxKeFE+A3+gkK8u7KLjtEt+uOih5LbNLYqSBPb0/UfxPXeiic92XlISjbjjvVBM
xvLV24mFqofwWsGlvIC85uEkMaKjG5MwAs7S0HXF2csljTVkyYPmeFtT+hk6ZOAr
SllwifJyDInriVFSa9tmmfD/A92pqocqgQ8L1Dpf+g7Hlc0Gx5OjaHTuAY6f4rox
Nqk28Iaa0FgBf5d+4CeO9hamRuPRycocQR/34x1TR2w0wkdoERWLTwXmWZjooHd9
zDrKUGe6O0w9lriqZxNTeOgz7g8G+2eYR9wL2WLJJAncsXbKtCicng71wDE2rdyB
DCHO7r8/+N1SzEKuIjvDkiax/0jnrubeSZ38Ig/PajkgX+xs5Hbnh4ou5CWjLQ/V
JbM3C86cEiPg/mxzmbecu9/okytbwD+PqiivGf4eMjEdLIQ7UFIA8bnhxdVHNzGW
hkz953MozRrwFJ72UQBRFst0GLH++cul3nMn6+KYh04fuFlVkksX1gD/NdJdhfKF
Es0FFOewybXzt5yLr6P+Ldoa+GqhCiXnuQ1VeroEnBYQOYp6Z0jLFaRbonExmuyz
DWn4twhoVwNuHdJ8M7HL4rADfpTXVLin5caOARi88VxjOvb/o9Sg7Gjlh1VoBUux
cyiXXgE3YCsvJ/gNTaqEB2r+3a98aCodCc4E0XMiCO9HVaytw7z/axhpvMEAq7IP
zFWQFrJn+LSqPHIkGIoYgIPKdcXR1x8f4X+Nfg6WbwAw55QblJqp9tTe4Wp7yPC5
DGC3MTUbIfsGzxmoKQHoVZ+ES3yqxCPhHDIv74SIm9SjdwmRGjLCR/lxD9j6xmWo
eScDg5/JjUI/3BBj1fne8zvx+D3iuq1OhjXJvazu5cqzWfvJqjns5eNVh0GzSXIB
nkwqQ0LSoE0+hK0ByldeP0OMAxGjn0SfqBbn2KBIziR9mfQz/brpKHcOfDchZ49S
ag2k4Db4d30pA3RrX0NLng1oY5+awVrKNSf+z8at0utcj8JQkQ2Zcjgx/42pYaLg
izoPNMywjP6rlH1uXCsttwWMfIaX6CeyZLC5cnBeh7Z92+DYpBSx7XX+J2sojYU6
7X/htwts83yGpTPNAU16g+R2HLkXUuN1U6CeZUIhfwS3pgr3u4HR64hj88834Zqh
whItKI30GJgZXgud1n6PzM0mIQUQOHzAUt/t78tW4d78YshcA4M+KUecza25RlNC
dKlOm6hNQO7FFWGOKadxVnqYaKeTTttDSeM/jPUytFVLgObjm6iV7uTcoX4Op+CA
TJmQQAMJuvTFuv+34rjl4/AXvBydxcr5nnQOzvJOWWNtLSkm4evosEs4QOCj24cF
CNqJ3JwK1DvJenRVxHO2smX6xrhL7Ngo5O9WY75VMfdfFeCaXoHgHxWDa3rNutTy
wx+SqxfF/Ew1q1Km9h96y79sMeTzBlBKVrYkVNNQXWiKGV3GnQpqhR8fybJ/zc/L
JQHUe7thp3BOtDPZX6GWGZRFqW9NDzv3jn3/j5cs+iQ6pNW+xoXNwNmnEH3VFlUf
tn9qT1rCjH9vmAQUDsxaKXNWTpBUIxhaMecJGqA6QFaP6TSxMMzoW1ZxI2U23oFE
IaNOH9DbqZ7Rlo799Zk/hS3Pys7bD8lqnTToOZVT/wK8bLK0C9XFe+Q8S+lS5jAg
NRP5IHHDis2SihHnOtNX4jLZzns97TWU6Sd6e0zz+bYVJ1v6BlIBf75hjC4DY5nR
R+8YkP0swUGoPYklOsScBni1gWSwmd2UmWwQT1cocYlyCc0v3JGrL9MNn2ij4oNJ
V9pvy44+wmL4AeXIw+o0ANJ6j4bkTjnwBuGPdXdD9HTECJAKcb7jGlqccMsrs6D6
5fuFgeLKrAaPvkjEIJSObJh/cUC4AmGhjjQVvFvlppLasctLV5e+dIdy4LFiafDv
6XyhDTWYXE1uls3Sicx1R5MWbcDwRTzBZzP7fzxf9Hl6j6jDNl2d6cKtyLjXeSbF
tTXHGBZYiKWO5Vfj+KpNOKWunGxsarZzgeRdyIIKvUQ/Jed3mUCERGl+0sHSajCt
atNKQY8TodchlMIO1IF1OwA5FGjkiiPBXOGhPUdmP4YPTdrIIcDSBHetb06vFEr3
+7Ap1x1Oemr21Z6l7NXiXweAJnaqLTDkFftBYuocYhYYn/zYVDqrqPqWYeXIWCkw
dXz6muZ/zl8f7YxGLz5I9JXXhbRGNORKeuxbUwDb7LahdOEE8qS16TmPtrFtM+5c
84lMW2w/eVMjWefOAAnT+CsXswbvNBGeoCWpvDVFWE62I6UnLlUVpDOSuK54k3xd
mvPyGISchLxvxjrUzKDOtAbMD4to/AvODpKN1S9tWedNxRS+t7+Mg8Lw7OsNlCL6
8fnuvD/nS+fLYskn/qV9CDVZA0uWy6y/0QIX+Ow8HGUmIVBo6jJLtWbYFq8/ASHS
8jqZloDpH9AoVkcAEK/97GMriyyqoRRYhKEyU0I9DAT84hgwMUCtvIoPBqUqonIS
28jdRCdbMkjNLvCtMet+ldX4ntfqKFNCHgGdPipyXLnAZYIhVYqznqx83ipHpLqI
LVjg440wHO1yoBx0IG2j6fx/e12HjL3Ya2JiFPUVN+GA3V6dP3HeKpJ5Q8JTIZeC
7wRULUfDTKviNHH0RXO4Da3DPvEaVFOlLZ1GUi2hB/u01O57pXP9EnM/gddJUWLE
JFIDtgAyz2SsNpH8765iMoQ1B8vv09FmFGafuKYtVn6AHwgXR/+FOKtZn0B111+1
5fPef8uX0GDyzJKzJXHAIiN1gc/Qgu6jiuTeiaCuSZvxD5KTVTIpyn8nbvu+aEt/
6TLyRZZ8N/oi7H5m5bhbVOH+xHFU33GzL/nnVa/SD1YywIn4JunyauEXl/AsUBwk
29lFZWJdEcJYqXbsawVI+4iZxJVkodVCF+a9d2m1B3rCljJyj5bfFRMhqAanw271
0O5kISwO3+DoXbveEBcpxLGtnpaZIIL3s23rLFCF2o//InGntJRB8IdnWL5fwA3Z
I/9fL+xAo9/+iSpxtW5fqzpA6jo7og5kZO7bn9qOdVwv7q+naXqccK58+LrlC1If
4ncN+yLLt78UnkPIijqPcUNRujSFRolDoec4K5xv+YVJsgCzo1FLkFlQEDpqtfhC
5Lqd2LQIVv1I1LeNKpXbMR5uh1IZTZwwICuytJkHc4BQP1JeHNuEotVKEY2CfaPd
xD3sUtkaYZaVClSFhQOLZJcHzAWY1qEGmlutouWqxKYEujsFaPuOvGNbxkxahksu
DE1ubYOn+Xa4XSx27ZNYtgt8tbL17YWT4zwfehblU2YbSBQKMVR6tQ+HwvyF7HXk
bvEDQE5KeS0fg8jXR7JRI6EiAOpyLbakKYwBkjbQQiJ0qivnIUhDqGiBNBHgbuHi
wjlXfDGq9cKscIIZvFfSPFrigsRHkdTTvEZQ3f63lfSlKg50zywlSlJqagGBBht6
S0evgjYDy53Qgz3KsxomxV21743pC4DfMQunr2ZTHK+plhWVUaEo6PZlKkbxv61k
zzUhG5VEtT8pWDIuHcGrAghSOOmrFMFeUnxN1SG8INIK4fouverQEB/ZtS+7R10E
2bzjD4fK3526rn/Kb6QpqX34qzXoXIIsMUg+FX2zyA+sXQz9qKqf5mVHS16BAB/q
5uS5F9VsDNl5Z9snRDOr+bv9xkTHxswOYi1ToMYAMStNnb4XPvjqVsBRTKAZ2SXc
blePru9ScPBtJdS8Tq7FUXO90Oi1ZyhfZoz4RV7nR2apaPmgO0lkuUvQV0SVchg9
bmBau0XiqQpuaKI5UPaXG2c8tYNUDbCRp8+olRJ6CunE26PfMHlIS/AihHqHsfdG
YYYLQxNW99zxWQEDDyjKMLGeWHmrNz2tkqwwszw3Lq2lOBPhxdxFo3XgfFlxmOOX
2mVEXOqoxD5+z5BjdQsXplrss6wg+tjBJXU21/cT2K+ZmQxUR5JNBKSg5AOX+j8Q
t2Bnq0+54Wg5qb+d6RutrsnJuROLCAFprGOM0GC64JfQ5LbosDSh94JPloI/REHS
sYx1N3fhJ8PJtlaXBGLXeZpYYCLq3pKj1IOV9n8lvT9TTcC0tEpe1SKx7gTFiH6f
4zwguAv2O303x4jOhMRkFF6TxPQnHj4XJmI8p/hVRibIxJsuSxxJY4ucWkcn2O6W
n4JfBeDSBpXimJW+1LHN+Ycl9qiF3D/sNDLpbaG8a3x3dyCbdijVifsYxRAQk+PL
xeZ7YsSuVE+O553bZwANRu4KwRn5uuTv2DWIwqJi1T7R1KJOe3/h/AXF4EOClXlc
MyAX5bPaiccBSxtLkFsPrNIrw8bGhXA5qlO3iCR8JT5GYC7IftL6q0uYzb4XZLkj
5jlCbIs8jpn8kVdu2M3z9RuAof0yp4IAdDwjQoMRHqi3ORD7NDewX7jq8tR05QrR
ObuVAmqa5sCxv2Z5mDSCKxbOsi6ebRJbAs3Vb+HwA7uCQiNKolPn6vkQI464V/jf
zMLcRbg92n5vtB6A87tT8Z78NNHzz6StRsihZ3CrEa3a5KzMq5uvqeqxqIRxYEj1
ngnd+zoXrpCGNEKWDoBsUpQs+diC5PECFG81ED7ftH2iFHe97B71TFhrJEnmZ5Pw
cqRJQQMHkzrXo5vBf59SvZLnlmLAWIYFPmAdfOWRh6FOxd4ltBHGSpmUqNIVKRLF
XPbeCUKEjzZLdQbHYe9XRm80iPyARV5KUFSrdQwQp2HrCQvCVSHUGOTBACa3Vtgl
eNwO8xsGpCn9UMQvKLIgKCYnjELjpMFxBNX9tfZb1+hIkBWXq4koBnjm1/XyPABa
bRCdwW0EGq6i4U6J4Oz9nAjxOGSKars/1M4DFpNAfBd06tRUbqYaEojqDw/wK2dB
Rg0HGLsP3QOTR4dkTG3syatKh38gAazpI4m0Ujb5l6CckzHPSpyK48YxihqXjIXe
CcIS7cXKvkewsqwHRs2q6Vet9BhqJ2+EXuAf19fRLrrfh+U5AjdkxccGQdiP0wuy
C5laiwTV9+7CbGCkSq6Yx7rh+0yGJQ9p5TQaig5H0900Ugka6vPgtiMxDxjD75OX
nX+fD/NZElRP16prUYdgLeu8Q57X4KTkIMrDHbuFPNkEbvlnj6I1nKfeSEYNuWqO
rvt0ALIHeoN+AKGvGVb+JjWYRRq2iu6agwIee5byFD2B1qzJmLXqLDwvsc2prglI
3ElPgjMOWqAsi4S++2fiPjlkYi+OVZPDIbyRu5B30KpDY2IJGwDrGgLqsJ8BmauC
hudWwJl+FoWIAnTlD3E9FgWjTZU+kLrD0ndKCGyM+ML8Gwuh5t556llEuf6hZC1+
EPYqjyMnGbXI20pJpn8PzSC8+kTUoKrvYc5M7zk6SZP25TUFwN57P1tAqcRZXrYz
4D8JN7cqpVXYvND+MT6mTs65m0/vI3NYyuhy4Bw6I5IdumuBwYpi/rnJyETLY05r
PJUyNPac1vTJme5QwF3IbxSeZ+JZeUwAEc4RuKLdasIiL/MqMS3Na3COtYsuXKCr
ktQJtSzL80Q0DsvWl6tz68mspF+/rGgTuq/uL4cpIBNcPc1XB27Xfv++K471zw2T
qod1PPbXr+UHJ+/2TgLpO6D41GYtG2kUaGvuIDqtDUPEpQAOlwpHUDJU0vYtcGtE
sQZy+W1jLLt1uXPW6behmkRyz+0HouO2hBNY1PGs9KDw4mHS0HOD5avVT1aei2K+
x38GnF4K/9k20hjNcTgFaNbYYFkY6ZwbpQ+l2kmfRXBR8zcIyTBRA0yUGBXPX9Gb
gd/HuYNEowte9tMrcscAExnRFqlmDJcbkGfhTxo/xsdBtOvwY2cHGkAyV016spR4
uoF3jAYKT0hEm+6fhcRYkXozgvsRZ70BnBBX+w5RoKJ6yyp9mp5lMMyNb3yKc8gy
ZFGoTAav4g5j8rX0MLUBkgf2hXuoAJQ8/xfM4/X1boCXXOtdmzUPY9YI5jLY2Rhg
Ylsitll2KheHlFsqXkO9rima5N1hrg/Yc3lmofLuWSf/KcUZzp5pS3SnsAkGW3z+
NiCfL14uwRklFhV03KdAG0p7iwK/l315Ar5cI5vcbXHhzwk8YXVRVba9a3K5cz1Q
gCe7vwfL+yzAAi/g/b5tx/Cdiq+eNjI4VZZMjxhl5fN+cWV4JXZxvxVqY5TQE/ed
N6L1ReT2LJwvxmQSCbgT3Wb8dk2XOzbwZlJ5Nlp54P4rVt+Eoy9+8Q8tQb5OKj3S
hh1NJodekfr9+DRsZUOkCUzmuqI5KE3C5++I5sr41pIHMb/qUlR7/+24KT040e/t
YxBDXHTFdfC8Qk1wHklMU7aAimITcRbBIwetXwE6JxTY26hyu6dHC4Pcid2mOy/l
XBYelBnwMLRFzXJuI7zSTuMdi3HxFBeCdLgkQl5FUVMQf6yr8fGME07lj0ewDnHf
H4czXKFuHWap256r8DcvXTMOIHsI5gYwgJ6dEgtQMis8Gtcn72AZS4hYSARUrR0I
Pd+tnhBA4xQ7ycpB90sDpcWCevNclPV79YTOJCHIQCXVqt/atbk39Kz5RDmKM9XX
TpXd7aj0n2edBKzIH/LN/mDyJ5kVH1j0V6I6sCKlpoDP4yXrBrl7ftHD8FP/ZQd6
FUKzL91bitcaTslDgmKKry1dMsGVMR9cloDCf0ruRwp81Z0G94/5afMinOqCZCuz
NFRAVUHM0h2gP/vaLG8Nz8V5fNq+yKIZsQlqVz9VwrceZXct1zDv62Z/lAbjFfe2
iofYGG2po0MFT8Cb1cBmQjDNdS4X3Y4cHucbp6SDfaeeSjLIIxi9VUf29o2W3GTu
cx/iLYjsPLw59RD+snugld+KI04PXm8DwRz6bAkucgP+sXZQcXfWpAlFnPI02Ld0
juOEYrN6g2rXTs5JQX1qJkcRCVG4nwasqCWvLz8fN9EH8HqWOjxbY5FsO9sWx1WG
Q1LWWAgxLYZUQutkeoHedYBJ79lFExtFrzlNrv+B3YBHPJwTRSOVUCG5FLo53pOg
yL8MJdlpArShenNcZ/TH3r9E02X252y/4Hi9Bh5HGTnt6k1ob1ixHnqTU/N3qmEw
l7o5fzVK45hh03bLLv2CoKHiZT09kf7sJS73i0ID5EQWIwkwWcjfV+O1PP90kEPD
5BEvTYqYlJZ7giBnCrt1IaxwFGoITXOOgdHlEiSOSYFFYKeuDBzndQk3XILzpS1e
O4McYeohbVDgMFgOULRoDQHwvE29WIilk/scP9W0h94M6irhwkWWYu4l1lVhWw+j
gzL6k5m+aWN66CQ/IKsMRsmJ7RjSuQuDOn3VSKQhuAIWHTe9v7fhMSn5ZoYOcVZa
yftYY0yfq4n0xNFfSrqiRcodDayd0XlspOTa4De1f8t2FvKfaQ0dMkG+NxBJfr1u
6Kk4a5ih8fyQyjmsks6wwRG/rqdbawehvzpfp0bfshUFRebp/EjLo6Z1ot15esc0
7URfF1fCSjo5q1k1W9bu5LNLRxmvRCEDqxV7rz4gLpBXRTPh5SGp5HdXHh+nthoH
02B+3mQZhzHtrq98tg7zAcEiVzXik5avUTGSJ88Bw3CXYeuLrW/RLev2tOrfCN4f
X42MOAu7AfMOHIjVGwj3/7Qegsuly+por0rpDablo1dJtLToC4gyQomyPCFsDm25
/4jRhF9wB2ovJ3k22f/sOv+rIm0sWwsLoR4upcbl6+5OuHq4j7HKru8VjsbC3bNp
Zue1sVltv98JwxfDlF/6A653LFB4TJTUOe8t9AIfNMs8AQGyQfYB+V1+qT8iF3UH
P2XqueJbGVLEC4+WpxTLjqX3R5scPHz5tEOoPjN6YNA8PoGOvFJdRMlGDdxFY5h6
AoTeTTi0z7HdP6nzQpesk84K2OpNYbj5tfp+GL1YKKCvy7uKLlxg5ghEVLibT7AU
2IV9RQZRn590SrPjm5i9JtNP34W0YgXadqQiJfT7P3xZQ0mKG27FZMFgRagarNqD
o35cGo+NZ7DGY6O1+nRULJOCggkSrqypx9wuN2Vhlpf+XkuxGrlFjJPQKZESEU9k
9ADmAB+gXhiR2Weeq2AARRFgh9+TzS97f69qmZ1PiE0FlrH6ZVrDSHGZmWQTxqQi
a7dmyNLqTFhYMFpCpSYPwwpiLT+Gt8xgaolp11cW3TALGnideluOnrRQ3405cpRC
DxGEFMyFKQXma3ipYrXjx9Kbf1OKe5QT1A5tuhRLtKp9m6ZTOxPm+2SlYg/okxEF
3doiV+pIImIWlIc6CAAJjwjlNeE6mD2NsdFMdfA5L8v13X4zFSAbAJFAdwJOPYbB
8P/otecXETFDBnft6imftgTPYZA6QkbyfnOJekJWOdnSUur0IRqjgHHVSArGYMXA
FsD1iVqgXVcct+E63cgQq1KouexpUyP1lU7tYq6VVR9A0WTemazJpkwVw8HOUFTt
GEPboPnv/VCVzcoVSc5uuFf8mq3TSvCiUBquBseoGeEHv3i6Xmb9qjV6pXQLL/gp
bD/t4QCnF91Az+tQOnNmlT4k7Gl73SOiuNMHIc9C/6nLkY8kEB3g/jLbSUJ5E182
eIpKmMaSGnsnp2059aCuzQ+jFABvnzuEphefmx00Seq/j60ODdGu1QEWa/Cmup+5
TUm2AhVeR/kkdJMuqxFu0FasXEb64WhvCwySGLWjVh1po3x0M7uuLzW5y++4Croh
TUvC18Z9rzATrlU2H8PNJWqrhpePd8VbksaH32TFI0smF5kdbenAT5+xvMe3quyG
BRNPyg7xkgowKS3LKEue45+BHZGDIKBYABgO5/VAOyqjDqPpRbkptyOIZsiGW5m0
XvAxs9FMphDKuniMJ+Muw6WqwfKkNRcLdCTe4oTF+W6mNFmxRnCTXzh09nZUG3xK
vwJehToXoXdgUSOY9LEVLgGKigVX2H6obnbNTwzf+p32qMeDOC7WdLfYQHhGrFOJ
6cD/iFjLbQt2Nkh+A5eUV2uLZ5Y7d3iTcLzI99u7Jy6dQioNgIRPx7zJIodRdmLU
7lN8CqcwHHeBlRCig3FB9M2k35/W/cWXw15rmZUR4jXuGyJj/A21i8f7ZKkpS3nZ
8mkZ2MbrQFlcquiV7rtBVPZuH+2JO53/kPxGgL/vE8jIfEI7facsGl1sNnhqaj3j
W7XK/LS0hYAzrQRb5NebMvJwF9cSX6YImqkZA1DCG6/gAkbCM/vHA9bDw1DE2DlH
zoqZncd5CJwMQ2tVhgK4y39mjs9NHa5zCRcFqPwPZzxqgskTRiDEW/8C57hA2APp
zPQomp/Pk+b0SOZvui/QOyI6u6hQp7yprAFQ54u0P8igrcY80/2YLN/rjpUWCj4e
RN5pMS2XoH1z0Z2IHvrcZcebMfd73+ALeMK4g0d9PhloNwnz99j0XD+vLPaTdFPW
vBnP6KAMXKK4TICoxBzkiQCz7qbauHkPcb/G8MasX6IUrAlPgjR3Qv0O5XasB7Kz
HE5BuVO7N3x5zSNyMj84+Ja0kvfwQSCsdObfE0x1uGk1qPdpobvEKV5S4ufhnsHE
c2pM6H9Mbk2QLet5UVBDvwfcUVJjGx+0ayN5ZgJCNcvC3+RLmNWw//J8FuMTIHHV
H0xTT39VV2wsy8RhkKPf3JUOGKfSQuKddWVglYCuLwSsh3ICJm+/zV4DKqa0eHN3
DGsFmy86Mv7WtYZDkuoXhTnoLKlNy6AIdOwMn2Aq4yAvtkoI225vAVffvR2hGfcK
GIfDgMJvyMxQsgtoH3JK7R4TfTRO/rehI3n/u96XUR8Q/TMWr4tZkya/Z7HWIoJT
gvztpG1nLYT2V765DXhTc1I+gyjrdLlID/24qIoi8PDEi0xNV7Aws3dp+ESenqkJ
56Yi+Q5GdT0auytygzDWlc6/ypC5/UElWig2UVZY0Hy/gZDJPeSSXHX59CEwBYgM
D7cy+VtC1bWCAO1VFMCNuiQ+vTILm5aIqYp3F6NNAByU8SO0ujos7fzF5F2DPq5P
KdhYUeKfSX/j+vrtR1DdZETlKvPMg6Aq3u1m+SLUGRFxDlB4mn+LxM71bwivtjrf
n9n40UcTW5+DhecUO/zBJLXby2IobkLDfDzQgCLh06plx26RE1PMR5C8Ad4WstyQ
87aQKXJJhzYlDM50qaMT0sZceu7MMQNn7IJXYWfwwQC8TFISln8SiwKJje0XAoJ7
1CBBEX5fia2o3fwLImq9T7B3UNDXQ+anxvpIfSOKnkNCezhVl6Hd1OIu7BgZ7zrm
NteZi3//YQrPHvItWG3H7Gr5Vh5CdY8ucZSROVobS76cx5msh8FdzV1wj53xVZYI
FLaV3wXhLKezf9r7JxNmH8OYMKVztqz/E9hFf/JJDfHlARaW7EHm8PCclwMF8Uw4
zEF5+LY3uP2gC6jHCndeA3b2Q0KMQBgeJgBhYSUAz/00HdhblORyZ5TcpntiXRuf
ed98AX+S7FqqV6KED3c+Vy1NUIXYbcoumf3KE7emSpGefVYD+U1HWN6pLRd1Rn7c
LFdrs+Lm5djY6G71JtA+wUhj8m055eJRnjDmQ11iQvRqlpSKZ7ug2ZCYXABgaOWy
2h6j3PABiTCCQGfoWuaK7iEd2EUgVAvVfskTtHlT7F+49i/QgXGw/t1rEOjfIJTO
0wxH64l4Zeuhm5i1W2xgukii78YfkdcAG017Q55/W1jV4bv2hD/RNfyHPYiSTGU3
WPs+kvUwiJXEffzy2hhVp1AHAbDCUEzsLRO+hVOxIpwR0TXB4uvhScglD0d7+Di4
5/qV9dUIDz8lL+Cp0NzDvfZk3hzJ5431gVTk1IRXb2faj/nRVm0oKJxbaov47N8d
iaHJw17shIq9OHUXJT/dbYb/0ELrGNfOenkwQaZTym8ISYqs9ENDXHaro7vRtMZs
aDIlVkAgDqC5z+SHIpeAwN3schAXv4Y9eByT5B3jAvMPiyF/koT5hvCHZLEwaHGZ
44zpjgKHVV29um2SlrR4/F9vFybomNO08XT3AqUtrDFU7TMPd4yf9aDvCvyALiy7
MbWE3sH/59wVe8IIHdfqoopbXBRmxt1TEjCzj4JK0ekUtO68G44c0oWBnJ8WIof8
Xzr1lxP157ZHAxeXbHrButUJij3FPzhpXpSZOT100iIm3MmjdtvFZjU91RO0TUu6
3LdqPDjdazjHFFpP3QsjwWEYhm16/lJL5Z44+lZgLQNBZpVnzcfjEPJJQKUxV/eH
sqKWJ+voLqcIhZb0k7UcZoaqbgEXGycHKndbkbiBjzuD5/473Lu3307zIhlKPUbf
PjmdqcYbhiTVs1I9BAXM6F4lciVnSGTOKfO05i2DdnGnO1HD+X127urXor5hssWl
witjM3+wMvHBjCPamePFy5CdOjtgHDh9Vx3zO9TRNbMoxTYY7EvIHZ7q3qTuPbag
S2yF4cdUIbJZTjWLO6fXAF6voHJYQtHZkEuwgMcVnBP2YEMGf+YJfa1Laoyv+MLW
lTrlO23+DoF7uRrhkc5kt5/xR4uc6MXk/ZwHVY9u4D1A1fWrSfHzFr6YqWcweSko
Wr+vfVHJkxc0icSeKIVWqpvHssHknNdH4Fp4zQVQDIy5oj5Wx/H4hiDVHa63g/fQ
DP/gKAoz/lS++VoiZS9yheffnZqHubV1ghv3Lcc2+r4NcVqZ9vl6XN0EbnZRBA4G
DrQbHvBtAClwNiqBoDjXysbsJy0gF7tPyeFhkk5nSRmDHOwR3cmttUELIHww430E
yMwCnnGkeYJ4kCetqB/1vyz3J4+v4Ug4+WW9xBijaGYod5np1Q5xxnmbCv+1O98u
FCMFpsL2LSnRdZCQe0fPu0IajbAF9cvp6sJJ87C29bY1XmkwHb2Zx/muZPJpWu3O
s0UoIhNyp1bgaJfda/e3iXIO3bZibzAgV4zjMg+Izx+4Me/z2ElvN2/cHeHfCrea
KJn+yqemLw3nhmXySSY22JFrPZIq6wfnx0Hu1RYUgChdCXgPwhfHj0mtcaDHMPbt
eBzmMzFtOPR2MR9nv0UyaHqUN8xu3SfUmZtDcNe+5lplXWXv8VZEEy4q3Ko6chur
xzd+1eDy4mq+yGBeqqJBafFUvjo9s9wjnQirY8a1BASR0NjyZHVQlhhSpMojaqxK
nB3HLBsmL7S3ICSDYyiZ710AincknWpPW6BTCTHyDL2jpDijVqzT/V3Dz3rvoTGc
RaluFwfcnQycamqX94KnAjtjr1jSs8mrJVKWX5bjucYB4ghMXfG83jhvNN/ale+o
P5QSHMbqRJ7aHlVmssjc9kOlbLTGsRS9ADu3E+34WEdPMAXeUGOJi/On8E9BLFJ7
+rUnl8hDT/qTrdY+CJUiURMUyHl8o4CnuhvYRPKCrEG8juvkiKgwQR39bNvU9iii
2JdkqOm7BNijv0RTSe1G8tzlPUkumwCdIU4JqeFZBOworQU69zgL1cxm8ac9dkH6
9/PGqtJeKd1A/l01zci5lzu0H67Bny+XSjUPR2fbXxp0RfNMbauzhaQ7TUXSSwwl
/gju3RgrE1ZQiAW0FBjru620oBojjBN21b3580nfqa6u/zAWnRJ1aVhRewGdmRtj
f+u2Pbwrn6k7w8r7m38dGJwh8ANpmEdm7VBRuqPVfrngjoozSA5DxPcBjlANykEz
+DfOW4CEzJi/QY3HEJ8AICNPR7F7PJK8X19FYCqH3OzBlCpu/yFBulGl9ygE5zXM
D2OUu1uowh7Z6/stFpxfoyNR6B5QlGLX0PpSTPSeRgTZ/jjfrVU3kJeBxxu06FQU
h8TyIM8xWUlm3gm1AwU42rhQPHnm0vbUFCL41+5G6qq8WR+qqCFiuavGdbjA7oNT
0na5PVIhq3g01kyp40gq/tmdIl9t7p40E7kJCkS/zi0kTxY2UxV6HOlXvJRAonxs
TrI/8Uk0BosVMCRS7q04gyJIEzmGCy6BNu9B3FBDottdr7RFQTHRIogZErcjXxm5
pM8LCOEG5PfC+X9xvHmbAbpNalfbOMQ0/A2GieHitS7ynU3ozVQmo5IugzW8rW53
h33HJYIUQVF39HmdAra03Gko0H5256IByHP+KWXla0xA7xPW/3opQXOfhzBZz9IJ
6eLOPKepfzPYJWY+razDmCFC0+8lmJ6zSWAfCqcgRt+Uca0MRvk3DtJiDjP8iD4e
0Cvbrt04cxVJUmvOoo7DkIwMsaLo5YrDxY5KHK9A7vellm7ewXL6M/Apac4LbTFE
XGn3+rUe+Q3AKmw7N8yr23ZK02zt5Or26FNHXsPW2dFzKUwtg/1sMIZ9KBg/I3Qx
ZTUHNU6FUQXE7daqTJpOfzwBoFEEBIqzzQLb8tAP59rzE+MaLSgK9+mS9Cu68dz9
SxfcbRLWrih9I0rSlzUhcL1gq0gnjdtkbYp8kLDHoHgc/YxKB67pFSO5OnkSk5F0
bR7kvdq+OSDhZk6MjFgDAxj8meO1bIz0jvMiowC6toS/3xxb1Q1N1k5UiO6OWQNc
MyA8zLjViPNyA3gkLXWJXc4IyyTjh2/q3KFho9bvFc+ctTYYY6b2lekVApCirzM5
xA2RbDRVE+fI/syH7LQiZqfG0hchCmmlz8THFQGQt3TsIzyKl/Dc3G9uDqiSUufp
7xS/vN+yiTrT0K3385H7ouorz8Vf/48O2z4cBo48/3ymJXjsos0nFfy+iPY6vYtE
QbKH3+9IJlK2mZOwthocjrLdiJGYedKB266LQoa0kZgQVT4MEGT3xPdDkX+QMtkd
iWwktn3Gdn7OtatdYkH9UiAd8H+BDaiUEY9QwtoEOo02vVqM8+5kOekFjhJMkJKT
a0NzAaF9T7phcoEyOnR51lLiXOWd8XOEZeCkx5P8ORVaDORP4qeFvHmRvk3nzU/x
ROyYJSFIfGapVztqj3//mCQe8FaoLd5QuJVeW4trKZ1dJlN6vuXEFYzqAMHsvZtM
wfEld89p6zYoWmNCMwsobCQqUVXOYGL9FqKPHppC2XZCgn7ynq6o9O+/Xu4KCM0y
/HjAzUbDwMq0G7dgDXPMv9G71JUmmc7W7p+YCEGWHwkrD3GgELdVPUhKv+mEciBD
m3nawbKGtYBl2A5Oo/OJ7Em/uKS/zbrZ9Dpa6dps8kRxzXWvURBKlm1YZpAWa0Em
WqkYeESglfbKOyIk4DATRxHIxUtLtstCYwoSRbATT91Gw1aDY5YE6Q0Er4fHCNhk
5D2woOxJ8Ogt0bpa8SMFvyhBAKn7FuNOyP351dHz3t4ukZ0tst/v2w2dWgjuAfq8
PF0OdIOmollrg+1Q1uPZJQqDFG79T/cuN6ZMQWVyH+HHJLSLpHh9JwumyvjCobre
KDyhE0C50h1RP4UuUNUiZUXGdco4cwXU3YNDv1Ea9YzGS5N7ulPZlkH28H0MYTCB
jjaBZLaQu6lyFKh7rIxwipyM6XPiJAO6SecPjaaGPOpc8PhJ1M2e9Ds50fIDSaPJ
BA4Tb/mNWM5jCgtzDz/Yigcx+gEB1nMtB3zvbKMmaCtPiPFtOAzSE0pOyrJ2ck8N
PRxYgKN+9qUs9J1Uiz1vwnAj3kWKohDJFXiQOPoEG1jIP67HERbiZalj9JoHetvb
FeuTXCLi6gFs1+qSQefM7JD1UFV9eV/FvqQY3SgjLrv/95MvNdYZOhhzinzJgfmO
E8OzuZzOxlwhO96s9xr418zaVU9JFh33fZh1ghK5zDj/eDuKT8AKajpKBc2qptsd
omLKHKsXZe/2XScG93M9zd1r95ZMhYASBBHh+hf7z/LADZPj72vbEx9FzJ5nzx8l
E1kqEitgOqNaAzZOk4tjUdbCr16UXRwuREAGxdL8FHVr0TVvYeHfVscU/GfWxFoy
1Xwmxvkx+ImnazjAVQ7qS1tYDI8zhjZFpbItuQQV29B8ucxe1HF43ePyYZmbqWXJ
L8z7SBUr0xpGJkhbuo5Q3B1/KaHdIUIGHJri1eKXJD5vzHtdtRjm3dBvPD57itoV
5p/kEONZex+oPvN7iUMgl+ZQLUq3o4hVae6KYbOlg+rkFQZFZNiAQoZHfa+PwcPu
6Yz2PcolO3k85v3+llkLiQ9EgC488U2VeXVZMUEMupgIVWsDaNnZiZVMO8Ua7B/R
1+870MvR4ZQW2guanNMKXSiRLlsRLGp1S4QuQExz3LaOYh/qmZIx0KFZO7+XUzXz
n1uEFPt6N0ZHbouBtPZn7ejpkVX1C33gB5FOzVHbK8hkOqt6hgysyLvEPzYoVuSg
DMjZ25YiGbnd4LvOTkofxJGow4hMqfwXoOvczMnMBzOfxcYPyJzDIYfRQkwGyX+M
iShB99WHnEEm75l8WXuDMW/nqHLjh4csX4WooP38k8j2oGJ+MQ3SjuBy3Vt0OKDo
y13emb3pM2S7tvFGIB6xn4ueYRAU9I38PR/i8KVbYCy2TNEq9GfItsdmGlNewKMP
V54zLyoQCy9oAsrzlfVDfowDT5P3tYCRt4uzS1z6PlSqMpyyw9A6bwY4Sr3xeGl+
8CM8Qw4G6YPgoNQPwDmchiENXbrDjdnB19FijrGlg+h+ToFL6xXGoF9+PCHDHNCg
ejXCh+bTxz0njAWwdoCVhyghQ5yiN799zvfD4FTOA1injflPw68S0WeCpyS1cNfm
GdDNH0xwW4r0Z8CdmEmUVhEmMZ8oWDCPibgpQZYN712leAfzZzBEiDhrKjtZFYxA
PPnIEN+eTJN32dsIp0ewdpdmDmmjb8ESir4ww82QQLc/5edd7ApvUyNjN2HOoEDx
r+PXMXDvg+8KTGjlFCIV8pfDhISi9HaZzPjlJk1+FbvauK4VtF3Xf1+tKUrC+Vxa
XcNfnmOLpfBd+ofWQQOfa5Z7STd25d8pSyqKlJ0hqo/WUWinrVbL2IHMNqrA8r2v
bCFLFDYx44BGdbJRrm1DRps3KApEIEBggAQa4RKpGmUEqcjyzTWDCCxvuWcSJvr2
Px4wuUzenVoyif8W1SDAuzzm+ObKz/7JJQvJuyVL+ML+hnlQwUUCwTTRLqDa/Dz1
wPbGC2s95ugIxsxTYKAU+hqqjslzWOU0zqf9OB806udXkNWNtfBGGjyhYEAcZUQS
c/qwVVFvF71ZgT6erHvT7kdQ+lpyivvI25MpaPs8qPC2mzydXHXq9MI8TeBR9rTm
G1Rl9Tzh5evugunfirFwGTdDsf6LOpoLamP9NsInRYnTqBSxIB70kc4rO4C/fCPW
d6/3FBG95zhLqYZtUTW8qTe2w8kRwABkcn9K12SqDZ1UwK/KCRo6s26u79LUHFKk
RUEEPnxDSu45sC2CEpYHnyCI0Tc/MvP5flv7UsB068I7pdD2A4vl4x1yHTCz1CxL
H8f4I1Wc+6IHFgJXxteyRaIDsT9fG+Ou+lx74PLklZ0AIN2PFmAKekK6YxP6/Qnz
Qm6GYpBGuUS0U6Q88pJUdjwcLlWwDijTWRwpMnAgOB+1HehJiKZ69cJjvU6DlWfS
7xrUIdprb2YIQISTqSKsiCqTGR9PdgNGsWbvdPUpcha+H2x2FJHR6fQAKHXlvrqZ
TfI7aioUBwTLW684/zes4GTl4drfszDvYzR9mH3roHix3YZ4MhJVc+U0s8hp4uSB
WoUUaOSIYhWgNoMM6DpfDJs/pKiQ8XUhRKALdmuKLfsvFMnGKjA2lUWZ+n+1hPvM
98MPdtAA6mT9djvVRUKnHxsSjC66hfMBRPlYJZvYzm4kUFvlKuqYZ/yCvW7i2bfV
wXtJJauEBfadnlBn8qeH/qPNdDQkIFFWNHItl37YZ5uuhPpoJw7AGPlVgGqV+ovn
slqgtPWCz2YWRYZhVot1pHFQM1fgwF5lFODctzJE/p8DzRjAXQd5f+uwuBKyr+/L
rHNA0+WFn+9WiTJABfMMY8tOX5cUyuJUQWRDF/JdFWlk7TUaYqvpw04IeIrbxqnw
MmT3zLqSPRDX2sVW5rpquUWUdkj8dVRAbwspk9I3usMKdzlDGMo5VieHfG0YT/zw
XBAp27+XvlO1DPPbQrcmyUDlJJndooZstQt+EUlFOE4R2KsPOe08GTfjKuy1LtTP
WZufM5Wwtz7yfKFaYYQJD1Peq4YqRDYVeY0oA5QmLXr0xHVZpdqgur92bexZLZ3Y
k7iM1RULqvjYPfV1O0sPSFvXG2X6FxNV1h+Ahu3ZFoCanb6rAFwtF5mtC5XgOFzU
xhtkeILwr16bDB/eHPRURwvZHJHs1e7O/ppmBMLnfRysANoDv82DqFf1CKJDzQa0
5RswKTplDqwgcRshpk4GuZKXPUcpJZMf8KHncVhCCAc1FzLH+1u7EEMal/rUdeog
d+zW/vQedwJAPFYxk9hLbWQkczqx4dGBmU6oITYv2ZgJf7Gn/BRxfwwu0eixgTqd
ISseAsrTmOI1Qxx0prgj5A52XPsbDl1Xaxf7BkioRUlrEJ2GjURJTANMb4itn/D7
DYrmkbNUEcJfLnOgwYP6ZbEd8Kv62bliV8VRBgujc/3hYy0hyNcviTjOkkNWPPEg
YJl58d9eQnSrPVK5ME8DNk9cpU++C7sSuSqtvy39mkQgRML1moGF1pHDdWEhVY8B
SkPEmsl7wUxaH8SlEnk0aXzsSeRG3saZvooddVDyuvebaJHptCl0xew6yZAUNNwg
Eiy6x3t5NEEpHaEY/IYZDb6H9MJYklwcSnEbMyGwrDKhYafrm17VltuBIJb4LiLs
vWkhgfaoMFU+WLUdSYF8+4nm8lptvpsEWchZkek0DOQExj0CGF7K73mVFGAeIE4u
+uYQfqTugvdwqVBMNsfRN4yXMazjNRPqOxvhs5hW9ryMJWbsOBwjdvbqP+9yklqf
JMKsCnj+dfMtln9aoMIXtCDVKBOcV6bmL4L5eS5t0hBb8kJn46b72H2zGzasvjso
LoA8DF605cGfBuxhkUXRMwJF16Qyr7IX1MRyu6lfig1aWfdlpTKk0n79P/Veel3y
nwJi2k8ji5pog3p0/IbcK0wOg/eqVaLkO5KaxL3DrvCC2xeTp0HM1ZciKw7SzYM8
AwQWguzrLgCXMhO77x2aJX2H0H5dOYtPk1ZLjZqdt0x2EbWAcMf1IbUQJ9GRPiR3
qNXvIMom3wUuQUJk+O3Hgq3VcGwTo2StKcWyky5aVmH7e1AhwauuQQvV9ku2SymN
xav7c46lDIXXR0hPuGTxWCQnyakxP158VYn4kn3gL6IVfAmMuQYhD1oIYdBWaTxf
pEAQ/s27jW3UJxxxTTTrZumz/NFMv/eoD84tR2gw0yy8TCdoX4akwF3i3GQQ/mnp
dDUcST49Nrk2Auk1V9kXTUZ1G/OH3Jd3pmVhqkZM0Ppa/enOxNHwZe2tL/6tnmRc
j/QtmNhXmQ3c+kzBneg14wUClrikxXpb2E9W6YI1PDybgxz5Pn5tSUfy++x6zrUk
/EMd7Ac6oG+2veYgm173KdIlnwfr3u7Uubz115gwoF411ZTTjCCU7rPJ/CzwzWgP
L9SIAjv2WVvQRoQ/vDiU8M8iy+kXrKeRgFdUC0Q6il3l/+IILQU4tbIJ3p6jlXrE
ogjkJ3pGy3qcRBypFPhrXv/g7ebULoQp24ZBe6efokGL43syIDmx3isLVCihMTcU
wAkHRVc9tjKkqwMEIkUvsxgE1zxa3jBcLPnDfKgxEc3EXNNGhBJgikAg46rsfVSH
UTe35j5WJ48ziiYVYQRVG6P0SD/Inus0Codl3C/RwKwqgk15pzyrykgQ33hhwEA5
eVHA8oyMYSR4mXEIMtiiwtsHWKgUKO8BMD9icYPzwpc/hDaknGc9u0zdzEonUlfy
CPYSpW7b7IDs3AnvgQn+cpeHXhaw4CNOpG9Qqf/w/rX16Qu9Cp7IMMX8F3viUkB/
g65R9NGRzYOtGJTKNqhutxdsCipIt40jc3dNdrMF2LI4k7nLiRa+Br7dws4vipuv
LKaCbGMqN/adm2s8Hb0aQgam2ED6rlSm/G973eEdCdbSebsUbt4yFxlFsvCuvxMA
YAtpXzPQnXQTAvjkJ8MX5aH7LJENQmLvzYWnrE61SR7RX1VaRcl5dlyINckEVChg
sQZ4VgiscCDw0vzVrjn1NDYRIaLcrxEDWRraLWtUdKg9KIn2c1cZ68IVYTgpv0ix
ZBYlJRNGP4YY7Gc/bkVa/3z0w2Kf0/K7FnADrmBAGWUgZj63kqyQkXp83ozvIKuO
QfMjsoF0ipSS3QgzuBa7Kr1TqPPGZvxHCRjeNnjCmfeD3N2ZxtnB7qjpNF8l1Vev
R+G7nQCMqJgIRfHs/0KD2bvbodjmV/lPmjsDiJ+9ZilwPRLQi8WifONC/xintQZ5
baJtxTRhf7BvoL5t+ILGQuf1ajpGzTEs+sVuDGr+zaXdaOtxjYXU00FIwDd/5PCS
f79tDky8PfzSy/ZKk+rSCQoA3wDKvs3CFpK+EhBgYKwb148CWer4ZgG3tRb6webB
yri32oi2WI2Eug+6xpy/2AuzGEHrkERwCLMtXydDRxLLmdvMdSekhztjyTgFIuQv
xwWuQXJGBxA2mzp8yAN9Lmz4AIkMTBxDLj33CjPkF2c3H8sLs45pZ9yK51dfHLhV
zkF6w1yjyBwGpTI311cKsh+Mnw6+QcYaVwI7Dv7B26SLdM5ZY86D3Yys9oVtq/HQ
PTmAD+AEV6of2fN1wWCybpF788tSBzd0bPlYJhMS1EI/seXCcRf2+GD2SQKUEmbp
uXDR5Dw6A2putr9hf0nJ2pNBzygeoEK+0bwNKSkQnZ7ReaS6ApJAPqJYZFi5r9jA
NkVIvFqh4FNd+xdUlmz6eybBHwZjAvtZGQYoXUHAjed9avgy0cqRTFX+sj84gzW4
UQ1OQCdzuq87+f3Qr+N3OJ98gz9S3UL+/jNSM4Ns5yIo8+34RluwJFTwvB9tWTZS
zkYleeTzJGCcgaV+HU4adfVw0Z/Z9uuLHrbf58uCKj24iytJsEM4tDsKssOdWQmY
amo71lgTiOR6MnrYsYDc+dF7Wcb+U/m/Cza84huyl0rNtUPe/jU1XnUlTWKJ2a3v
/4nQM9Ad70WAdRid9vDjl0072/qYntmuDl+KR8MTf+1YBsuFgDLjExOa1G33kZzu
B/myk4TYmmKsvx9NqVGzXKoRaOU7fglY9blyZBUdoaaU3IUO1Y5XQ2uZve7a4xla
4+u4R2SbMHXIiJk9dYqN1s7zmUJ97eJosONaAFsNzV8KLqAXlfWzCSGE7Z4V9dov
4Tr5/ApFI7iLrdTBGz9E0aZWpE3mfKFj3Zm6CHuKVSxGwnu5FxY7WbezYlHSjnZT
pZLfBEbVajqNLaFcE+2EYnk/cCli70rWo+98a1pOWzP/TGPsSLM4/W/CiVlwMGpQ
Qi4II0k7wZCPDr/OYtMr7bd1rdnj90wnlDdQAPS6bVobaVKT/MwNcODBHpdx1Spo
xUrCOwRIrk3BYz60gUNRXW9fRvpculoJ0VuhtM2N49FmCK8BtQCEVvKAcHs7ASmt
Zu0R865Iv5Y8BKFBXF8ZLo98xX/MMb8zBIEPqvv3RJFPW+Dr4fiYntW5zd+gVXra
OBhgFEMwklfaA3JVAlA6otpR7ZddoSoqhIF1m541Be5OG53cL9ZlVjkAW6HiLbBP
cTXRgTRsoA7v9n9qePjq+vqgdDY5HkazH2n7WEBdFmpkZD/0pOl+FCqiBLS9WNQW
yS2d5s1qPBZuqnmqb1cQIqqmuiAPK/J2+G+cdQLIe6uGobxduuTG056wKzktuD6h
MAtSJ8I4BH8MBEzG2L9sIxavhJvX1KWbStMX7TLIehVmjkKAbqZMTmDJfF6VGPwi
Fv4sohxukCU5Gk+YOf7EBTw6mrFXFdm+OEF4IDXbjAQPhRn1RUQ4S5lAKxgE24g1
QmW+nTPmMR4rb9f3lLUNJCxTyvs84LVtPSIMCDAOWXj2XKNzssGQ8bVj1uOx1+2s
hTC4H2788Nmw5SzcCWI7+BWNoWLxmjU674jI0nD15OtoC3AP06UgLx71Tao6AjBA
w9Ok3Lpr4XmhSWp9z4pz5FoZedKnqWX5Xc3hPd4Ytr21IHKII7UeuUrFfNOSn2G7
4xhi/DCb3kAhXXWR0ftttwAbqE67s0ndckdOiGjI39p5AIzgibdK5m7fko9j9PY/
YTPIzQ8iSEALeU/bm3dkW0E/t/Y8c4LEeh3AgYK5uSf1rhN2XcmwP39andMCf788
YVPyEzlYJwM74/XSwjXAzBcW0A8oDRMWygB8poJXoie25Dbv4i22FShyIcWc4KYE
A7QqkJhvVqtPCt/hS3KI5SXS0Zcme6yhpajmtHxsQGdJo74a7wptTfvhljnRl6tk
Jjd/i/EhRgVxN6TgLmlW8jmE4OAlv7zpSPNMHy1/gdWAtWPAme/4C2r4KXRhUPYd
aNDRkaFVAjYXXt21L+7vzIpcnv/Be5TVb42+groPSVYDy1OQgGJl7RW05WMeh4om
0pOMrfOKyDAjaa2GFZUwzxceHBxbqnN9Gn2vBMk+O24VfGd5aml81zLu4nYsdISf
j11MK32pfkNDba7fX4/c/8g3bQl1cSB7E9DR4zdJxLA6aNarc4oGNQIFmb8g3w/1
2SHcj4FIxEhQ0KqGXCmNFALck4T2hDv/yR6aaUZmGEYRfYSOfWjJImChhvrN6C6C
3if/hWip/wepGLKDFVuxKBagMBPwOXSthG0US+j6VjGyEnXlR+lgi137vOUdatjh
/IOv+I930DzaGwe3iVFrBOsVJ86w2jMEizv7S2RS3H5TsEzC0h/7nPyM5xsjJ3Dl
88QqWk70GYBzRkwRznE8iiKLysEMVqgAPTxkYwHg98qcP28FNF1claqtWVQecGxS
fyWuweerROBtFfQ3n/cgpcIkj+Kb6Sq0MXrYf5bX1VB9R0P+lxMgAUp0dYYyvVcD
73RuVQhLZ+SgcU7yPEZ08RDGgHqjgYbc4GmBxdYVVhKceFvpY2lcxYVLhPHl7gTw
2cOql9t5pvmP44XButzYyqhEymlvlDMmvY12Ik1RfnVaLt/SYnnUvw+nSRu6g5mI
nU2Q+WACY4ThIpsyTnjEIvdG0zuwNpy3hqGZgZGhdujZyIB+iCxm1zhA6igpdIew
uZ0j0Q+WvClEkXagkzVQ17sp5Ou0iNZcC03aF/VexEmgWu54UtRx/fOh376utENI
yJAa6cJkFEs0XCpv+5hfALJwZcicxFB3fiE0Yk/Atb/Y6u1x2MefcvaD+sZ9jI6o
DhklmP275PRqdpdbQS5fLtpK8VeU8ys0UHT4y3+GSuulufcP49ofhuDZsADxk7a5
MO+ofyEiMZhuYbHY+3zC7WS7vRA5rzm/jkbb3qr7AzE0nAe7KNvQ+ubNX9cxDYoY
rZ+mXYdDCuCxkUGbOtHAirlO1CvhtQC3SmkINVFrMg0ouUZmNkekasRSjHe5SjTz
+X6OogfMD57AdF9afr36XQkLY9PDnyx3eSdnb3ITJoBLE5j5JY0fVvSxzrUEBti1
1PntlkEOGWSLjkxfRFMQwYwdgbKuH23/hE7GE1bQxwkdAPtoInY7S7NwpxPrsPMk
0apRREkriGXco/W3b3EUijvH3REAtkMPHKydTnIXYSEZjEPm/WwUinU3uzAVA9Bh
VWqE6U7qkOJrGZh63/AuQTdazfpqAll4/JtHBwH94QuGbb1yhMWAVgEhFJaAfRD/
kfd+dB9mSLX0uYLnQbzrVU4xvUk6qnomqLqB8IVIhgID7oGMIMjGjoyd2DKdl8fn
/yHEGkne7Sen4yjSJs08tx1VaVtJl7hIWLAt8/uaIAxhrjgyVmPq9J1NIZElmrfI
EsZ1R/scu7pEkOAviZ2vlbJyicuSdXI4G6octv4GtkEcIurxuCtRTkJmCzgCeoac
xiDtA0GCzsm6ZnT10Ec8+l+q5jtZH5I6tvcoI5CYOcpywl7tz99V1ihxcvs5xjNR
HleaUkaPdabmRLDAUjDcp7KycRk7qLCvwPj0WDCJ5isR+jVzaeO6f1Dg65XpWzx4
xQlIqY08rpUkIb4PLCXls4o9/dwchuQUIjfgILK+lujHO39hY+7UQg+K+ihBt7gw
nSJrIQcVhPbA+FQV4xjMPbhQdDPlbtNeiw5Z0+yRXIoLYBwqpOCBe9NxxDXjHyz8
qkgkLvHnOgpLWebRitaFz5DXIaUrktt/pngHepwXV5sdFAFPmK2CpxcyXEyoxiQg
8bl+yZxtdXyFhaud6yVgFwqIsBscN+9dJ7M6uTvpdmC4qWDKQuRbA20zgQlyOt0c
HFa8c1u6HpfnPHzhWzu/0V/KzjcaR9Mz9KMn32YdaD0XcSxLmpPERBhvAcIli1XY
4M6PLVDpfp0tbjbUI8bMoQ5+rGRm44Jw7jd+j1dFI6ERt61MpHnO1d/42RrKXMvj
02Ci6CRXqirH/+IAgA+36qktRuO26tx6Mk2ctv3ZiYkI+go8EB4bdOFNz0x7xj/e
E8L5aQ3xDAWVaXMq5jvLmiHhTUHE5t5kG6VqkXUFLAGVNAVdVSgnyUQwhI6TsB+L
MbC/qUkPooH+TUiiZTuRpQ1/4QNdpfiiUGhNX3j8Hu+RQ2nB4jj0Fw2+jsvrlday
c0JpoMdjssRL6UQLi0Zo9E8Ed9ecg7SYkDDvz9QXLIjvnTdfVOaT2J2uGhU/3dWH
mxOj2KiKuYHG2BvGrFcTTB/5nWy+NDJoXimSKRFbMyOIBWbu46Lmm1NX7hLM9374
4vZJwYnwgZqiW5eK2fIwfFgyzxkdOMxOJxMIMK4JlwjCsv412TakAIz2ar/IPWE7
p1/nCcNzjxg0/s1XS6tGt/B570zZwBygx1Q/HLoRESH6DKJruCeogIt7eN/K6mJG
xeIOhq/guMjY7I1ymgsrlOLu/FY31N/2n/kiPKYNqPrd48JbvFRmlb9wUuN/Vdnw
NNL5yAUJS5gPaB8p6VSn4OOutfNIWR0qB5BTD4HpxF/wpeD3KW36VqNaKwh9E/cA
WWQJmKDi5trlN9C59f0EPV8Cf46EzmhzVYjb11VtThfKyA8YihP3joUV4XXhaGxC
8orpWp38b9y+mPp/hjzii2mYi+Ih+mFpJ3n/lsZS8rNwpf5Mrcv3mSTR2O7d8BtX
iSdBjh1WiOPQInSJ+Zwilx7DLG8aWsljOKwebFHtmL5HpZoQH8VhJXT29a7eEo2S
2BcQT4OluQZ2s8Ysh6qES8KbIYu0u68nHlcfux/RfAiS6yIAUlw1h8SG7Y9xvlOU
NA4ozr5fB94TLo5rXDaBorN1S/CR5bW2ck0CRnvRfguu/CCMopKKFjgP8w0LgF88
bsYZ16Ec6X+ZywKySjNsj38KHGZWlmIfeCLXx8CZdmhuvKyTE5GASB+7Yz2+A6FQ
i+lKSyBWIYPC/PcAU+V/rhwNe8RZPxbNopWFoAwSZTJNORPl7KaUYMB3Ubc/KowK
4QeGPLAACGY2zzFtTcwwYcviKod5h1x3FB9VlwZTbnJ4LAsgBDKj89S4/LS0Gjhz
OVpe62ohvvpiGhI6/oA4ng8msCXmaiIfHGz6VIGNy+eyTEfNo6G/lKSJSl9l6/oG
n++t5T8J2HLgEnmvRNVT2SeigNRlAlzG5iAj3+qMUqA2ZwIzGgulDxGcLxNBDMHy
Eh3UI52W2hC0vO6iBd7h4D4BMa4rqIP2lDqmg4gvdmW7odRGEZtm/Fjwmiq/FvX3
FLFVM/lik9g19/Kqwvof4izE4uDHSh7i3qyOQ2RGKm4yNjg43SuJfjAKOaJfVGNQ
ghqw0pSqOPDt9WH7Wp7ft5N0Pcqkj/OfnSYll06wDRzpa9Mglt+F/LaPJXK8ox2v
hQU6yORRME0UyUOTTpQgns8yTENYi5oTz5BmxkMeDl9HSMKdTxFqGN1LmIdostf4
oMpc8O5CBLZU9Xggn0Hou2rYVS8nkNwkw+tkic71naKRcjTBNbKaJe38No9KhoeX
qxW7duXxt0deJ8GdGUWlDUpCNMvlmeDM/oj4XNUWF2Snzx0UyQqjTJTbdjv8/KbN
6VEIJymFo6rp4Q6igz9s27/jJ7IokBx06+/OSsDNaU+RhicgJbr8c1cHSYSyZiO/
0xLBn5WX9VZt8Dg4oXL4CLMud+pB3mWamnDqaiOBSS4iJQr/W5YSI/HFzKsE42+e
xr1Ufsg220VoYWq3cJSZ+fAIrVfIFsqSXsdhkKNp8IHErsOx9lj/tkALnb4a0vyF
LNaBP6ieFE4nn+SVyIWQVSuCFfTJ9X13G90ihTNPQ0STb6oU9x33JrTqaNoizgYU
cfYwb7Oncc/xQHAXUjRpl/iOHKjTqMyt58F0Pr82fJZn08sfuTHM9u7jq9wojK/O
Zk9vp8pbL0AHVByohHUDtoDndjbtjHOkieduEB+ZKYlYgdVoi1Ntx2HOslTyA4Co
TB9HqBBIcY+VhYd3eJoF8KFknAGkSLnPnhUcqjML7Qg63xXEEIxmjS7ddmZ84Ed0
cDWEM6rbzum4sYGr+DSZXeqJWPKFei2NfeLedqh7dEbl2AJObF9xeSzOrjNjwzg5
MRP6EfA3AYmgNbuVi+8TJWYsYTcB3j0IJjFdvOin1ijm8D+mf2hAk9reOg2Gilll
2O3flM95/aYAcJxqmnsbOXH4kfM7DDbuTVcX5R54QJhZnPle0q+ITgjybl6bJlao
eQuhIDLfd1jnKNPcRN2mxWyfHY16+jIyPd5Y1C6kSSGRyzlYHBkoBmzmVM9AQq0w
/2RGu1bIVbIuh1q6UcfduRY4cY2W90WpB3I5529Cwa2nyDeyhbLvgcaSTsHqqbG2
Lo+3XAtfjjqhHxJd9XbCrEh8srGekyDTK86iUta6GmhG5qhDD/wl6FZB6yBvh1Vb
/WLU6/R2OeMER8JF3woZO2A1dvttGrJj/F5WGjraeoOUgsPITiEXyOYDU+UpAo9d
gxb4TMoZ/y0bFQ9VB2G1d08ZQkoipCO8OQz19qendIc57FzhbM7BWcOPhnbB3zgo
rjEcsF3l35VZ24Qq7pQCLP+yg5g0694YN/sIqLVbRkK0xaNXQYdk25NEhT4hrJMw
YcD+T5zP2ZGbW5eJt9K/h5WrKXYhI73MHQzD1lj4HCQc8nFAEyDeB2oD3Sv+ay78
f9XQYxw3jsz94hecpnwBohfnt1G10NkPw8bLGP1kirNceF4fd3nQZWaSEUTKJy+l
ZXNnsnmrITW6NzFhxti57l+9yulXCD0VcIm+Mj17FNcQ/8Rq4JykuuBN4YAy8Ouh
EtpdjFA2pMf8Avi4QUfmnqytXYNpncSnAiA+Io/m95nNdM/SKoKo1RxCGUqxeTOv
HOFRABI0X4V2OuSnoAQyfxC0fNqTFerZv7x2ENXa4ZBJGwoW0VgNxYvaS5TbtjxQ
KjhM93VH9hHf3EhhpyMVaVSAIRGPRu5qIup86qwU/n0xRbIxw4cwU186a8MtW1eK
5W5Xjlh8gVHUfO9ETjYYe4YQ5MfUGKKZZtktkAk8Qf+ms1+X8T69nevtnpbBOnWr
Dml9hWt9OLhppIduUqhdsnmGhodTvDr4Zg8tBQRgCZqwGaYSwnIUcDvxHtYVsDM8
zkO4zMz/EQjBcWDMBdvMsW3dYle1hszKHt1enxJtA7ByeybzDkgw7bG6eAf8YhGT
EVDH2lKKGd2jwARjcDXKUzZrAsR+Nkw39EgwuF+AF848ydzg+PWE6Hsn/ziB9S76
+h32mI4zA3Ss6c6dQbWwlRy3mUUYlKHwmnQzQMIXZKh8lwz9f1rclBpv9tFt2dd9
krhRBrK+PhdJwMgavMSJJq46/YyGqZKl1i5YiE3XrHDqEfOXZ0o7dHFrHgaw+Rin
OTgBVWNidQXfDMxm3Hh3ltH6HeaYk7KGiNBR8n+GngJKfielvD4iAk/axPQf7vSi
lugDfAK4GzaBQNK/fabunXQbTq2c7D/AsXpmD5QSbot1AUh9Y5YBz+Xv7JiTPovC
Bst5o0nWGZm7qjAf3HkzghhnlZ2xFXU9kAuTh0RJYTG/1w4A1i3Gl8rC15U0GHGA
IF0QjkCq2hVL7Bv7DLFjPFMPAHX0JQtUwsQwEictRbaCMq+nrG0Yk8x4x8XCCa6j
2SLOpbjtdgiZdc2pHWr27vHfjbNN7t8n2VLcg56GyM85B2Ox+jZ3WsodmaaJ0rkn
hTdWXQ+kmsrUdHuia906DAm7NoKGJuN9uCBnfKGoRwH2aDU02jjixN8ZafJBkh+y
jlWoiBeVDkggzS5oTiZFNp8CPItZ8e8YT6SaWT7vcmh4mujI/7LVKDIKT4GmAZhI
vOxsuU+HMs7hzO9ltZ+DgNYXNJvNxt2EhPsgW5BMwZwyrLYv/6lRV/mfNdz7cLg1
hzbbU03EosA4d7sto9vSOp4x2ObIC22CYP7ISz40HwesYKbyup80etzDr/U7fqj1
l69RXjyNYQQe3lUsE2G15gooF5vdmESbphrsnMeP9rDKmakZ6BysgpBazgtMwezy
RyVtREa9DXlmUWNbyA1QD44NsN363GGoa5E83fRJg5/hPytIebJWnT9+hhk+Qf7L
L77q6pvGd9fidxkSGZE8z1F6meJsBJL7juODfU/yBiQN5BkwTSlmgS8W7RzNW9j+
OvIRMRfi0YF+E0a1c0QdKXhAkTuy4sETe3ZCiEqADwX+CK7V2wiCLQINtEpsBWTH
HnmQoP/w8NWHL1keewjGqUWbIwZ+g1u06t3+dBz2aARDx8Jbmhf2ePl0aKWLlFYo
ObwSEhdoGmPP2NY6dT8I4/R9skXCUnnSdOUTVrxRV/LHrq2NnnFJaStWy3sG1PMt
Jb7sJGieUOZQYzodVptDym0VEApVzRLqU6sZd4AC2X28PgskNnY0MPqJl2AaC5Cz
jRH+DEY5pl6iisDYuob74SywJBFmdNX6obfpc6DJVSmZ2zt7mKz458cN2HrfBej/
hhj5DeCk41NtlSn9+5Rr32jICzY/wKEqUJ4aWEWbGvgX/MjgbGBDbmk1mod6HytL
sdp/d+QUdDOwRtqS2bXUzCDruSWt7flA8yMSZM9Bd81hS5CqLdxiiboVkO4FRsgO
PqttDWBKfro5YR+JuwSreV1eWTrkM0EaR9kJvCYsXAttgfq40C0dvXbb1wAWSq1O
iM+edHqsH30xSmaTqo/gESW4sluceH1tY1XvOAVfDzX++znLaZzGHuYl9JaurGCj
W2eQ98BFTWM5uvhvuk/8biDTgr6lOvNnCWKUriobFvFI4AofZBR9ajFMcA//BZl7
KcUHBHm/ZeJJRQxMga1s1yw2f9X6Xmi/LdVWiNgHK+ZCa2PdSE1xk5F5+9MUSB98
tbDok43YZA6njJF537jQ74Q7kdtfXgWsAiDeYGKBAfJGQcJx1eoB+FxgkPeZTJeO
lMOsqWyGiIP1m2odjYO9HBOxE/PXRR84eyLdS/nqFiwuu839QulkZbclU8gtdzTd
+Vaap0pTEVRswUJ1/mFpEokRZpXbk8ebZlMpwsCBlG7/uDYYj3YFXXb0PfPKmbIt
j6VmjxlPB5HI4V2kj7suH4ljHHSU2lN6deGjC7I3rKJIt5uVHv6vza4p117uo5uv
210V2eWfAQDpxvRJLhTGSwcrCoo6AMDumxTmVdqUkblLWHwEuTN1IQgZOcDoMCGS
aHwpdvtuX0sspgmahIfLJB4uP+h8xTviJfyhvAqnHXqfmTnrdnXTuWwGfsqf0W+w
Y1TebEHhOCser9qf048+8K+6c8zuVBj0fQToxQ3/sYz6k1/WkXaRc5zLZGWQ3WxB
MyhVtTWWI8hhZokmkl1vHlp7U/ylkYrE77nzjLB6iW/f/M9HlGNCaI9GCyeHCSxI
3jYErFiW3LwSGJDy3lKH8V+fOrqtPQBeala66UM+FNpRJiYygP24KqRk7AY+WsQ9
h7yosERtcWmtmurrZoLYQ/jQZaPhPWK+FsuFUJr+jiyM5dE/lVH6+wXRYF8u+Uox
VzYRh6VjFIqYXO5KnUtes9CbTiihxkx+xTpqFQmMPqdLAHvqT9V4qslKWC9nuvl1
5TotxoZ4B2d5hfV8kDNyuf9+zcTwaUr79q7ApIgLAHFzFozHmHeTFc+g/fRguU8K
3X+2nIjStSuBpulOuS1IvDl5pZR3X0R7sWxdydpL2OEtjnsxCRDCK5U7MOIL/fMN
WbJoID6ClMmZTDG8cVZMW0i6tBszSf+/hdeggC9R2cZpGnBljSFYSVHZSuMwsATm
CZNIHaumnDyiY4oziEYpbkdWuyfSkizfAWOAanlfy0OKcADLMwK9iubj38JdEXgS
r9V4xPjxjftpe54/yGg/uwZNYNauVjxBuOhNIvgZaI+GScugXQzSp7sia4pacI9g
KHTtZrMw37oei3eyd9ZhgKPmWZT8byGxzrosQuodEsCWOl+a4f3QwRPSP+U1bT6O
/zbau++Xx01O22niti+7Sl8Jr+NfektKKPiOZWfN9z1slaJsAiX82Y9biRnM7Te/
WTSbg9Y5YywgAxioSUROIR2fyD6ikE3v04ErNKQoRaGrOR74TMNlgYKtAaHsTBO5
Sw92bV4waS7W/IZdoxZqDY0eTSMhrK0qrKudFLxh4mukhE1DePBV+6AXLogYIGpa
GGJQppzPomJl89Jv983r/Wj5quReL2CdyEOY3yTP+Yp+LvVzmNBxmgCDap8OWVi6
XBu18WujjjD6QlbLWWolzSANKoKPth2tSbGMGpNT2C7ABa80hgqYsxS3qysjFITI
6pp98LuC7aaLcSzi2DZczqlHCRpR5RZEpfku+lqOapx4d6Sli/pfeVViz+OVX1Le
R1dqb9QziwdFcoiRghMjuVtlGmplRetGPZ4DS8DW82xGDAIzRBjHFpED5WelyV1j
jU7Lo46r7zDnskSC6uV4Ff2vyHznmUw3xdSxy0zSR0tJxsvS4dtVBGorlSOEHbK7
9tGHV+mdpQ+WjxySisE7Y6rkeHNHmekRazgjamQNvpWPb8nuKKkfYC7EekVw5qdG
FwVJe1XeIIZaFUQ7+eSsE+Y+54E/ECJqqoMG177mAqYvhgCD0VWpCBXU9VdK1p1m
jiTqVpFRompOjwpnhkuUM97SFN1r+XBwtkNFEiRyKmZBYPjF47ggAcFT/V2DO0ga
8ec2odNIHamRKOAY2rIgbBAD04JoHnSekt3YyGfub44nKcv1rsYdoAkawyk8jO38
Z/HFBHZ0/LOcFySIa6UjcGys+G5NGpFKEaxfFjptB5PrIBl382KM2GZXj3fgSwVj
/dja8flLandjNLV63zBu9fpPq2F6wSxW5IDTh/cRVXO5m+Ltbo6XkJUVRpiYWCt+
rwn9HWtYxdx91L7tT7ahcLIax4fK3pLyWXuHiySt0L8ywZTvfuS+nv0cgBq81kMM
qqAeDIEtRNH4DwahQVWWSp+173cCKqFAB8s/apPDVqM/mLq0l+2hJjfz5pQZED0z
3Yb7C3xBYyzqTwm5T8xiPGfZPmUVy7vsO+uUVqGwqA1V7VE5CbV2RydzEpqeNSvf
bAm0wq6gSdyFxp7nokZ+E5TPLNHBhMP91boAdpGNY9/Y6aaZ1MLmYCfpnc3CJ+h9
AvPr5ZxGdKpLBkB6C5DGHafWXvUJBpwz+PO8M8PHLK9yHo8M0qLKsQOx8T1e7kz2
4egxbUb5QG+BwfiO+xJ0fkOhUOzf9nkb5oRKrh6ewvlUAhK/ZE9cF763zxv8rvBq
QoAs2kbRrCGqymqp/5vJcbxPcTyNEfDctu2AXdD1JqOfDhkU61Ci/a3yCRZaODD5
qp18XA+0BOe/FoSMfV6ctYMD6q5G+ab9Lm+V/1D2m8iSP/J8n+Uq5JUQ02gWnWmG
Hid9Hxec5DvbsQur/pUXR2SDqAGD7eE4+IkVIF37uStedof6Z+ZHMRjz2g5kqT4G
5lU2Tdb/yqFVmAznuxJXaj5TikJWuIGS+bgidfY0JOjXm4eMavEE2F21nsCDNdX4
CcdUPu/W6b3Dt2RgH3fBTpXBVVlYYt/6kmDz77GGwto9gS0BdnKwWJkZefl2vgfn
Ks+xPdBcluShXOHpfCvcHAWkY32vjAD9AiNCO3QSLkCVSIyV5jcWWaoxt+zHxJHE
lWqujpoZsa2CNFZA/r67XKazAuWbqLqbtS4WuWBjW0wYXLbjHixKY4AKC61EI9hB
1UJpnLR2o5giPNqDsHRnMu80GFrinO7g0IlF81MYHdxtK3C12sq/5FaMDrzp3nFR
GCohMCXqAy9R8yz4x/G6WpX+nRA9z+rnHGBozI4p1IG12HPwPRbUY035b054UaAO
Izu+JHr20u4sOS4JJniViEkKfU/cNIE2MKyQLda9L/2HC76jwWYjvaiKIKiklFs1
X0ahd9TjTXwzUu2EolwDluylEPaxIQycHhC9+jr6LuCAUp4CHYTU3EjJmVtwXrqV
zugskjywe8sRVdwB3aksPmWWP2UTm6mOjy37HwlkJUX2FP8o2fUKaaqO2hzqN5Fk
HEQIsUziDYy0OcEDqvZxBiFRKVKPRdiqK9KSv/SolaRU1TLklX+SLWHoThhQ4b4n
E5pJp+f6j6kVxLL09s5kIpJoCr5sOZkmW5OQhWEZktJti1nbzsDt3YxAflw+ZGSw
6hqeG9yEVUD9IPaWVe9VLPXM9yGBuilI2oexJW9Ig9kcIa03Q81T4sL3J3HyP8vQ
cdQ6egRmpjjKhAGR2u6PIcuS+WQVne+0RZX6kpHsf29juyzeQ6G5T7iKLhefZ3ct
SGy0GmbvMsfUBBRKvv606n/evYosSwUAKzwabwyILRF43POQb9l9C4YTF+jphNNE
E5dbxo/EL+QnF2qQS+LTen3YodF1KNHy+xjUAczl89MFnvwC9PUaSnVT99un/XAy
C4XqfUK5Bgm+JARR9B027jw34NuQL9h8b2yTFpOB+gmLpQbxzFea1wjryiiYRH5I
cIy55g3oRKi3Ob/zuutXBxBeUJLRm1hf5KoqmHtHpt0XklyxSjDBe8Xn80WtGdbF
yFkIR+nETz/9DDCq+Goj+iGHgh9GohE1xE3PT/AG43peFsiV76dvcFfd/ZLZsEfX
IajsvqSCnaLAuZt4NsC2yhmCZ2Vhvn81eC2tQpUEQYUfxY80vpONFqu3My1rqFJs
vl/9c+zY8h2DqxTbR+kd2CHZsh7fwKlyF8x5LRjM6o9R7bXB+0K8FDs6MNnB9fiY
LR2OxZzK0UG7fBWOp0B+MAv9leEcer0bsUq6YW9pFjd5zvz0tYV1Jwf+emUq3l6j
f17YQKn+KKrDR2zweZCcwRDYzPr2ckjg/8dnK+gs99u+2DwA1xEuqhwiIq1Wrr93
lJBIfCgKxma9lUv3NL0d22MwxTsWnLCIde+HtKRy99wrdLG+4i2+WkRGUMzYz24X
U9j+LWLHrjqjxSEq2I1jnAV4j/1aVsxDZRUlBJDkqL6D4faVhppny8H9Ylwfx2bz
6gGwiRHgN7xTxC+VsZOUdpV8+CbQqe0IVicoY79fU+pXKDyH5+fqb4rhaXu0Y4KT
tDiqGwUbfGFnUQP0O0ohegBOcOmduk/bo1NOYm2qqYQXUKV21F7ueJHkn6+Vuxrg
m6Qj19t4wuZb9yIq4OhAQ/2CRUQBRKnjW7gK2WoC6YU4tNomHEt41hBefnQ63VZn
pGtxG3fQnVnyovZ0VJWWvMgfXWNP0jzyZnMTdDSLIqVN1edCd6cBJTTfNW4ssqmz
rMoGMW8Jn6dCkLKCEGOBYFo8GzEvXaXaW/vXQCBDyte8SnglCMRgkojIBL8mZKFn
Lit/nppddTXzV1Pc/SicBVwsVxrMjZpR1aJm5uXF/aIAFsWT33DXx4GL1Pb/RzqR
BsKKZFBMjasf1gTtzUxB2GTePGG7mYjhuTZnynHZ1jJoiMM4bcB35NPTw++J2GrU
ec1Ah2TF6wPO6I84v7pRtw121tyYH+KcMtPfxSSXKr2zDd9wQUqFe+DvXMDO8qG7
V3ncUtAdzJu0JxE4cZ6aGIsQvFPRzONMxIPBYX5mBA5gNCBue3m9lB5Dj/k1Jgjj
0F/9nNEZe7k5AHjm4kToygOJ+Z9TNK+oIW/lMqV867rd9rTcSE+GTk8Kh54y73Vb
uj90Pdq9Nda6vBIjB5Pe/XnXFALeW/zmckIf+J3aIs7JPAMlrDUBIcRfOeSj2sSl
ms5L1TrvodBrHQciDyldw5HUKqlsFXFkDPKhOqUFs3hOwOaR+/+yIjMDNP4EFtbt
t+Ie7EGSxnIAsDYWELpYeEG760eFlTWQS8I3Iclfz2SWGkklI/Jr+nOuk6MO+w+H
0MFzMHAHKOV8VLogZ9gYdB7EIkd0eDwyVUVIjrLaXaMDHRSqrUVus2tYt85hZBHt
9WRjk95iF/QuIBY767IRZTbjyeaY2ROr34AdHO1Yh7m5K6IFCfbLTQWAk3y/V9wx
H0SawFCUzmjSou2t9nKJi4GT08zcsfoqTNMTxvnDLd0OUvZHc8j0x4fYAg5hSemz
PfTStEHHfHiK6+65zynxcliE0obk4eAf5J23vUmrJmZoqNXbHxK9zvNNP3S1uEB1
A0VLLcHnJ8j9CJofE6PAgUx5uHxbCqAn/hfIwZzHWlOqxvwRGhxYWeLn+0eIsTSl
3t/LsbZsVWYSJjFnP80cofLpRS+f/tXNa/Mvv7HjUgeoVpvrazsW8u1aawxzUIGh
xR1/5OXT9f/Yl5ULj1qjUYHkEu3pn/3QldSHpBhe1mqmuGq36qsCApDw92f1DWzR
6FgrWLgcvPl44IdiiyJ2HG7UsouiAG9sgOF63bQ/LVomKCY15eRxzbkD9/GL1SA/
+sVXmQuuTbLNs6UtmecYEqWr0ZuV+FKj9guJKFrkVwMkZXwEGUyWIIEIr1fgGkGC
QibT46uqozEF7RtcB5lqRhYru2CdGlmSUE1Aia3iUo8bzJsHKZszVzjqm34kreiZ
yNJrZrbW36j9tXKgwpWbF8sVpw9TJH4NJr/StCFSM3Iqdrw/Pjk/qB3dt4UlGas5
BY4JbI0Af8s5cEX22JQqBEruAyH7zGttRLQiywF0ouAY9F32mdCmv2Zp3Msm4WZf
d3NbTAsfP2OxO6/JfwAunsH5jJIjX/QyJgDap6QESsuasddvz+SHiV0hO96PVpDR
J6+6BMhVd08N780WV5gCR+hoeRh3INwaVNSQmBuikznq7803BX4Y5nwEv+qEe9ee
ab8oze0OvtLlpdSgrn+C4ojF/GazS7VnRaXwv+CnOf07P4cFR/cUnwfoBrWywGUU
tBgnGS1T8foetUy4C0SN21xNK3mUIdtMw88w/oK/tYmuz6wbXYQn6n/445PdaNhQ
Hof6qOsixKirvrLwPXRYlfrcdY1Xlhe9QClu3/PZ4qtggEuHqwndOydF/9jAOpsG
lVZQoMmcquExwDRyIR/mN+MqD/fiL/hEolkKYaLCOwC4Hqjv72lrgzlj5Tqq4Rb8
U0vM8MPDxBIJwpE66kP4FHW8sv3Ru+AQQzZ3TyRXrusmk3oq9RcnUKppboUo2m0/
Nu5FV8M23icTOG01UA3x8AkK6DXxK1cFdN4jyE4tJMyEoGfI9sT3JQB5BAEXLito
ZZjU0BNEy3ZMrqSH+MttuUIoYkNNMvSKRnX3hn+JUCbRkUsvcNDWGfVQTMXeRYev
17d3AE4OUaK/qPPpJ/xp8achMKA8A8/m8LlQiCQ30XOrrmAA5q1TaEK2BR7RYXt5
T4zUN1CLGwZti2Gd/qkExIiGkF5/YaSGvyLCRyq4NK+pnniPKJCoRUvnfHbGyyTk
x5LpNrt/A4RGjgLt54UzqCPML/2p8/tV6+55VtPRMdOVshoRhgBjDOusbgsdji9U
gOGyu578b6oRNtwIQrhKzzG9SpQZEvrxePZFi5jzkfZsnSpi647sQUoSKOnL0yit
DOKlUp7g00xb9ejVuGwlTfcOoPVBnk65lWRnrLEhXe2Kn3SaRI3sTiiP+Imyfhit
nxPq8uC6SNCBZ4Ok07rmjnNUF0rKy7XbJf0pQZrA/qGdSKX2HDqPTKsAZyPrDQWl
0xd8AzNzG1jzXSjsxOrH8PWMGlxgwaEH1YJ0Iu8Uk7e8RxJjWIUxCxWr7vRd0XsT
gOJvGXZwDwWsGOvltyba6NQBTyQ1rivSj6SuPRsHGOTpMfkFP0nlwJYP56Mu5Lbs
6n+c3sW/ZOGjUyAsZmH2PaB9a1EAAGAqsJUzURfv/QVKAjhcz7bDop3w0U/UwZQg
CPk6VG8sN1yrNoggTjrMu8YNSQAaFrHMSy9Q7nEv45C+wWXQm2w5Rp7KrV4RFuhP
imi4rU8mrKc+oe/x9Tvdp0lAj8b+w708Ap3gvMrEuEaK2IpNEKVBsXmt64q2DRt2
5efw2y7/chm5cee4ENfYqpv5aIuxc1YvG3kNkd8FYOXdvOm7CBp1GUE4u7PyN/jJ
3U/KgUQ27+h2OXj7wgQkV26G9SyL9V9bhDH4saHPGOhWGJV67Amxn0H7vcYuGEV1
Rhl9SAAv/fYSieepnr9Ow/M0e/vXWFR68L9Z7IF5RRuiHU2wW5iK06Tih8alHBaS
lPNOUCM0xUZoBximANDgHMH0P+lkhbYNVlKR9MtCW7gW09vC5et1sXZr4aJDz8Nw
OsRdK5Qe5zcDYHlMy5BUUNhLIz6Kk2sRrN+uu+HZpfP03M8tAEL2sUqoOMX3VnAf
wKHB6tMoGhYrZFaIhagVTH5vSNepAPjS6QnWAHrqmmNSKY6yEnaysJmo9aYXuDSD
Tu9Z161rN5KMn654XHqgwZPnLNHwWqbSUXuZCkQtANqxlT6fxgx4rYQvIaJpn/zM
bjdMMy6L9swZ0njiolZnuSedNZzlz0HRk02WzTnYNPoeGnbNAJ5c9xb4+vShvPwT
PFJxBbUSQhjvZ5b46hm/PeqaUGH5QqLr2l6xjacJRIGXmDU7GLHL7fyriTUyOxLh
tq63XqTQuyk6k0i5GxUsiL6ImOVTisTFBsSlfWmgrk3X8uGOikD7SrYLffISPK9M
dy5aK6/B3RtnClT0L3hIJahdkYQD39cZN1vTDeZF8qFOwCU7xyTGNkqj9FoFfyVk
CKTlvxP2RFJMoIGNdYEVNe6HMKV3Dihj6tBPE+QWF3yTByj7MSZ6Z8tgEQvpsF4r
w1lTwbkr6AZJaaxlB7w9LX+3ZtP6aQeHlKzOcpVJoDK3c6R/q+a5TllFsP6FkGMi
GY9iBbZA5XxCiNea4m7JSebVHtEvGxsndafpqdaeoLHcT1CnlKPsueLXIAKvD6+h
AwJeMk9O3fNQBbG4c99V+2tu+uVz/bApmQhe/qjCzciR0gb6s37MJYjMOjzgdV3O
9+D5gEk5pfB6IYaGiFSn0Pf/PlS00OGKslXqUX9NjWACyI/NByOCjO5oWS/or8Th
Pvr1r8COGmpPdke9ylqYnpqjx2prqtYgptPHiwQ2geIq46oJFOymtevBXRu2KC33
qNX581bFJ9HVaLuDnSqJfywCM4qo2lk8oZuMGQi79AW+8geqomLGnaHpQXaQkxbH
X++yud3ifQkRH96QcDC16gSlhXJxrHMTU+/qrwtYascKr8lHyOtOuKa7f7YgDYXx
3boir0HPA27UewaH7ZIET6NcQcWQ0zdwvZUcbNNYz9vxFCYXo8c5Bkm8ip7Q4LPW
D89mzktUrAqjzAJMpcp1GOgAWgk9fn8/l690yHXT3v/5dccLC/CNGA0QfmPN7sZt
Hinr5BW0B2YyyFx3PtPHPGNSyw2JF2FO5Y1GPgfkGB5agQL5w1MfS8tJGXMUfLtA
n/ytmMGO1mhjSuVAKNPOQZsH1gjG38RA0Qq3MxHAkyqSn34TWA0ZehpqIed1j9wp
zsclCVd7Uf0xP1yKoDM+k6uBwVzWQNMngC0dBAtVceVDsI9R7VEBDI6rZfXkzrSS
AUqRZBTirxj17wJ6CXtdemncXTHMXpKp9uQTBoLsGcQiBbZBgSMqPjHMgv+Tl1gn
h7rlWg5hA+750PMXqNf4YJouvk7gSIN2O54/crvOvkdr3TKbl73FxisRd4XLLLHF
Gaau2tXGdeRLvlziLSzLb0LtOmLIW01QJDU02g79QKLzU/kz4ftAn99gEe2woPMK
utLAyhDo2zhydZgZHX98k6FLzC79SEo/bc64s8C/MxdVHmMhj/cR0atYWEKxhGtJ
hrajUphb6cO/Tbwcj/crCpR/AjEtntm8oWXdL5NcnoKtdzgaXgZWEiheG6w+3DsQ
yqKpzpWy9T1uOWzg3CBmCykOfHgxw8QQ8dKTGzTKNImXGR/0rf89GKkvQ04nJOL/
X+UjTXjVFFj+sspLKDm7rNYdrBKx4+YVx2yutnclZyubMUJUHBopSbQyuUrNriJ9
B66sn0eDhoDCF+MpXv3lGKxyU/EFFgunboLdnF8bfzlbhXjOpxVjYn0h/RUY+1vv
jUN6wBR55OYbkZQfhPSCm0z7wcTel6Rcs0rHh9ntPYrmm+CW+udhJu76jtRCb0Zn
MWpE2OesgIpTWUpyX0hJlvB9RmUmN5oxS9+TzXLeOelQGkctXewVNJHZk18HHXSH
HD7hmm1z9c/9HQsm2SYZLRLC6j6aYjhgwADyHLZMw+iNBdjdcdTGql04Qdt08XK7
kUbYYVSfbUiEr67bWNWCBbMPRWnwthGp8OwCMfaE3SeyGeHqO7Yd0FIGSQG2Ts57
VS8A9qC+wMCaOPHu5KrVyWHbHPp2DLqp3i+w6a8A1oo6UlQLnklvx3hOjWlCtfiI
WkEJ6peMqVxm+Ny1SughvAGc23XM+dcnZC9nPls9q8dMD+9I+9P5Tu+QXR3b0Cn6
zNIc5DZk3hFfuJiywDvdXlZlVspDKiA5HhLcoRzHt4tZKjsEHUjJ9WpSfFS0kjHA
ucmHdHATkU4HszZbvr9zQp7UEPD0B7HQj5NCMns+5WJIxVC2ZnEzfXP0RGWWdzDp
UfRAIj7DJFXLhLccRJ1Ii9LWF2armqOnqM4PMJdih591CFboGRIwJ2DUaHvuHTUR
LWrIOtENRxk+XJx1tW3OtD1bt6OB9sy9G80jI934F8v6wm2I87sQqhuB8YVaoBYn
1sWmI1tftTliVjMuVNUhW48uz2uM1qLXtn0Yak4JST+sfrWHSU2EUqU0J6yPVc0y
9YHvWZkXDqEkF3soF8t0eoTE+ZUZqIzdMPhlI7MxosrgoZGNk/AaDn5EPdYcA0Ua
g2Gc9in2PrFFricbW9Ey4vWX0StC2lu7n1YVHq1i13haQxoYSeic9jWvoAQQzYGE
H2ZZKFEpxiDRrumGYO1TSfL4qiAPBgbgU+1yUAxjU1HtLjI4DjLZsEI0Vr3ejHFv
oJeh7VyJsYXaeRrfSp+vnrbT75+uSG8FUjaIfuncB7gT0w+rtQuS0y1APnFjrEXH
odxQkmfd1hVAaFHS0wKQvgRdnlqsopWhn2B7Smj26yUWwF5veN3vc1+SnRKUeqQK
Gpm4BX9phNQUQa1WpWbBUs+uaVspEnkeN5UsE86L/8VFEErHP7hlpF3MfHdWZFw8
/78fygUp+4DWoltItblK8n58gXNcoM2wrr3VsKBrWZbTqQCP/bzLcjhqQVbZDdM2
6xr8oBn/ziTG6L86W63E8WDB4fzqL4I0SI7cZi5ly1DMnRiSYEnfjBEmSCvQgzyO
+buhlMcIfUK1T38c3eZ7W7oe4nEdeo1wRkpdN0HYxXY7UTxpdWupiszCpR9+8Hzu
u1mlQjCKOokavzaZYYAS1zIIq6Mj5b7Pd+NM3LypayQHDrvz6+iWRAFMY/SNkoQH
qS8qlmy5EVBs6P1WUhqVl2B3jKleX+W5xoawl8jws0bvi9YoxTU+buCwcuH86CjO
4aN/KGMRDhSPWDKHNCSKvANRxqD+nyphaHG/lAmcTzYF+d90VhzI9QaKpI+Y+SxT
eUgHe6fYJulTtWkjsYGONcZ6QsTRVDSFMqSCq81YHrjGC9Lu2AOXMfbIURNnWsHB
CWM0g+DGRud+81WyAzVKlrguqMlerDsKWY1eit/UbNRVDglPgwsSTNIIytSL14HL
B8PHD9yB1dmjZ6oXH2ds6UqhLa+yKiVecHelbs+B612drefVpT3iNUPT0jsmjT3K
hUEeBC387nmQUYa0uJlC5xl/yXmZy05H4c2GzbEhf1obq8KMUV0Yytk1EOU5Zbz+
TH6OtHpf/rHXHig5vUPIJBym5zMEHs4SHBFYgOuA5/SZkJquH52LVVkImqYHo5LV
WU2siFQOOygHyVSvEdCad/ViQQ+bUKX/Pf6TvRr3vjF2HqDAOf67a+8FxmXeucT6
b795/dSTAPNJBmvltta6H8bd80+3OCANRL76HoTGoEej6pk5Tb1tAWdrwSJf6/NP
JsWuJkTUIFrJpvyo1YxEbP4IVAWJVf29EYRYV0+19AW8g0d8UlJxyj0h0p8rcrGz
V/GLIJlpn9dXjwEAYcszkHXiBjvlZvAWQZB6PZVTZr2c6xL+BFlpPSFuFQ+xx62P
KgyYWloavtl5kb/2bHevQQFamiDen7niXjKplq3R2tEVU1LenQvyeIyFmEDdpSUo
gh2wmC6Fg8HsmClIGTX4Fs/dAW5kKYkjMhLbqf4MZqPoFIJfzX1rmRGcFbz9ZAYG
hqnt+TyFHxu62Jx+kr8j3c+P5hB72OAK6Ngzfv25h27Drt/ndXqvLsK+Angc04Ih
oDVYqjgYqyD8TRwlKTrIpS2BbGQ+Az7IjvLz8N7v4kMkt3lTuzBOxPcDEPAWZeEi
E6ke9vVuZvRi/WoUjg79HF7s4W4ARhrnBvN4Gpmbe6joKINE1rHYm5TLmFaK+3Jz
o3tQBN0BH6k847xVU8JbIw9JufFh8YAmMmwAzWI++6+bJy02kvmq1+qFouqaz496
8gBU9KtlHEy6qo8A4spnaGX15/7JyhfDeksg7HszpCGYhbCWp3l2NWbEzcASC2KO
+89r+SGPo/hYxRIGJucmJNsughL6jgyDCiyi2VlS8KFM0CX+8AoRQLfbTcpD1uJe
uUhR9a61pJ8bENf4tIxCcQNuOPHR1gR1KnR77EDUZW7chI85S0qwEeMvGDc7oBTf
C0+iIwEzway5JdGTDH3kk37lEQwSTYdDIFW3mZQKRCa3/Hvi305LCmmtp88ry/UL
cprdjQvYncdt3ON+qXRdbbHNROmlHkvvmQ0u0D1TJxjUmHKab5oMMA5cfkI/xePc
PQcLM+2IUKmFcbJGvdTTYuVtaxc0nu4Dv9JfXmzeiJuZGMf/YgFmFEydWm7Up4IC
oJQqB6E4hsJqagGpKLIcBjguFDQ8VvwkzMm+V12sG1r2m/FIogN+Fgy+d8g944F0
THmt3Pe6fxPToM92nGSX3Gh0iIW6281U+9lAnDequ4SWHw3tUTvNnF3tNHbAYV8V
moHcqWMIUV5EQH6mc5VuDQitCzaznXfmPw5dxPszlAsb/Jt61f22ftwl0U1ja3QD
UFkPhBZZoBmF+gI66DpS+FUWSZ+6W0/jOHXzUZ9irMbUn92HiUsOlhZWRKsHKOKd
s6pGGKS3huwd47ObURmwssR2M3WML7at+LoiHFhWAaf2upsu/6R2k9VozV6MRLF5
swHucDYcE4GzzyX7mj6sQERZRbqpimTZETP8+giA/yFDS1NRyXA1eVKH8uyOsjHZ
UGtAGw3Ic6Dtj76HrGjd/5SWvUWE+EFaC2Xri2o5H0/tqk71Fqhlgbl65l+v+/b2
9oRff1a45es/gq7Lr/GQ0DJLlSWM+4LJD1sYI531+TixsD2GpIW70frCvgqOHwfa
uObMShv4VskdbQu22n6/9l7va/Y7gkwqWw5aOq7vjCm23VmDN8XLW5YG1oNg9lJu
ZG/4qMlF+Z3bNqE9RvNNZod369pxPpgASdbfXGhWzk07616+iuNwFHyaFubB2+Rh
+8tp8qWW+EYefkieqSdX1ZVd19fBM+OV1421CsKAgJm1FPdCOhzZa9k2dGDlvhBl
NekrSGtQfQsKpgb5XPxm1DesJ1q2tzFXitRrOlVbhpGmZ+pN3aewV9InVdaNQy7H
U8EKa9vEF8IWfKayPHU0hmkn/6oD8yWs8miR4C2+8pHDSVGMhpwphiYVtk1WnqDR
RjFR7a8oTKsRpY3FIDr1am/Vyqc4GxMgNRWvVDvOuiCcz5VVui6LNOCxYt4foH+1
WOjQUvC+deTL2lJMyuc7SpNdaWU+VDCzrKFxNYJVsD1W1fi1nNezcUP1CyktwrsN
TYkce5PoKkvFPJ4DirNjCA5qemzvt3ea51JESynXHm/efKoOMBH6tP1vyjiQZ2iK
5+aDHXDX6isXRMhTiAZzMyDowuA6FpRs7ZFHt3L5KXqT2nPR2NePGbHBXdTHoyOL
w7fVfUle60XR8FgtFhFCRkk3yakZd4AQ8fg4/s/OyEyJD1TuCAJag5MyVQaRtQwe
RVq9XxygGXSJTvJ0ubhz+tYaZCRwvjYGe3tI9YD/RgQg8xPC7Q6mNwjBnv7c2Raz
rq00+fW/5VZeIi/szaCdi7li4y9g1AknlrDhU+FqMdOSVvmUUEefxwlr0bgr65Sp
mlePpXRFX/CD3MCqjHe0Cnroe2s3+TJyZbA1N7PwBuooqiJQox0PN9giz44Hdprz
/lpwKK4CQ9dsw4/Dpl3UwsMtFsrmWF76sBeZhi/cRoKxapewPCqRbBMeXI0mmFE9
8cEoTL1ZZ5g8lDvaMKR1PvWel4nTowIyTRNhDhHlPrLSL+/FpxAZQzVhW9xRftGn
RLc8+hgmO2iUYRrg1oemglRmuMcVE3+I4sZV/lqtlTirR18LKDeM+xBGdAOfw1iR
Yw8NvEGbEgZyeJ69RbCsgpItU16khGlz28hGwx317Eg0ZeG+Kt6KZ2+mQFzaXuLo
edE308cLmb0HMqIOxVbj26XII2EsLKfwmhgRB0TVj2v8PMrUgBYwyoheFugehv2J
TsejvW9hYAjz+NElGA38RZLVHv1WEKRR9YZ0UNADZ2YjarqXAFNza2cOeeEYl9ea
fM++aLxRr5JOGy9jJfUeSDUubBgrcqkqgRa+VxZLA5tzFnZ5Q/jdc4GuJDFkhjRa
q4OdhOSMH+/80yTl8CW2AeqmwhvDchRnc5JZEbB+OkjMghn2fGkj6xmKivuDHNHI
8NfLnGz97gaLvQgyB4lpUhaFLnNch66FEEVmChwmq1p4vd0hXAmPiTkOw3BUB7NC
0vMdS6hhDyLOh88cXN/fEdJMtojMc+l5813j0n+dY+5hBqosOLJjounoCH1TZYH+
0o0acYwJy0RxTxr/H+bEJoDbsky3T13WvBFI14TyLgS1u4s4qWQOaBiM3jZeSjGv
xWdzn6A0J7t4rqHUAUsSsaUgWmjo5eiaUAi9sCMy9/3kiMG3OJu/LLX8ykWf9Fvt
klQlxu8qva6rzkY7za+xbBTi4l4EOamSxcR6hBDuCndQEnUpxC2CaDL5xYDbQ8Mh
+o4UndFznzmsmxng7h0gfWdO1ci1eI8Ey35pxciNIeHhHQ3S6gzF6gQznzo9ls8z
08dxIoUQ6UcA3qbkHRQBpWvk41bw7la7OM0ubvs7C4UKufXs8+HxzzEgdFEHtU9h
NEwzJwjUCcin9fkoyVLt2wGVYb/+XjyQkBI0M3NyKkzyu6fZYXzjZZrxAjKihq5H
rrgqDKv3f7DdfhxLaqmutOT0HbgXQfbr0XNkSVWse5vSa1UMKkYhGsBWhaSsI3yh
DE4h4N4q2uwtsaHbWOznfTxoMHdrdXsKRGBqWLdiGQonTIVRCpvBsFj3gFjnsSMq
RJ/zRmjouNHdzXh00yvsPwtUxq/zAhaqfvCDpBqxFbkThryz2iU2muQnZ7nP19tc
mkvADnQC1oNRWMtXgfAiacVHJz6fDgsaKPKSsXNrWNEVHvCaSLxGgnDoiBDyQyG0
2CcvKz8kGunIY8FVS0J6t4SxqDrJHYiMNFFebWSiPonJb3+76mdv68G38udZ3kEe
XRXZzKWz/HKOSZLvRCkgQMofdzxsuwhQ5PVVBTsZyLhXbOlWavv1D2qcfzWHHS3k
ACPdewulaZLv2A8spo7fZES4OFGiL6HBoG8F93ZUpgzbKuYLlLTRVCHUsfDVnri5
n6Xt9oDO16pIHunJ6iveZX11uOvJKxqVczTg1P0N7jD+sfgckZ/DG+zXylSH+ZXM
BMwdi1ytYeYPnuquJSvgz92QDFoncelXj9/prOs+BzFUhn0bEzMonCqlmIY58T/N
eQk/253DrmSCk708pj0c2Om1rR+AGSrKZhfuaruR9ZjX+7T3rShqVu0OKfaomvO1
ihjJP906njT731pwHJXi182A454Ipv/pKaF60jhkyNyev9Sxih95oOXdYN0DT2vi
7NUOrWSxF9dqovWiVfyUGGDtj9OvrfgTf7OxrOXx7xkJEEhij6N7j39S/RVMGj5b
nB3GVXCXInpiwjvN/YeUy9f1L6VepEhQs4WCnyGQ4McuinTNKmGOFp0UskNBb2QE
lQEJ1VuV9EWIk0e367UplfvNqAXR6fcPgV/uQkuZQW9V5m0+RpgBr5Hp653UZpfG
kLtn8Kx48g89IUZ3Mvts5Ss8EHeFeENCiZcXyc+8SoE9x6+UshoH0AaQdE646Txr
zfPvo4FmxQWK8mhPxYDwo/TdxofY+x/K3hcDviiJc2MRX8T9xAi2jc/mgVYlJQ0c
VszkBypL80rJ+bytBX1UTPBEvc0IYxJQ5W+RdAkdzVBBFn8SYG6n7aZCC5DbD6MZ
MfeAAzvLiwMhfhzUeZvftIwkaemPH5rDYWkIwQuj6jbuS4fp/AOSShuQlZ+EdOl1
qrNh+ilgX5Gkndz6LZaaPqZOZlo5zqfWjFcWkRs30K3ExifGIIKKqFuAvpBHqO7w
3U+ZrLbTNKUtNGJ3D1RaAAO2a2cqF8YTH4FdmunOnLEbnRBNrgRQj5Ocojx4OFlb
EpeSlc0hlbs/4S44pxbHyV4c6SlGuFxfOAn0fV1ZD1jv7PH1zO8soAi8BMxkDDNk
8dAIMo24Qg74CPPEOFlhFLRb6EbbVgqd9ulEVSJRip3mDd4zpOQI53/Yha+4LjbG
39EfnsibLX6iz9ug4xQulV1J5/Qpy4sLDwM940ATV4JuNLDb/aDMte/FmaRDtKTT
uScU3Zc3XXaQL6t/laO81kXjNue9Z8vfAMTWLK2YHrDQw+aNNyyBk6yrZemSkdgM
2xuUX1nqxn+/IY1USnJbNqrzx6/m9oAgSfXeRFN/kbWVu5dQDSMvkPa4b1FtBRIo
QL9T0SjUaEI8s/rR0iG0XmywbfkL8eOjAkaMf9k84CTfLrwhxRxUfP59PSr0MAMD
SkN90SSxiv5Yn52VqLXvI7S3tLsrJ4B7EDlhJ8E78bR9G53/tD9M7784sUJj3JkZ
p598/Vd6u26oVjkkdwutbveAFMkk8A/0hQoLGow/vUG/DmVn4VTcw8EemYuUIKDQ
zk2FYL85Rxyidn8iSWx5kkIvOcYJ1isoqKCf08C0JTWTNsCzEwpntIpRfIKs0ZaJ
pF0YCdZmQm439smI6NbXbiqrdn4Dhqo8QMvI4Epkilrv/XK9aiIfkdfyv9+TctcD
5GdWpIFTVtI3d+0k1PWnT9MlHb/3oNKoErHVrcpf3hGZBXuHxrIwW+lw/XIBXr+U
jtujis3OXXnzAtXFwmrTVcuWqwLtQBDxSxShie1r6afc2pPFqVukitLhbu1wFKXO
lSfvB/ZPcWj5IYNVLgGGX3u6bk3WXo9DoxqKSwaXIZ4g9/oWTW4e0Qw11OMUO/F+
AlW9fVEnX9MmtsoZa7njHR/IdRrUPnzTiqTnuMudvpus4HYb+TYyLWhoLN1O0y67
O7NeIEKptBSXn/yQzKYmrecsL/6ggg1h5s4DP2zHokmtkFpCVc/VpTVBMXk5cIQK
IWZTm3xz/xCrhWtQKkCbfneaU8TtEE5vHcEhmSBDxJdpK96ao7+tIFDAymTNYJQG
ep8J4eEQnqmoEJ2qrmw5jl7v1lO7r2ia7KM4QS9U4pllH2XLSyQUaafZfXfzKexS
h4WnnUHAthv/HEDLJxvvxNyxgSNfVZU3h2dU+lugU92wegooVoo3LgHSMTvB2TQo
7UD5g14rIftAoBUFYBFqqNrpH+l3jf1bSGtcMRQiBbpO0XYxRZx2pliCRWiL5ABW
wO6C86Me3j+2zwZsWt5nhJ/L92TJAPi1q/BSVKVTbykVm6zUo7y5NIq+0WzK+rZT
K0bCQebX9kWz08X742n9tRftupI6liRovaZFNxpLe+mfxWcDHzDUmShiNgNXsSXp
8bkE5XlVf6+Zg1FQQgvUKwgQbSLxrTVU/iCoTVc/+6VB64lPcJ4UlKBUcCLzMswx
Y9xner4UgSYAlaEk4SjXl9zQmUCJWjLhcir8N2nyzXxnFvjrJ+lGngaxKWKLNbEo
eBB3IjulJFokdfavk5q8MrHbdcKeSl0qasDu6Mr4vDkRYi+icoGskF9Of8syz9TD
Mjw8urS9v1C8ai017f25BywC+CgQYCN5oQNZoBVWg9VMeFwavxG4E6vDaOoJacsq
nyUYUXcfBUqBcK525Su07Dxg57l+SbhoaTLewv/vPY46FMfLtuEyw/PnvFahlQlq
GsECiRbauxv8bMzBeEMY7M0bBPB8vdW1o6ufhayeYQdtK4C1eSdCsUbOmeJsUapW
SVjx+wnoFILjuf38uXeEVxdl1ZW39TnN3t9hSVuAsz3KeRees8jQo/GEtP2eJkS9
TulT11OsHNtuv6tckLJB1V/FRmM9jSFhL4EbhBY9EqwLi0c9dnSYoZkfOpxJP2SU
/A0oPMk38t2o4b75a66NiaPBR+y8X3OA5RJpAqwwycZtCcN2P+GRDktPZmMPhRw6
HxPqij6u8sZIb5Hn8FLtW5BWxOts9J2UuRX8Dcg/USRCN9nz4f+otuJlBkO6lZLd
YV0ErYTpmLqHiPeG7uk+Sr8y3azpKkBKlQvo8Hhs6HAc2IF5JqzE02Jdsdy8SWRt
xabzMCCrEXcGN0S0Xhdda+1s6D47TuZPk9dSoMC2R7wGx/pTrahDxwB/pDCtJJwi
nOyrtWWF8y9h0gUr56+iBj+CaRwbpiW+lUc9VDTQ+aO5ijnWE3Cu0IKY4Mgsd49u
Yp96aNn7N1Mc5GyUB/PO/YlGjgzr96H511ahSHup45Mn+LkVKPuWh3g8RCIfbVl9
P5RlperuRXA7umz9q+nheUBvl8iNzN7FMFfDwRIp00CNcBp2mLk8YcQuH8OOagGk
dn0mCYJnMo7FYbtjANHZzrdSqaJr2b0esyffGjp3muJTE18aa8NiL+Fcdgwo/pZx
2/cm4ZAGzSa1z/T+rGLacJAXf0obzm3T1Th/pNjBSOdknc1wwShIz/HPSHZFKW57
US/A3u0SF4nYq+GWmU21PBy4S/4rUb6RIV3s+cyt5d3lGi7U3vwFvz21Ju6vFRPw
bELSiVq/nS0TLgbNlqfj0y7/n1L5S++ejzzcFHDzxFEKWiP7va1cAGLWb3o5po/3
zBhGDr0Lsp0CsaORj3kWbPslaLAx298k1kEcif1K8Kl7XIVg0ixtp26nHbP69lxc
JFhFNA8wdrAIREg2aHtPTpCgl21du8xMLp+fAVTSHZ6+BUjF8vfSUGDHOUYMt4ff
wXB1iTRR6zDCvGzUh9pWbcijlBGMu77IS+M+md3UaivpuIt2NnKHsg6zTeZ6+A8X
lZ5bdgptcP9SVm8pi77j7K37303Fcvkr4wHGi6CCDoSmYabj4kjLaN08Hgu8DtG8
bzgYSrMZvx4J4l0pJ0GVA2cuIYtrwiJxJjZafuLl5qcdhdimwE9/TLpH4g6uUEV5
2FJwf7/PBkiO49uiy+7fIXHsm8rWlrJVjhudoSVEGChZFfCjt3udbLWzja5VhP8+
Y5Bt+HW+RICKSCGLkycAscVZrGOP+rbmbsCHxgxoR9cNLnis5t+eMTd29bs+SrLi
QPyjmkpPo76u8thLC3tDyAs8ThOb8m83LRPGQuIfGr3e4trZhU2skYeSdJ8kjBqf
iDwGcnOI1GOe5gqlE6pb0MWgFULJPt0AWxzl0x8qy+zbgXbI2yYyj52luAth6Awl
oPbq65kDRC94yYimc3KxCHtZXM8gqTR0Nf4WiFzrcQ2sar3kR1uzpmPE6Bkl0KS3
J1E8wD9nUU2TxM0t0W4s9RUVrKcPN4RYonR54yKoEkdo+9TpWrokk0uud46s5p7T
C9ngEZuYCZznUctjkDJvSyegrSPg5inrakS/AuROOtZClv8hbuCQjtgxym/4AR8T
YSctIrnTceNHvhf+isfvx13h4yE8K0+MaHWVTaJs1hFdWFoE1xF0+d9WS4fynIuF
lazUsoTxXnRwsuc7o9WsvQLShchrAwFGxWiNvP4XG6DsIzCYnxxR2JmuTgMt7u9i
I2ePaBBFtjDV5Hxe9rlVvYMAaDyOkomVdgXFqIJGLRual4QKbhjp227NeEPZzqVb
NpTRLRW44A2DB831o17xWItYcT/8kX4CbtmeL7v/SWIj4n5qzmWSgCytBs8t/Ep5
LJ2+4SXLCw7wrRwVQww53ljfrLNRVhNU/3CGvPCzIc+Z3XZaPCQNsxIhW+R86d6M
tnQA8QqIpvNGFIntNEOzkIhUD3lt6r/SBSWMqHH71XTeylOugvvYbhl29a6LBDV7
OMPKgILL+gzwLTzuL2QpLvf1YdIdkBgxwdVyr5/R6gaApbR1ZYpnbNxn9u8M/b5L
+aIKsHjS2iueR00KA8iEDsr3yiQb2IjD0NN+HQbKon050/nIPzlkzW8mVuJ1Fa8T
V/JQHYfYONr0YH6tc7Y74UZ1aeoN737MG37BzASzHtaL17JcDPObPU3ZTVwsiObd
vqaa5N05GxAxd51LlEAtXWNz4hyf5X8JMZF0jyqDvCNlkXGEyXpaEefrvZr0a0Af
2IOA5m9Z0JQoiMlpHQhVfP42+m8Qw8XJxEXcZDb1+s7TivgphAW24FAPyiOJ5QU2
LXq963VUdX7z7DU10sKqaKrrzkn95hbmORjQoSsanS7/mB8Gt4C8ajeKsP0RKmKJ
J9evpph78j1DK0OInzO9+GrUbErguzeOEhBbIwIcSoha2EGdvwrO7Hd8Hh3kglrt
zae7A0AR/p/mxNYXXYn0F7JMYbTVN7W1UeYnbzszKtl+v86yXZKlwqq/+sX57SdU
PHUhtZyMB4pJ0BPnwd7ob8NE4P/Nw+u2UbIO+eANadgJqbld/Z7XUOcr1yB1ajpm
D8ZpjVIuz4z6aChbrz/XkeyISzZ+nm8rLIagSHt0OVy0/Sifj0W0hpajs7fi0RFl
nqE+Lv6cZv/nsvsrJ9M7pqJ4HNDDSjyMuW4CQdTI+RARjPzrd/JgWIJtlNAy3ZrM
KlVwn0YzG4rVYaIMrIlZjWXE1HHQ9GC56+odtGTYZHXvrcyJyf312eLpdIGZ7p6L
9BxLq4emq8b63PN1J3b6mkoxpf1UcTEZNImCD1eYH2p3HmPvta6a9rarnHQZzkmP
1af0j8e3KZHpQOPql19WdH5V60luJpLOvIkBJLgGQHdfVdz4OR9dEnZD+8sP3CrX
21BCoLfx20uAda7wnacauogIEF/LzulD7/yDj9FI9gsP6tYFHeXksDhmzT5PO/JB
7k0fph+ma4q48hZFJHLGEwOeHfCxfPUyI4lGrI3g5RC10NOfVf6EmGPRaqpMGbud
RifTnbvpnwhg0GjpauZilh7liPOou67qLrAhQa/V2dYvPYFnLMTKnyVEwIx/E2T7
j4ucmbR+Lb/B6U9fDeLZZ+CK7vJ39516DNr2SsK/JbrBo840bBlyWeOBzXYtSxT3
dQKu89iiN6nZDOdACEceZRzp+7WOztD49OlrQxu/MpuuEDcHZNN1K2w2/H+Rskl3
VMBqw225MVapL/Pk8leFAJjqit16hjD0TQbxz0SioYn8nZM2CEOLsMUXE7cN+w8l
Mk73RQSJdEBpLUEUW4VSnw1FDFPUtz6CYDqz4P2Smjsvow8ufCHPbdIbWPB2V2Hc
gnFgTbLFEBYfo9dY/KjCnpsjBMpM/tXEcSvLzY6RgsCCJjboT0Hfq1ZyA1EaF5rO
V+QrwFf/zWhxCW2WOXiHiPeFvcOeIWIdsUycSKedVOD2R5K0kdNrE1h5pdSd5eeH
braqdGOlpzDMlMiSXs9O9KfQ1r0JWjPhjTq/R19HhSIfGD0SHQuTZgZwUk1v+zRR
cZhc8P82+8Ufi6UHHvUCneQ9dhe7vNmYz1N35FaarnM6/NEl/CJTkmni2FWP4urG
9U4ustSpqY+4XQ4rw1m2ix27sFC13bLulT4+1aGEUBf7aB/B/kTKNwUM+w+udnnS
eceNldHpbFP8WWjStrp9lPCSSAgufgEiOC+SmMx19r9BMqrM4uhQ+2ss1vEwnsa7
Iw0TnSh5ss4eiKusi7Sj5HaCPhm9caL41YkjOm4ktANFIsVFd+mV8PMSXd5VsQml
LRUmfGNx/mqV0V9DZrEFUqOkkzUj7mK4qMOuKiR/UjC0VRGWWdps4Tmh3V5EIwh5
6s2aBHY4EuCYeiTsn4JLsQ9ghZYaZvFih7Ejd521BxWd4itGAia72DrGM4236cts
SsTsTjv1WBY6iI0Sl9wnVxWRXRbQyl4hL8o0ktIyeM4/QybdbT83+YJ7mzLyqdvw
01BsV3E+5zJ/PIFmgzHt43+EMNrP+MaGrq5sfBwwpo1jZpFnwAKNSzd0kz3tWrze
qP/bQCqtlfmX9xhF+fwrcBqrdgTny2qNAim7HJNbFbNbqHiIlQSlxyVW8XKUJlG6
TkvU9RDrmPZeK43nK7h2DUMldnQmCJ95pgdr0mbyzXOxsPPgUvGFeOs59uhCE7DC
2Li/WO/aihsg/AMSq0bOq6l8CMZMSAd+aQDMW8XQe/ak/0kwE1NRz6ZYBUbditQg
IR1SxfO9ArLAHdtG/9XwfBcxazO+F/uC6jHSXBqrE/jl9N+eDnMKYInAfeHKCyyy
w5MMgIaH9UnaS6K6uB9XchRW3WAKpILI/fFTMXFdpxAVxU42Lt+SWqmKjpqIUvwC
X5rfFi3bNog6oOI5mAo7ChH9R0lnix9v7WqKl7cczRe8/B4fYFsqpJ5DC60dtHL0
V8Jyl+DLSpFpq5Nwy1s/46xWYipx6Exi9TznUQX8SJlxNifpwikE4rNNe9CRVYOV
ZHJINN06o1bXPb0c8PgiVKJo4Jn4N+LDOa60ovJnSNm9gHz2tdL39HW8g9EeAhUT
6OHRQn/GSSxTFxcatnL6LNdM3mp1Y9cJL56NhhH69lG123ZeCYsmHDC3V+8SIIpY
a6AMoDymcOXc8ay0QyHr9QiR/cuOb5nA8NQ4Q4i2xgVYBTm76dw1bxzSAC7VukzT
yKiuem8AkLSljX6Pb/4h4Pw5SpUUST9vs8x/OgOAnImXH4JytI5gVdMlnh+6gz6r
RxMdV4etGEz7RkyXufN318II+ynzy7XsuSjAGFEUH+xP7j0Yot2RV0F6V50APiPa
0L2aRghkWKHbDnkdZsmMtXcKH8OjlKLq5SPDKofvHRlA9PnbmIc4/frRaZuUeBkc
gocSYDseKloLvBVrVubm0rfzG94UWtKd2JOWXRbBrCk5eJWXqiGFm+1yJesMbryj
OrpJrgD78nR1hUUEPhwFhUO3v/o6QqB7cwvE2guriZ/gH8BbSXGXUwC1rFVDMFyc
8cBNIjWY4kzlbldxADwCoETd5w1DfwrU4QvEffGUDwtSQpclXDEWGjmoo8JUJArW
To5m4/I28f7l4pMbOF7wx8qpfx6av8ivKG9hWyuYnk4yxD/im5RpHfYyrrc1kw/w
+5GZvEYYZM6PeJQ3KrXsbgTjq6peXPiE+SngJx1TmSxmClyWNGO+6XuauS6kLgZD
g7/Z9lAg/SoDsgnf9zhCp0BH9ewQfDbnMxhKpC0Sp2ZfG9Ec0JpUd5JOyQ3OShF8
h+lnInQtirW9Nh3uh13+TDtdumi08zKyWsWad4deqIcT3krTcvk5qU434N8dMkRG
B4BpgYnRiVciq8lZVkyKQM+t3+dY6f0gmOltJrhE2frKOzjj1VTbJHaj4I5DfiSj
2vIV7tNQcL9Qo+o8v8z4mZGO8TkKgXyzl3LrW1i7oulThTNB3V4AcJlMxwTDHHlt
QXfdhWE4yty7qro/AnJx6xHzJb5byXr7K9/9f9E7dMdmJeqs8eawzzOQTn38pVgj
hEuuUzS8omiIPxuPJugAxRFbJBWye0R8CoTFI9GqWqWdC1z2f7e1Lh92fI7u8cEJ
7nVaNf5/17eUxWqpK8YqldEmD5m/uD/XxulSDTwSRWkgWU0LfHQKqq7QfVK4RkyK
lzbiO3e1rKivNz1F/bDOme0bNUbrM+GwWsB2Jcx5BKEcLkMqQ7alx7THyc4rgiJZ
g5bZ5xiR/G0nv2BZNEOrO4rAh0DC4FqCt7MqAO6cQaUU+4OisDuRgx4BZXcoogCz
vetrL8S5jQ0e0iHrWhx1Ei4DaZsyev1eQhgAM6clonMoJ3kfTpBUUCvf7LXlcgLv
xWbUb5yyU5IpxP7f1IRJrlCFy8urO5liI6qAm4L+NI/5JOM7wkdgwbDpsneT/Ndq
Sxkej2PefDBEnHSsruOk+tIWK3av2rUbqc5y8wlLFWl8BQ6oP91B5Q0t29EQSZfl
7jIEmY9kPrtbxfDfZO4t/7QLNu2oO2ZOXPHXUXpSeyEAYofB4igPTGCY4Od3/ra8
8pd5PSYZHXJPTPiWo7KEcdNKstcFM+lIYhSsEeMp3EDF/VdW+1LA4igFVTFrmwba
CZwxQzyK9rRD0ALdIDCr3X6n5f//n0VjEiKRn2P+uTn0VDHMg/mwXEOujMFfUrBp
hWaEImT2UCtV1TFgpnPxNBth7HfxJc1CvoY/KYctoqeZPnVBDow6bsYCgztPtY0O
lVjLSc1oVqyRilxEgzChU86E46w+bq38CEuK1+diTAIe9ox2ajAMEtYwrwSsBDhg
lAZYV/sIPTLkXHl3es94p+07kJW7Ntws59mYBF5ZkVlnhLY2hfnqyZ/qaDsu3eE7
Q+GMIe21tQZrVwZUpRd+SMW/ZnxZEGPkkB98AK1LIYvxBUsGA0ZwPvgIE3Q9JhqS
9BvGH8mSMk2zXLU83M7Ee7AFe11IEqTfK6h4zxUc3VhnTyt2GApqAEENuRda5cLD
myF73n7uTNzX35MKIbTslG1VDapmBx1h5/+FsJLdWdYqjYBgV4/1MbDdVJ/Cdi+U
jaQl6/u6TcWbvakunI/HU0GWRyCAH7I9+LU2Kc/edYfV3E3cErMKgDanAJ63ALul
NLt298LOSAFg4o0rZ0cuhw8Dtbm1ZSr/Aru6v/cNrePuzVW0Q6drpW1pqyftkvC6
ndGPnm6yX+2kbLJI1UNXApVFDSNrYf7c6tX7IvD7rLM7xWtNWCQtkb1SldGe45+7
cpZENMdDqKxVXewcF/MN1OgRmPfeorEgSKRBCiUmCWqWn6oVHE0gukWWrLsIwEK1
0axMvtRPh35aNP5GRJYqegUhLQyHTWB+pGPBZyx73+pkTz+8U7Culu3ALoLvDQIm
KWYDIlIl9VEMTuZmSFf0aeCDBzQwcGdW8npyGtLyzuzt4DrTR+q7MBrEXWDtD8bU
vPSBywi5OVKdECOk4EXaB8YBhZlrf261C8vkxabEl6JRp1xm1LXvAsSKRX3Ck/2L
otboWKKZb37trutMfHDLvbKR1yWEQKxTe8bWQyBKFIFvJnL4nXqTkXgoFFm+A6KS
k+yD/qtirGa4oIUEDZlKwlPfCVOAFa1bBKEd/FVQHAXqwUDo9G948DnV3iEITCWP
a7xMNox6bjAuonaq5BmK3wB3wmWnFdtA3no1tgdS4bSlkETHu+4m2641QJSfhsJT
qJCeSwsrkh70ZAhNmjHvRDi8yEDP0bEHc6tSuDQoHOWqRQEACM6XCKEijD7VjDgl
SMQnrcmDb0kCrcm1RgLiM/rBBKzu9IsWjwWefkwZOkJtzLyVnE9EUkcKNndezBXa
iCDEI0MOBhBxWKmLY/6hvegSinKWEWxra84fX7kYft+0MnQ9c6t//p0au25rktNs
Swwqy3jF09f6RNGDgYrQBjn3YQueI8O8tGXq7GPQou0BXb5Cer1+XXEsvF9pzu2E
7EksMl5dufttQdyY7fU55H/G8VLZFPbnhSyRUMfCnZ+apBkHrrd1JXrkY85W6FlN
SZA6IzdN0RUaFVVibcBOqq5KKIBYS2WTu9XPnuShp4BMAGasc2SDRoCkK0o4vDTI
AmlQMXZSeKbvDGz2Ulp7o/6D9elhIqla+EtnrHKQLDzLz1WbhLFmm1aIhDuGpVP2
TxpqTaDz+3PtJqzzHvSOWVxuFO7FyfIvqV0p/sQJjY0trrjKxHwsz287D1LYqQnV
QYsIF0QPPWsM27/WqWSQ1tkmTINW05H3/LjOQDjaXSBxtq3SXmoZLWVDJZDU2WnC
gXU/ybI7RHHNyiMOUjn7bXZ6+tUMDaPpDrqbKuNGeGQ7m5rV+yNDF1ZNJJ0pkino
SVkxIb+YA1sSuyrfcaYU2332Shpwf8+TF9patRqrWyGazdvWNVYhhHMe4u20MU4q
X+82XMZDeJu0RfZBWttPCN9uK8g+Q4nRT7o1pUI2BsMZluienyqtUXcvfuNiSiSb
UBG07FBU0vOy7WjasCd4oxhJJj/25fspx13EtXYX+jJcbHYapwSf7ivvI5IYZBoh
S+D9dSzrTla+ggCgV493XoOzJa1g1JqFATXoQPmHSn2yYaTsFrEo4fvPeGY61rPz
CrXRXVs7x1r4AY04QPSIA3GFqeIG8o48UaWTrDF3LT6keH8sz46fK6LUiSODoOiE
nnxjR0g4go+MWEDdCn9EMB+6/eK2Hl4w+L+7pBlpvDvWRva7v+ac/qcB+dCui3h9
nDui/gDtC0oHTbYyW6Cms76cibdVZPPlvlxKjUsGyYfodq+aFiilSM67N/EqPCM8
GEjPfT8zW3aD4jH/jAHzXWV7/85NXWK+NgFwgYhMt0llXzZTi+p0eWqvb8WVNokO
uRR0bEHu+9efgSFk5AxtSxNJjiS5LD7E6cDa2bqRdPYoydgy5CExl9r7KYcIEoQe
YMfOumTlEwgYTsPrWGapY/5r0vVQwfUulxWvSy0MnIS4juNeEdkAPVqbpR9fkNeK
eADux4Fs42wSkqz3e6kZPShVL57b0dLqx7Y1SBThb+3yVZ2oLUzaVifWnsbm9kfk
Vnt/RzsLJIFK8Ffeh9qMHJ6v5IzbNmEn10Pp81uE8F2RveJqD5IM4xobsMM/crWl
o6xDkr0JE8J/XGEYckMuBiSxLkdSnscWqO0vgD+uHuevpbn9bBaKNLGs+EbGfsln
1bJ7y1A+XyHLQpWfqTOapoTkhbA6lwR6g/0Ss2MVERLt3DHqyH+aSLPFIuPqtvhm
qYeb94anacuebvYxdDqcSvnnyk31P3BAHhlydbnj6s96mv2C66wZ3uX2nuqCUkzK
YXRgRxLM84c56+CoMOQggfbcLgbjdAmlIeDsJcpDJ2E2Rd1WCSmC6Z0zcB24HYmk
DD+D5V+8DmjGYigaDNabgfSBGaGJlIrerdse8nPMi4IkkQiLdrWlmc79mdLVc/jW
llbf1Jw/g0baG1zjbBDUIOUvzIlZifNKjbpep3dhUjCapUN/gdBb+J85FzOs1viR
ZNICONKGcX0QCdNp/nVTICe/j+0DwVLhj3Ki4zaeuLpO2v6Th/GSppwJ/E/sqKQv
Moj2ieWmoHqIrckuXUjk8uoN+1MLSc3ttT57Ho5UgyfLCvLBnLhVXF0WwQ5LiVr/
an47VYtd3VlUTpFvD/JRwPmumI8vqOtIVTlVqsegf6roJFCvPzmk0XjAIdKNs3RT
jbAkvisy9JcCt5LYarFlQRTWNYT4FDvkFLe+yIdJFkpLdZmer58R9JsSkerSKlwt
dh3Sd5U6bkFUaOqpyfyGg7YnwsWZsxiuyje2u/hXuNaNU3zSgbAB1ddKS6/biFlF
B13remSj4DgdSLgOMDhXylHAcLvuMiy/aE72el3k7Ar+jmqdMwU5/fK3+rspOsr1
Y6ZLUL+q6h1Q5ePeE+EjIXVZlcmt/ujCK81Yc6R8/hObPuxS1Z7JpMqq97uAJWED
/E/AU1bCdlPsWRFtD/ULzdVtYJSgxOPsYmRiUiVOwAeNdlezUYTT3ryUgF3KjhGA
4JY2VMZVEVUosO+3GhnLkNbBS00MUbGXfe45m5rOikBEsBEYo0ycsaK683NYcigg
/aS2oOntAHAxIWR6x9k8x/dmSyb9FNYxqPun45GP+Ez8qK1prL+3bQuQMM7ai7vO
wE+oO4Suk6jcQgJu19n0JTYSLMl+P9OMH6SRoYOPbGmkBgaatHkpb8rPOtrd8p3g
ri0Zzbqq700sDOIZXd4rzqH4MnY/2SZaFrOULfCUEcrPrmxfR7efbzClkPH4uXHL
cckF/xLI4CaerIi13N4A5UL9OJTPOeLAK29u6gllKdtrGP8acxy0WPcwr3waPzCc
u7zNr8jBoFbGKbnhO/lIft8pJt4DxBsknjphDfI8sSB4zogsc718wSsUVgyhkDQO
KSn/tchk0QO8HONXCYNLQAXAPR66VoZ3k01Q8RxI2wts9HvOEpsd+W//eDoKomf1
46z5w67PZlt4QDijCK5sqfuM048p1ff1WRMFQ/cjgY2hQ00/+aIpmLjRpnoQTZT3
1St7QWcoTueLDYbG9bS3aSALwYsNhgL9LNHI3pyWBu9I5JTpUCbSke7YUl1c5Tye
aElKS0KBmXp7Q0G1yRm4lmMAiKVEgsdcsvt7/z0zkfSNGNAeTtOFMEu1g4JZa9hm
u6jTGlwJs8GhoA8CtbT9kVMBy+YvPf1s7gEQo0TYDxlIVb8VyLbep3qcc96jHrSo
3QaqZ0N3RlRVl9P2jbMwuPwkOQc//HJYcE5B+kA0amQ/90HOF7vcl/2tiX+JcV3V
3tXlVw9DlwrdZE0zCij66VHXKLOFOGFo90zuhI9yrzkwSZRjtfXPhMvWmgR161ji
2VRR81ePSWPYZESXfH6Srroat3GrXC1FJX5RpH/OaGA9ijc2gjdFQ42G2KWlUBvt
VwlQLGpEBogWAwr/vwPT/3dm+Hw8J+XCvc9hEatMJrgCjzZ6Br3FDPUDay3ZyoUh
OXVtDyLs25XoaxEjlyqsq0lobIDcMYHiwHzHq4TY4xMiJ19dccVJMvTuj/0QCcGM
TjlqPW/MFFHW7qWDKRJX+M/S5ejVaEZ7CvqckuzWuxyZxLV0iQ7m7aTldSJulBFQ
DFp7eRsNxCKLgkyWyJdZAzGB3Ydkg/fRCcCVFEx7Ea2V7xhZ8oSWhHkqb/YD/aES
krF7OvsfZMOS3c6qSws3Ne9WmBapPsUnBzdMl89TXSxrdNZ1WiyNk/EiYwPWGf/H
sbt1hXt5EG2l4801NcYPuoHpOUYzL3IZp/nHD+SNZgbyIskS3Ukd9szsGYO2RYLL
fi9tzjhMdGZKglZk00Z/EGks0M0nmxn03JMYiCMcKru1jsHsQ9Yt4I4EQr5AMK1h
KyrKXqB5XUoW9EIw409OlTATdtyNWv6Uwn9uB5nzSWsV2TO4NfOx4YVw630DLQ3n
f3vQHAZVPi7DnI/RmqZMCpCUtIZ03X4SuyKRMwnvCt+IzZydSC/F1Lgzx4CWkYnu
UWLkEy31GSLqt4yzHm6xMUVe9+e6HOcEhUIH7mbRkId84yBjV2h3vIvoI0Wcj/PC
xuJ8J0bbSRo3lEV9S6Fsj0WWZodYzA2RfYlmS3psoW9ECiWn0krO/79CqJt15CJQ
zFVhav3QLGUwra/BiEzYd+la2DqnqZO9NBox/MN0ZnDTf/s+/YwbDRM1BhzAvGfU
0yQq9TISjDPZItmOhTkcnMTP0BIUggP8X+bEgBjF9vm/RmjUaEpHMw7wS/qG0Vnt
zV5v4m065uzQeurhqrbcQvsHvDc4Nz79JaLpERcF7Vc9P42zVcpHETZFRvQgg7BN
qEMloznWWaxNPPbKhuPKDvZc0Ezksn5CazwtLFvQAdhAcUXXWXKWSWSVFOziyPjG
5Fk6PnZ2qW+pWadHsbjjnlokab0DdWlUiKyZqU22qr3/VUGaU5zpqko45qIh/OJh
sgF9ke2hMsTtgx3Q8TFhi/1x/r7YiFlggi2imDNNFBg5/RcaQ2fThuA6kyRS3Zjx
PhzSXTPfGPhm8/ld0MRLuQbRtkqO8Vctzz/M4ZcVJEQGKXM22d7QuCWuPuI+uLEe
ugjMCAmh23+/eiTnlZg0o9UebVSeGEr+2tL7pgNzSyEOtyK4o7Z9MWxSfZLJG61P
QZBSrsCKMTcedmdym9tY6tWMC/KoLMxeZex9GNPN7XaIYMPf4KBawmvSJBf84Fly
4ysfvo0832BENTsRycFamLXHaAluRwU3CbozIDzASe+KNDNrb7kUWN0UWSWlbXr8
ZQ9VfDcrntWnZIotR2JgVQegJBEr58akneSKUoGcnQnJWucMhQdrZz9UTqVmor2l
01hK8rY2usbe1hW9PEgQTmN2hhE9Rl38vEFJHPHBa/OvOgvzpqWiSm8aQGhF6x70
9cr1h+hNgxYFNgyxUdgKaBuMWGALvXn9oBXWYpm10e84KC0TYh1Kgs1LdRhAINGb
RyQln39dzwJjtDuoiO9MPR5dN9E3bM+Lri+aGDfygY7/RMcwkHclSHoTFYAiv6SW
9LuSt1Ph+cA5rKMFWRqeW3amNY0Pmv52NWR9IWo/cs8DklubQfQjUcVlX3GEW7/l
2MQJpEXWLdgtcTHGuB79z3srXPLX1JfVqfYXJW40oAj/fX4zxf/tt+nSmggIlZsW
prtzYraCzM3JuhIgTqkzWXsgNzbtej+lrIhDvvSwoQxU7WSqBt9YrKimn0FoLrQO
Rl93+NDiXAGyFbl9cy2S5j75OT0kOfZn7B9a0S59dFpatYsHggjtlamUogiKtkMj
VMzsKzcF2/DaTi6z72ycLCRHgcroUCVtaQPH0T9V4PH0frdZIteAbz+2J/6XBs3k
voUDu7vC2HNsdLq06N46Yr3E6q9NGpe7Cs9XRv54SyCKo8xvvnFYh3FIZka5mIFb
QCGkmG1jws77SRc9tnprQsnhTqP8Ob4BP+Zddhzq/alhImprh5t/ktSVte6jHALn
KduwF1kDuDQBKj2mGUqjWVYP/ZA0CXXhcbmXT4oaoQmLsWWZaqetxo3ckhWD2CxE
QYWF6kCpAyqb8XSKLpwsUHX4uzPgoO0n8TBgz58jLXuzyZ/g6PxVJyfRlpbZa5AC
3e9i4H/J9yV+tEumcYEPKZdCFNZOlCCKfaw7ezevOZhjvlyN+wTqj8UmCGvOn++x
ucA2nhPoMcwZFyvvCtNVhlR/dWwmo94vZyzfWkM3QKxRn3mpvF1sRDMzkVc5VVzM
IWPMszztjDrIr7RRZHMoYi/l/RtF1dNgOVxJD+8lo3MBLOfZ8uWoxarAhxB1cK58
Ew6yoYdtdIh/WMZvW8bV5EOVdV1i2IjoewgJo/ijNPlN9PMm9s1+W6v4d1OdXS3r
JtV7QlnrlUq7oe8/6CsF2lrx6zeruN+VOzuAXV9deGG8T4XmVbQW8KY6uYSNzv+6
KabPi4d7gbuH9QReVBi979N1v2X4FSe//Rab2ba+M1N/hyyIMd6KeF+9roZEh8VA
7AavQMw5HwxxfDnubtDBTERHb3vjl81wYIf07D3s8xabhFmBir2AICwbec+aoTip
vnIdRJ8DZvHQ9rjW7ZjgiulUe68dbeqKVBiOrwpfyyAaz8Ud8WwOLdr0EhedJmKb
OzysP+9jehvg3oudzSWTtBDs2CHJB5/aEJB2i2jw/7EB3Eu7t+CuelgEMOnxXN2T
7YGAfPethYI2+G8sjh8Z2VIq7zQPq4od9kgaXfHh/1GJlSgs3AtijuHDKQN0XiDw
tRhCO8W4jZ4GTS6UJLfAHNvwMTpFA2FpvA8O4HcpLZqVjIoQivDvuZEBN4bsKLC9
7kPbofw0hv+rCi9ZSDroIrwlNhCwEnt9G9s0iUFM/VjF6TzavGhAq3QZZDqNj/FK
zYfHNkXcDzVy+MWKg1HvKFPuKlHJ+PYYOQbOiXYLNUpTIhop/lZ9O85Y5S18YCTD
/kWjWbwl2dIg9XDrUL7YL0zQc47k8Qqk08zVlyqEL16TbRKQfwM8VMFMEtyD+Gx1
OqpQQ+S37buq90y9PQjBrJHhOROYqVqnR6IXWkZGamq4COJwjHIG3dRNhnrx0LkB
L3F+JHfZ9RnqIpx+aZw9pVDMCYCAUB9cSfLdk/bd4nR/5SbeuafINCW3OzJWhUSo
26OFCgddA2L01ibaLtl1FYGpasqS40S8B+85bwqaiQIcTjBfJhpuHCrAwOlUwMRe
gj7uFzdCBJxwxZ0ZyjQEDUY2hNPm41DIwvKPVDMy2ABdfjiw4NT4g+7w0E5oaLZE
U1TaJbLAtWV9rgs75qBs8qpaQ02yXcuMEqUEVmRHSmaOagCbxuVOvX8aKnFjfEcn
g4PX6EYntiEGSZ7UwBJT4vVOFCrjMATW8F2qr4Q2fRMI3Pe+lx1W2PHOpgqYiNP6
7I18wZfJEUs6WXpLxMUZdEo6nBY/9dBcGql8S5g0NBcQ7EszeZ4zDUlndLF/6kFn
3X/Jy7fOM97jkqBy6DHvpGwUKIO9KnRohr0zrSPNU2cUv7lfDGotD4uBZcGq4Iqn
ouSWZdIqiseP7F7iqYvEZ0e6on3Ud9Hbs4TMX5utCj8v5R7V6iJDoF0kgpq/mGBo
ktYOqW8Vcw2/u2oI509kEginFBRm3HHaJP5bUvh9JDrwWfQPjlGv9M9TPPtjUrhR
d93/hkdL1iAaOnIMVUIDdRtdDMr+EG+29mEYDNAsL6d9H92gfHemdZ+dpaQkxP8F
YJgEXYPhuNZQRbkYOHfBGYMLDTlQNE6g/N25HnxrpN2ip0vjTI/TiGiyXUCFHnAr
4W/znzPeYQgXtUpKiSIGiwxUuIq3JINPq/RpC72QI+kZ4rHxZF1okKP37u5Yyeg5
ZkoHlZAHpAuI432Zy/i63OwYbrGb3q4xJKJ5C1T/ts8uLvysgRn3dtAgAJu3VA0c
LGF0h6hIOP5NnM6GNYb+wu6oddM2RszByLcdfLtXvgMph5q2kDTpnt7cgoks16py
2ZqOipJehbxFPItIwY2Jx59LLaIfeBFFO2CFW4NzJxqEftYJSKiEAmqGez4+a/Bq
dQafqJt5mD5ZjShQ0ZbBDdOtqZPeGcC4ucqS8YBxoev1dfCfNmmJ2z3/vDltlXo3
/wU2GvXHWejiDwYrkKHOpIiURV3N8lfscLnfAAh7nhmrLdyUBYEJ/vAv1CsVVVEK
taCBwz6+kR7c/G3GROxSsDP/ootXkBTIQncjEB0vwKyxLlpCCby1secIGCgJvufE
c2W2IOy4gc8IRIVHZJ2OqdDLMqr5bt4dzyqoB2BoYMNKejhT5+klHXjfuVrM+A/e
Rd25EIhqJ9C/I5+yJb8/SgGyeCHt6Rj2iqK/Z/QudyqfQFTeD5TaKx92ndC4xj+U
dPT0/SaZh3/gjetN1KfooI4r7UpPTZIEUDaQSaT6bMys2ccEPpxK/S77d7weHwBc
MItVkAL9bSgVBv2uCv2qW/tOPvXcQUstTWJEOTKDiyEkL6u1EZEp5fIO6Yx0ua5S
zHdT08e1gwtf3Cax13yni+M5E3PdoxHSV7crno5oPzqd62mrtCi8yPxOBzzokItM
aLg7f23Wz5L2OvF/exos+o55dqAb7hQ9La6xocpoeOkVMK1QlMkEM8Epa5Q1E2Sd
LI3IX/1n9VGiGLPvCCSHZxj53SE17woGO8J+QDuNcTXlxtT7XieIzl5H53iS3X9L
lTTCRQZmphAPKM+ZX7v6LXDSldhO83IC8mqGvLEqMw/QT5w/N5BicNxnVae0fKm2
5t6U4/RT/yfFj37MndMEfie+Q0OjvolTjc8C515SRsXzUY8N8xPNBD5lQej6INu3
B9KQgaFWTDRtwxssrmlB3KJ4jGSdOSJvG+vE4hh9YXtadxbsiYQ3J4deNW42mZ6u
rkgvJ6rtnzZNX2PDLR8/ZB725oEBG8E/CUQ6egMGgfbPLrrH1aTUdCy9SqAO9IFr
EcBgNaLrEPuz43xaaTnMMmSqMs4Cx29qIKbIFPgKqsd5cyy7JdPIr2nzFDtK+fkj
iuypCdMnRa/XidLY9MVPwARRet6sLOL7zlYVFmKiZ1o8fgI/VVElT5hfx3AyO2Er
mzovQCxGJnhxu8dx9Fsg6/ovw7qnoGXXGaJVFHpz/yQGzZSczlQlnq1i5QhjzDjl
4GoIioEnvM8lUViNIz8i64casfvbtlf6WqnuMWx0dU61Txwl0EOeE/ooxT6SOVQx
tkqqNSsXvlv3Ow86dab1hm98IbSBxZ5Mm4UnXWILjaQXhm3rfgHvaXXSc3qLuh27
iKyllg/ZGgPsLURVwo5HVlBebdRiMuUDS0aDXZEcBuQ9n0YOY8siqKX+ieOwGfqM
l82obIgqAA+0fK1r77tS/wfTV56+s172J5/D1taPwvNppZ7vEtKdyS4L1cN8I5jg
rkPgrlEmUe3KqH1UvnIO+XV/sjTSczQOgYBPjGm2HzUBwMpVOGSfv/yjQpLrH/7u
tTVG/w2P/TmKr6z54OrrtY9uciaZMF8cjrLDVvM/VoooyC9n1zQVMwtkVRe1/gRo
tsQJY8cFnVMsgm/4TJ2OnUr5qNM0mzqdUwFUVFBRSRTOfqL8YJj2tjgvyz14RNna
wp6reQ5Zhs+3ijIybULGghzGJanhAWAQqOcAnI6jjDJXyAPmNuWmGY8iQrKxySat
SLkoZPZmxbgIOsRfVPhGDIHOoomhTsLgQDlnQLLzGdMzi7pAJ+s5rRsdP5pzyE7N
bWcJvOhdgUGHfb0vkh1zRQQ6IMWGzUEWs4wFZr7GKidiPE+IDgf+r7ouybV40o4k
EgbMwpCRoujzAk63PoIVbOBzs5xNb7xm72A+XktxMT1DLMZ4bRI4HmMXz9KKWhu7
oqP85Ax+iBkrw684XxxcD43D64Q6eQmncuenldGLh010GPB5YzIhmUQU5+8Ixn02
xqmJYUDEVkiK+AnnvzE6zrXu/gKGDjwFZZFM/rTIPv/CwME7oflAnVGffZAxbIDB
yUOAly/7AfoB7zGujPUKHXw5Yhd6RYrqgVUaC1vQ64uzC90aCO2o62PaPIS3P8i5
L6ryipB9Wz81VUwYg7Sg9jeLJ7dPJuqK278Z70cnhsOpVcFjydi57lR/hgXGFEGs
ipegK7zNwd/B71afnR9qgiSfI1TUGsomIn4PXIxe08ZRL1m76jQwdGzo/6jRX8ei
PUKAKm1s2aCxF1AFk+oEWwv4SvXl1U60mfmd0Naq5UNNkdNrysRWIwQ5KJE2qBq3
RwYNoha2gcILf2iCT6PL+Ujc6iJajUReo1xqHeq0zQo+2gIShCs4rtjq/gsbmIkU
3+tOXmjBJXU3PMTqc0bg/KA1t0Na0ckBjFyQrlJ9Ia6roK+qIPVcSQ8LY/vL7NSl
Fm6DUql2q79ZP3K5rUTJ2XBu+BkBC3vFr0Bz0jTLCGjK9XRR2NPcQurf9ItyRiWu
zuyLXHrrymTCxqLCVrfTgSjjmNKmy0IbMVQenhDMrqRPwrKvdl0WbUXmrGNbQ4F6
S2DssA6WZ2y31T7+X6LLHyISuihtBxI+wrjBy92mRBfgkc9Omvpj9oNLp0F1ghTv
jpTUJdu3a82E1Abvr8BSZi73Jb2XMpGQX5yoKvmXKl6LQDgLp1M55rkA/qxqAH4J
nlYqXotP70TtFM6MXqx0riDbrUwRc3R6wFHcVhK3/Km42qYjC+aW6DN+GjKIjOs8
VXrQd1TMVlYflZ8TeX1nZiYesea3jXJEEq965U4JvSAXpwqhp2DOYTuoJHJ0Euh+
xPjiddicTibo5Ewa7p5CgvSjXpw+02up0bgH/FZVIipwQiiHwnrGE5ltf7mPX6Wd
qSiSDiGpXKvO7LZTIuDv5J2TiKI5kzI90sEiOkPOoqc78l6xI7PGIcWrzj9fX2n9
Vrbit2JJi/vIid7ABAILdyu/++/mrHAPU4s5H/QTBpTo4VF312V/cjDbvt+E7yyw
HLKq25WkeZ9WAJ4+YKFNAVEmqlT2R4YooNJKsQ7CorU9pKk+Huo8LRWWbpEWJ/Op
rB1Y93i2r4l7SzcT8tV7l9wJKtrnqfdcG3ojWA4DARMrAN2V7ZpJ7JuktXPdgI3H
PeK2885zz3dlQl8yEEYqnwqD8/jh4OuOlnwlF3DGoLOAALcU41k38xIpVkdFrQCr
cnv7GEw6DlQKOV8RBhAas1b+FBd0A9vOSM8uwNZWm6HCebWtrinku65b28SZ5+LY
CkbRih/ThmpJTeuVz3XBngkezjTQfk/E/E1tg/og0Psk5kRCZviIA2XYB1pjDubs
l6H1T48Y0cYtjeqjHstLmEkIYrRAncaAsORQ/8bFnDsM8uFkeMNZ5yOP1ewposq4
I605WqFOeoTYnzL8qMxeeTpUfwa/3cCgPpatLlDU3A0XGhumLzLwNPbrIMinx2s7
thqxdNOszrLDKcBsUc3cWeyqRrCFSBkCmGW/NH+3k6znoeFxIkU80s5bzG8DJz+z
Ki2fPjboKVGG/LkYxOnYODjtWppuzSE3VWqgiwhpNoWwmpBYHosCPNpY/fguC781
32CxDymM6UCLUemqiAi0xT0V7Gt/f01iI6gDNtIFgx4c581pOkwAybRjgB47dFmQ
jR3rs3LWK/N/UyaFsJt7ev32i9PhQ7h8r4qcMUiSJzrI45TXgOkqzMSNVBwy97z6
klk2TQjxJWMiad9ObT/fZpN9IUvXnzPPPToWIfa64Cg8fzLib4Pq+WJDHWOKtDmm
n0UuSs/X16gP2As6cRU4QVbIKGZ0egggIihBWvmnH1HrC8JYMCLMHg5ptKShYW+u
Hzy/L7Zin/9nED6hgbALv0OTEJiIv7t9DTmvDIoJ/tyfQv60GkG/iKAg6p2VEYXh
mD/wfoJ7n0N0JVSnbQpUssDF8QpByF+mB9Nz8FSsOi+xxDi590dMTNseMXvmGQMJ
f+HA9RxXjbimTyosSTY7wZ54pHGigOrfwMKwDusCZp6xUbZ6rcGOVneQ3OksVp7x
7b1A5llAFoGSuoPJfZ/fv+qBK5HizmMjwmwtQXqbEMSKcW0trZCDjihR5EYCYg3+
Wd1hfayrMi0miz1bYc7Nn2oxO/2vphGx9yrHCJVdtJv3BRhkr7Wj115Rofx0Jp2T
aBz22V1Qe/rwyKQnrNLA/Exne69To4DnGPMYDz8oMF67kTVT2hgPGGKdYa5XACGj
Sr2Wwsp5Wi84SRvlNXWUWNwDxDiHB2qHNGDGozkw0Uip7faw3rj2TaSxrhqKpEc5
ET1eLdaxX1h7sNyDO3JxEU5HpbEzThej7LOKf53tppqflZSu/A1XY5pRDU8a12Kx
UP+qGwgaX9/+E1wX0utOl0PAcCpPGOvo02Ey5HfVJqZdgi8TBG5jhYxIs+2mS2aS
tBnRnxYWSwRyYyiCHz2lJS1+URQ/lmN5C4X6RA37eN3p4Ha+tEf6vQkRe0lJRAMo
Zstas23f2B3jN0IN0jIfof6mQOuxgBBPKqnX8HfdsYDYBLUYcX5Q9LLOJhwNJJKH
qMXkNNISPdyvSvdZDs4CSA1AGxGpSxZ3EloZ/A2Y96lAAQTBuOIIs8qAJYHVkpLk
x86iBpZBU4198jxsrLfNZtlGCY2E19wMnr5FN5sxwuQabr9VPYr+m+TWkCcsfm+I
lKB6p5M5Jydlv8GRMa4w014uqVpJO1CBPGX8bfFe3XMKwjzSZeHaUUD/XMpEwAhu
VbxWe9oOxSrlq71/wHuDYbMkCGmOCeDL0rcdm6E5kJYUmxi4fpiVprxL/NCO1xDJ
moXlpRi9WNGitH6zJVls1qfNbFmDWecEggoMoJlrzRI9A+CU8DZTfbC26iv1z3MH
HTKYOlevH9CCeCJeC4gQY+h/wFmf6aglOLRft16PEr8o7A3P+KPqxf5NrrYW+9SK
ZeHzY2NZoOZKGf6BQqxUJCmWNZJpTvidulC8iDYo4Hrm+ez/PGYruPt9dsV0T2VF
qP4aUvQ7x7wLs+vMpD2xZ0nYphLr5ViKpouMhl9pV7A0MoMJXC+NRwtrs1uDovgE
Chu0gHzRDlRmEkNuRL/k3hXZYLfWgwqrg2NspvLJwbRKLrSGOADTSSYPG7cOQ9PO
x9KKJDCSstmExvaopXx7lbjOr+p719ecJpy8/IHMCv+5Wy4ntAVyYcZEv5oAvF/U
VopBGidwr11NUhumyoh5q/gJ2GY+cmxiv0VJUswezbeAevSwcmCgpZrJC3plyJhX
CK9BMoT2KPlf33d6sWqdaQBQQ6zXQWItD5xuY77DPJEKTOY2hZEvkXa17+WwKHje
xLpFsnUzcwEq3nVadYpook+9bs1aOATfPthE9chrRoi4IFyqk8b4ZCebMPDvRYz+
aKSe9t1Ddkz7s4sOrfbK6Isln60GwAmUCvYncoeAgFPxDHRmogfAXd8rmYs7x9+P
zqnhHlbf24AKq75FDEx+2GwfvCWNxD402jk1Sw7qbO0AkPMjS1qpybaqfnrJ9kyE
iqKKE8BeqE4ryV6YyoXsbTrEhTZGv32+xe/qxvvWrFcn3ViAYImFhunipE5sAvQ9
TwqDh350FsA/s3E8KQmFoYua7ATxIZc5Zxt2N2ydX2nSxdQM5CDUBI84LgUU5RnW
a0m7wM4MN0BM0nSX4TgIvbtDbCrqPxbOvTYzPI6py7P6UHPcGx25Bc+orhqzpZRJ
DRrdZbOsXWrZyCwDC6GVc9hYq59JEhO5ivQcAZ+A8FxB4fqsPnsrGRc/7jQakkal
+T2p5IiYaEONlaPH/6LHktPLXfEap8fdUvF0DnRINL2VmKIglkluUJDAKcto8+8C
SbhvGWHFjnUPucsqQ5FRc4TyV//hJYwo2QTqFMQot5Cl9RlQVArmsDwiuWyNDz6i
xwbuBodT2oy6nn7mAvbNx3T8uL4kaGW4kTGyLdOfVXkXz47tWwnTJycSc9/lX+QY
vMIKo6yZQcnQ39u8tU37xf4c/+Vj9XcCrUnW9mOxJN/Vu5MPbDnA/UBJxB6UhR8E
wMbl1UArRSCdNXIgZKZ0RvaKpsa17sDRIWd1igujAT9MF6VLM0aLeK19lbKvtb69
Gjbm8cUUiyF2LmtJzi7qspsBJK6F438X3xwKZveu285wMJmKCUp5wE94fZTa0Lpb
ciiXIen6GCAzJwUiSfUAHjyiUeLBrs4P5ZLWzAYWTC0bIGAG7Iisju3OpmIZoh2D
qn/1ZgtjSY4fH/LWAbopt3YAN1fimB4SP01yGV8cpWd10piVpQGC5tQnfOCxCnP0
eDzTWCX+F1luLg2WhO25HG9Squmgfu6HBp8i479foET1Mtiz4xrAAoKd/FQajy9t
88a8tUdSNCnmTyfC40trKs7+jstdppfw9oL2VBvc79lgDNzHi0XOFdu5moisNCnd
ZkufI1EVK1Br7PnJbHY6MDw8upJubEp1WMfP029/eEARzG1uVn3HpE2BmH3sHj5R
5Wt1o+obFTTpY0+vygKqBHPS5/NagC34bVCvVaiBwwiu++mmEoeMlXCmgHzf2Llb
VY2W7iq7qnhLQ55XmbrokskstfYXV0tH0xfW8OQpvTWdZrAthpv0JAeDpHwkRTqb
G4s38vxakDvguf7eDUUl8nAGmj63GE8m8dgYdKlE8/wuSA7mdGAGWEVx2gc3Z6wX
NvhPjkJ+FKSDum2H1/BbclYWsxWNyqaoAN9VjBFuzBInlk16+Q/xXfH9vvc8MWE2
bs5x0y7K5cvMKsbY+Lo70gXOqgAM2wr43zT3qiRq2GmDyxGSoSWQXA/Op5kOC1Se
D28Al+NDfA5Vp2MZhXputYIJy0B5kdU8zH4gmLoJr12Ubvq7nNPYqGucJPX52V+U
Aflz8UqdSuxxwM06hfSuYA0ERfwj/SNN91RJ19g4IZo93xgzEk6A1wQcHAsBRn7L
5o0evAfZiVtfHZL60J2DfjoAfPGo1z9dlaHvTEkfJIqK+V7ad05D5lCmhF5aAFLq
2CGLOvtYi4WU0nt68dLnTU8IB7bk+ishyzHfEAeKbu9XNmmAemHPF0sPcRZ5NStq
H/T5dLKkenTYQd7YTQ3sDIai3eQ8CgdDkzAQ3Wyj4gs1T0WZASnqF8JGBlhBCX8V
UwjGo1LVVWbG4HEQTFbIb3vK0E3aZZmiA6JQecBbyuQsH1PhY1r+rHliD5lKqnru
YbhOxpTsiGgpQ9gjLzKfPCl8qNc/fs/AQa+p5xwSkVcGV1gi8fPGUxxyKz6o5DhH
bFM5p0S7eVV9RBwmuXnbY+I38RY5gj39dNQQ3LylybXVI+LhoBwSqIuFK90H1Z7h
UUAarFBA+kG6k7kmQLC3RUeDRiPwPNY9w6nz6lnrHOoALHRlOs3TXVVh2UOcmKmT
2VLGr+1Fx2+NnWulWndJ3NuHMKtEfMYYnKxusq5H7FlPXeDx4p+1xxykQhXV6YED
7Pu4Fm+WzPcGJ56tKg+mQVUaWlqYroQj/3bJTZ39LNAoRFrJCAnZQbpNRSVLUv95
PXVBz/6AivJi0gueN/VW5MFKL/MX/Q/4c4/NVk7irdipq1gqPHom5L/iolgQnsBM
BCEUyOdZRqyQtD+npVgXympZjPIzzFw+oaeZTcbr25kWxkVTHUEJwTjbgqKbXC7s
WFFqLEDP7Ul9llRGD5uQGgMc+wyDwM0xmFDcpHVsncptuEMnoIokJKfPNgHFkRHF
zA+CDQKGrttj9CKBHnCZX018N6xByIWGmc7naKx0L/PPo/7UFRGmmCkKp0VX/eOu
TnSDJ8JqluzIEissOfOGk+2lxA21q5WviZnUFxWqYnrOeaIwVlpFZccFIJpW6263
79a583QpWWgcDGQL0PsfgG9YLrF5l0eKpUeIJ8XT7LnInf6CvSy8pekT8dUfRpq4
Y8wFyh3InDdBL2jaBBMTtsCNMGIVOaoMLMzObD+MEjSbasJ2cnP6eASlE8i1T7G3
/y3cCX+dxGTvy7IsKQCyaXSZVHhKNrIDvoQNM+h4Cu8AGuE3VcCcNVwR72E6lCHC
TVBYoHNzVYKhu8vy+M7iuhFIIHteB7yr8aVFFptkgXVZpJPDQIn7r3nr1r21H/OW
XvkHwmQW2erZZvUFO0Pyis4WHpDcvqO8WFgDFVv5/G/LGRxlFeUxmC1rQseJFDZ3
GAfL5aUFAOSVTTdRcM8aC9HHA8dDEXOXubHWKEQrxr7Yx/Tg7/MHebkmzX+HQY7+
IzJsxrNbTpTJazoYBP5xoJX1zHbByPksGi9STXRHntQaiYjp/b5HRQhMrYcSPahG
z1PmPuBdP7utcQWjjfW28iw6fL8JllCFWzEKQGJefnMvNKVG5HLR/I/O0iRc6OwV
PpIrbIxEJhlQ36myHikELvwRQANqPAc6jZGTuqT35NYwydIegJlROp4Rhzbd7mvx
5/PTL6zu9xYL3xhQqG1wGnLnruQkecIDz791eVqMWXKNxxznbi1oNRzFYkGwawHW
dabeRVpMXeB7JgcCxjVsEbRfhwN/eobcXlSLa+weLq3qM6Ne6HT7d0dhfODDZzTS
dpchip2l6jSjabGMOjCLUlW1SbY6ppnLmp86djXgPsl2FyuEjlOCpotHzTcfxO5b
eq7prH9HWurNRj8aRzgNdgus/w4ETSTaZdfWrCV94d/Y19wxu3nsiIKE3X5ikd5T
PMaygD7urt9U7HkY8lj3mgVHnyI8xauEFh3qVV1eYCW2OEWbZosDwNCCk+mu3eDE
eJFwBCz3mT7jYZjHQwJ2Hn7K14eisQRiJgd2AF2rZKSIaQmsEfc18uJifA9d4R54
PcLm0SYLLIGXofPb1MtuSZpq4oYJD0lBzq3l6et1DZhfhGDkn7DArB7TEN6E3wUU
GdIdbDLkGNh+qHq64JiVWHmsQbA8NSLEDL9tqGuuJCSTaX+kqmpYKnIwPfJ3JiDy
L5S0v5Wl/kL6kjCf8Bx9+zK78ElLuBv1zFIVGADNUtcSBeDH0FEL7nh077YvWn3s
gB0rqVix55F6rBjsXY7FzsMIshOXXK/r2FopdFQlOtFrglwYo0eF9V80apVA6n6i
01LdSqLohq8mNln0AUfzRbKuHcoPxSeYD3OkEF8errCD1q0JzoLjDGEQ7k4R2zjJ
5BDtsuNLQMB/81Frl5d4xph5rfnqoFvP3l5j294UNf1b2ESwiutU0CPJsR/8tfIh
5yPxgFStmuX9umU96bZkU3Lj0leW61cQrr/fxpje9fIsKkA3zcSlCbPQKWfeh7Pb
FrJ85Ueaf74/sr+6qN2Raq5KOtaxnoDL0CC64/pAUyTOyHdwbCNzfnHsy+6Xojp5
DjMnGlf0s6236DdXoMcdD/vesozhDW5MnhiBpsWrvod1xcmR5JfETW3RrIscdbnw
XDpVuG2PEKcBCqFzIWpsDNrBTrWzVvBhVaKNRvYw4kSYgFF4NUT45CcvkJOclBc7
ZxdWpa6bnefki5FZA+Ng9Oh+UYI8EHC16g4xk4lklXgyK9oT0B6vhztjzFp+VTaV
JOv1+S+ThFzBsMo2t0ZqxiAogWl8itPkneCavJa8vl9mZWDL/YVWP6rh5kSglVKs
pxAtIWsumFgiIZtg5GULxgnbUmWBSpAs7ZMBYxd/UkSOykbcVO3lOA0QUQDt5K6P
OwDK+re/hOVIwQzHJLGopD7tCpn3VTjvvsgoVzk4uF7HIgjOibj1VDL3YjAIpf99
mojb3AfZkOr1c0rkgZX+DrQspTLCd53QrNcE6fGGdP07XXLCnf2xNlqC5A2FEqbi
B164IpdIC6MvXxfjgZ9G1L3l0YSR+8frZis9M6hNxcrPx2hrU9uG+vmVupiRDkvp
oepKs5Vddsf8lSzmNIYbQ1NoYavit2FzWzNqGpao/tynoSDoytUr887yI3MwR6oX
VkWw10Gf56EhiYfz1soocTHnVbpbBzLU3zeHqPeDFlOgu6ahAX3wFXDR1DYdCsMS
+zV8DC2hIu8JITL59G75LrGlra33T2mhgR6sOttzIHP14ae5TTTN1HF8k9LBDEQ/
S8/5V/kiAeZ+lFdHl6SwkwuNAf6NicwEbPAD5CnSuyx2oPZnBKWc89EbxPMa9bBM
22JeiGTfM0o1AXnlwTolSs7eHCXxd3EK3PFV5p3WRG05spqV6hTdxu2y/XlUKYCn
GpIO9Ew+gUQ6S3uTqSWnuTPBWQvcqJV183mZDrKOHr1ls3ISwBoeXOgP/nH3JzUz
fZUb34R6ebj8XDTJZINBvD1UFBs1E94AU9y5+zVyQAMf+pP8wfUm9hL4eHcy9h89
GwbfnbxlCGGlu8lBU7AFhqOYBfwT5C3Pv4ruImU8payKGrgn6OGMtk6NyIlNySbd
fwK4qEO63PST1XUFbIyp41ulOf+QH242EqHvm3QKXfIgdfyktIRFCRZ+2RcYku54
Wf23L+0AoJ4Il2sS3dfoUdJm8pI5EpWLcTwc0iw7q3NtOKosQuwXrKZHZlOkrbuC
vKBc1OW50ims2JiTRq7LmIwO94GhdJLWUM/cLhMANW6dIQcoaPsLhklVKrJHls/3
zlxGBGg7jEdcAlAxv67myj9KliIZrHdWrL1CaCeqdZNdL14LgcYp8jQu6T8YiMNg
yXo8rX1Dz7/o9/GzCO+A1LiKhAjJ1g8tYSQzkcQ2xQLWQfthyclehJy2B+DHysPp
PwSYVX1EVvXBdRI3Xsvv2qpC2dlMpstIWvJwtAUrxR0XnUgyiRh+Qduti5ctRiVR
byr+x0D+OeK1netkG46x8Jok9sPNGlr9oLaoHK0uRk0CSUznhyyUlAbwrGW9hrhh
O63MoU0xg7GFdhntMwmzGJ9QFj8es42ttPUSjudoBEP7DQink28uD1IFAyZpRTTP
miABEwOChQFQh+74D13eisszP8YM6SG12KR5oj8iWal5A+zM/kUR6Ca3ZE3zngTc
BllRc868uZhl2nqZlCrXPDTpwTfVdCa7xbrMZWsHvw2OvA21cCvc/qNsuewVtWE5
AB21T/nsJHXnxo1L/93Y4bwPfA2NKst0JpJm7jqxk5tnUeQ2ybv9SxZx+JClEzFi
ZFZdADjqUPzcT4iGrCpRDWFv1m7NJdkuqSJlM+BMp7d0X98sZPouGcXqWqcE6vQM
CIK8qiYkc+ZuD6tKvReDUpv/A/lbW+rF+uGbQeJPC5K2pPMPQzwj6jf4JmJkjP7l
3pYNFx/M8bYOW5auUF+bApqwhKixBibQQiMxm4u5oYJo2of3uCvvlgC+/9na8d5D
bd5CnjZicPHzNNEh9Z6qhzurlkVlxd2xjMllX2Z6vc8K+b7DDcUYlqexP3lPIUsw
7B7OMzSsecxY5Joi//I7llBoPjQEe5+dNUjR0iKatQqkauW4v2/BALOpa79pYs1S
E3A5ISf96BnVPdFLYiPjO9944ghyKujKzk/LArA8tHe9PvBTNn74qFcgwHcJSYXP
vpT2N0C4aDSxGqkIC4Z9ep8e6KeNYx8huBobTEddsVyNgOLPEChE1MlxpTau8hlG
LB2urHgrgWXjM7sTfHi42exvZ+vMJQX5uFmAuXBSOFIBYh5dXok48fjDt8G4SyUI
z57WmF7a058O5RWt7+3ux3NLLEGLvZpjVVpl1TFhQU2lX+4++IMGtdYjeOUHBXCi
G8qN4sAE7r1UG1oV6JOtPi3HJHeWAGuPZR09vdiWKXIe7z2IKwDj0eHtaYsQnGkw
TQNBkZQvmp4rdtF5gOJr71T8leZTDNltxvehDSM/t+N/XtdPoI1c55a/Llou90Jy
xev1NzDJVdttZ101NigMQpoAJXKRqN094r8jP1U0ig58l7FzCrH3ovxis0/Ct1xY
9n4FyvppypGsCArisSWjdsvcqD04wKkocYAMhcENtDO4MFHuzJjGOCaHIP+snNZY
KpVHjXi58FKIyT4cz/Cph2PNX2sEnFPf71js38k1Nb74d2Sm4benXRWs4Xo8+Hvr
W9hbIQLVl08Ci7Wrc24ufeK/KLe0KS1CIr3C+ZKp0GuEFu1auqLG8lUroyyBIWiN
V3eBv7axtVb/jLYDYr8Kmf5YYlaQY8rXZirA0ANZch+el/6hFrKaEixEkwCcI0wl
cntqpg3mRaEz7UQShhtv8vM07XcBXYcr3TYU9ihcKj/GWk0oZi3eeq6cfKEMXTr7
19AlnrjkTFZFdBUA2JdacjBNLz1YYA5zBBAEtc/6UEEGdJvfmGkHUxaJTgljFQAh
hMq8o9DD7JckebQR4XmzOfc4F0IkzB0j1Bkp29hspTMpYeFhw3HbItC5FCwHU2Zn
3TMufQDfHkD3MATqaLD0lh7cKdEG3iEDbgjFFsrbPbBpnaN4DTVZm0f/WSYJLDtL
s3ASX4YjI5D5/VskBXTePBX45H/nPN7EzSQGMtDOBpzVBAuhLyPaol0o5EHwSzjI
uxnySQDMsTzZbOCgVHeMSVUsRw5EP3cYXOCripwqiqKVZZ85n0Jcsk/RFgVRu8JI
GDPvTohgZ5XCxDmnOPy8iZnNq9gZMBXRe95x+EBBiJ0yXnbNMfr6NfBfC+OqBPiE
PAS+wFuPnye1h3wW2ppVGq0NzU/qNKe1857T/1MqiI5FoWlOnz85zAoI6O/kBjOh
sMtspSb+mNBAsBfSUHoV2EArKJpSHLcd/QzZ1/Sj0iOotz4xl2aPRrOgGWc23se4
PTevccwmGSIYk/BkZXWvmLHsYcFCF4ff2mhQ3EVeRjS8LWgXjL008lp/RE+Ajzu/
23bF1S9K377G7ARBD0XJOqD+38rQjtJU4wuSWl1Efjb9VlQgPGchwtmkmniiP4ws
3JrikTTyWQaWSmWayc6yqLBAyLQWgmhmIAQKLj6Zvw1Bl2WlLaLL5gTcZjm01XAI
/K5eVGuJNZ00ixKkjjWG+6KUvxTJe4aEtR9pAdGsD8xDCEgUn+q7Ugo/SWQl03ng
Q4QMTlYZK8cQ3a6DXlM9sfKqUpCMIUxwOPNCylHB6sozSDfAo1urJGzqjYxoqGi9
vO2b7jTctAxKp5YkDK+NwatWKgQZ23c7VutpuYYmNu97XrgMB66Vuibd7YTNqeBR
lVvzQBon4e5irltLobZEVVv95QPDpdTuj1UorgP7V7G+TJsMmMIUmZUWS4Cec10C
lxHVHm3cAmhIKUxm7jM3uKGOgFGZ7bB/d2ysJWWhHe4i5FclsCxpHdr6OTcxHoZf
bC+C/zanLMlEYIC1UmMFQSv9vELwcjV1e4KlWhULFvJcRqVhBzpzHFBqOqCQ/8SK
1FR3e5OePC2sP8pfAmczCjhz4MABmpFZ00QjD+GUHa1OcHZ1x7pIN7WuV/4RYBH5
B87nZ2OGJjj8nVDX4nmqBAK0e9ANCl8vGPt6wn4gVlNAgKK4FwrozjCuVyfMryCM
IzEgbvODKJM44BVkED0ua+AuqEsaMBNrbWnzqXX94OQu4411yZMErqmz6rLQe/84
Zjw/R6wLfgBZdM/4NsjZ8/YUS6YiUabGHYUdlqzApwUh3aZuN/hcCYPF+clS5V8R
CZf5K6AJfms4hJuCLF5GvGLDNkB8IyFm+oXyNhxZU3Cw91FfbXNO/pzv9+z8io6n
jUHvXEzrUzbM9HodvwgkD0BY2UD4pIBZ+yrkW7cT3SUf/2nj0f13jc12+ykStjua
eMoAJtz2JPc93Pl7EChLYzYIfQE8GPDRSVKNemUWhtaaGrQxOm9CRgkwclMPuAiY
AZ0enwfv1nCN2LvvNUakMHMWapkqE4A4yOzJKZlHoIvMujCAExmkixXKqJpNEHyw
pGvyoOZ2e5BG0oYq6GbO13R5YWD0PFxoHLs7geaVwPYZzThUiOn5E10gjfILalBu
UFvTumlj3ld4fEjGuNbgbY+hYdA3w90HoZzJg8PNlwYEsvIbvbqbF/XPkD9uVj6+
qk+iuc21uTVJgO3Kcq8yYtJt2S+JFNxyoLUvukdZfh19d/ky09bhzD6b3KE4Tm43
xKrIAj87BZkHI24fmRxxBr2/Uw0W3EnNkAAJEyPhIhZCaiFx4laW1zq0Z/61C+MB
+urM08v7LedbETB3TXJsjFnqYRtdUis2JMWN+BzluctkvNJn99ffon6rYZm3eU82
3h9VWCkEJM8CMd4E1LjylF+56W8Nqx4uW8hQwnF09f85NQvTwqWaC/T8mQT5Z99b
3Iti9jUo0Tvzv0go1YaQ4BDdWawrgZ06jQYjkvdSOP/9gZ86I0fY6snaEOPeTzyG
Ix7oXxX2ZZdZKRlQJV+XEsFjJum/MjvqHRxbpWShTjxDOMSgxLTosIifHKAz6swA
TmETtCP+0hGJQkDqroTr7Xt7kcYAykNz2yu8hR7mMtfXBP5zajh3qfPqWnRGbOrS
eYrZ15QiujJ7mwPXzS+TB6mkvNY0DogJYR5ranQYxzGVmOTLxWz3iZonBoHVXt8w
j80Q5tt3HT8v3qIpzrnR+JQOP72XaFjiumABRxicQJEVlQJzcTmb7W3O1WmXiWL2
8fGTcqzoiI3ZXpVD3OZqvnCetfPk8kOUshWqoOtlew7WyAUYOYocuwSUCLajE2TQ
AklEAVOQIw4FAsjHFoNxNZihfiCH1R0XfgKNGtLBK1tnvk+otujNvYrzSPDIAbLN
PIbUDd5YggqHXX7yANLIEPfYqGnffbqf3GktS9roWQ2iskPYQD/LstyCA4C56e0c
5ouDvlIauinhN1nNtNz7NXQAs3YSbZ5Pc3qFEetBbwBQ7+Xnt+gU5M3JIUsdaPOG
3+eMauJjjY20k7O0aJts8JheTvr2xQP41w4hGOtUzHfj36MpeKzgG6JK6aThfg1o
DvRQwQS0WKKBr8UXzNBwfApQO/UaomkKfRxK50XtWWyoxvZoFc8n99YYoW/+Qm86
+V425qiRuvzF4gC9G34DHmb661E1K9UQrcV2G3OMvhbLOP5H+Z2j05tYtGJTkpRQ
CCyeiik7pvgY/mrxXwOaV3z24Qhb3AtecfvL5bkn+AF99ERSldhd+2bMxsdTcht/
7oeS2KIp1Mt0WjW7ssh7xxpoBmL7KtvEwVymGU6BpEas1/dCo1dYFqYuQxjIxrgJ
M/pU99tP8tDYxn4/YJsuA8apiVq0wO5Yv+o3IYXfNaAGq+jRB1K9cyDyd7CmIBig
YwRlhcyAxF21aOJjhrdQPBRIlyYCtuhWYwa/QkNKF8Vhqxa79gRqs8kQCPnGtMsY
E4QcOWdt0DZ9N+PIb2+SMnfgt3jUZiAXVVGP9OtjFw3TuFatCBFzkNIzG0Y10sDy
ej7l7TKQyjIsEtJFKShml77j9iBvapGYAyYvGVwyEfhzjZ9vblw0pLATEvulk4Nc
XzO8zZbIy5SE842lZo8Ar+B52hYVfIo5gypRp0Te4EJmBTM2dheAfdUrnn6ElU6E
eroZp6waZJwtGtAKAim70VtHfYGpnB5DTWkTzG7300/2b1UqKj6Wx4gapS8dAqnc
gG1ALY9DQnvrtfvW6elNP7lWnErilPRoR9/+NGgl4goFpp34NuD20U01X8GxlEuZ
9pYkVM/GoKsJfHoocZZs4I+VKXQUb4h5slWAL/2dilUriVLJY7idhcWQThlyVB39
bisVYUAdwXRtC5CcpKMCDIFNHoyOxIzoj5Oo6d/7zK/Cgvsd7Kwgt0M26jOe13U4
B2/JJ7RDZENoFx39Y44Ab93D0StZYR7YcI+0WTYfuubdIXggeh4du706ExL1A+Fs
aCDxIBgkt4OoYPxE1kIro7NJ0WFF3aS963/0RrUGgmoekxtdpICmR801sodaiH7g
mR6q2jbfDX0Z+0UMHNrGuSWfOY/qy1LqkCYwKAJez9AorLGluEkaCTdAPhL3zUjH
NnjOlfRr2/sh8Bl74nGqE3gRNo9xmyM3IK4XuipF3gEmphRrzSqizLEHtLw9ywmQ
9gCmz6CvcgmbwWbgLKxqZdwFBMpztQBFkoNwn0so07hoNJIRFAv5QPgkMn/4ssbB
r4PKgRVURWLRUR8bRv4vR+YAlsyt4Lmn5ZiZGENPcjO/Wj/VyZLJOE//gT8PzzL0
LVNrMde+MXzuZkw0l+n/CV50smri55oH7aP6gFsqGVKP2gEAvBLV5E8+Tj3DYmav
8Od2B00LDS/JL/vu+CrdaoBKsG6Zlw18OGANDacyyp926/feQSTL+Gkw9ELqH7QZ
PsxGR7PAqVbO0033LPH/CUCCeKI5FwyQX2HsruvzMTdalYv+i/vjiYjPPXyFox7j
AbR1cUlLodFQnZKvIOriFmPrwNb5VblbPAhW7jFuB5FKg4Krm7DoMBiWm4/I4YpA
fDXaAxaZ3jyE7lerIothtbqN36QJ4GNU+3Y2r1IPs4dCEf9E1TmHMF1yLQSZRB7Y
wDoscg+AN41QeWa0GbtE0EXOZDKqD0E8BlxWqiYJB/9zqjgqE2P2Z45pTQzl6TMj
H7NSYzAY1pbDCnBD5gFhxLZDcN4YJSlwmuH6eJ3ZMlYWWxdw9fBluvp3ePu/KJAg
zEmG3N5sfFvhMleWL+4ND5K4bQhn2OfV0zfzuc7g9MCXUPuKU736x/4K0Nx76sJj
0QLtGIXXtLM2Uc72AZoi4HIUOxKAtscWhpMHt35wCP1k02cKHRv7tefgSTb5r/CN
oOGpnd1xc4nlOt0iI292jnJ0x24IUWInhN2wl0ao/HqByE6BQSZIUFEf0nmvOU7R
LwMHW7kWzkU+FnAmSjZ9j0KZPds9W0ywBPJWtqnhGr68ozRJYg7OaRlXZ/CUzHVu
GK4X/Uuiq+AWKTj2RJboFafXJk/ijDhNwKsQb1P4e3vm3DUClGB4pnXrys+sQwnH
uizfzNZlTFrAOV8lBKkxdCBn7tDbPk4nONqUU/MZrUsb1DJ6dB6/rLRyP+XBADAR
GRoRmTywOYBU+0JbUVVS0T+aBCO8mTNhiXcByQESoqDsAkNIkXGiiP1g2OYgITpG
RghCm8ONCainSTOvM10pvRJF0ryGzQFDwXu4EFi/xSm+fQJVN+Ql1tpkTdIHf9OX
QjVk/Onocx7O6WEcJubP6bZMLH1UtQz2POFjlwUIWOyBDQp/GycK0KJ889wr78dl
5C5PV7BBwjx8tXWnfHx5d7GxeO/onO0Uo1wXlwOCs6OFw8+EFEiqVMCx455fs875
IKPkXROGf6fDv8G6o/8FqRLJ9UtuBwy066ndwdySIipZ66RWciPf/eRctfgyDzx+
F8riDpSbidUAedA/TELzbvApX4kkquY1UGrpHQWXckj2P6aX/VpOQ2YdKVOl4L48
Fwn8457xVXrwPQqS59RsMorPd6Zae8i1oHOZe0d5PmS/jonrHjaNyJ2E3avQrL63
5OpzXkjT8pNkCiJ7o2agyOlcjHgRpy0xK/MVsn4hujKq8wKS9R81nwe+19JXlMhO
MYVokCRGXRR/RAy/BZudTxpkPXqJWnBvbeZRvAvbsCpWBRn4f3YyZ2Ta+ASa7P4m
0Ze8QTsmOAS/IhcABF424bEV3XL141xSCoDU+70Huf8R7OiwvZy2pbZaDYXOc3wr
4m77HfXa1IPN8mVYfnStMkvEy6/YqQJCUo9XWYixyLoGNp5a8+9wA2DDaBK2ucrX
IQKLKhZMnhnFHvGuMPrN4SVJA+BhFgKUgKyPIMSB4jLNdW71YkSVcsRIUgbulzli
hUAxJ7dTKKdDFII2oEN/yUF9oHE2lJFeB6W6idjKf3vzpRLoIbb4x0Qq+5NEOTuu
l2PZKbQtMMGzEddKxhoAKMSUPVwSSkJG6m74Q5TEALSFkU27p4otJEFQqmk69gMn
VWqSfQoX4MR192v3gdhF54kAlSSP/U74rDdYftTOCkWeWpQlog+Frsb3OCBtf37O
uYxe0C9aM6WfoIQjq87s9M3bIsek0iObY0cmpIZw7O2C0Kp1UOV+ZtvI3xO480c4
7/9clKxfFSkSCv56CoDsQZAn3SuuBbBdMQlCWvTAD1PN9qC8IOt5pkP6lL97H1HF
1N1bSkrAj8/nBOnAHXGQcXUAxYN56e6R9EFUkdl1gdtU/fpTk/KC35NZK9wl0wLp
+HbTKZPr1y/93yAt5ORQt+AQ5UttTuAlnijnBPkzT08mqG4Mo5sQVy8KZuAlm7qz
0xxtHZqQL6zk2nVGzrUfYjLnwCZsyfGt0yYKO2tDPguQq3C4942TWm9TLbNqBGC5
4xW8bvt4bhgQiQZNQretBlG2cQimrRCpd3lt93KalO00/AqSsMITA3FKsXDT4G3A
nqpRqNXjaNlqxAYzJlvdW49SqQsVqOA0RFOLYHGM75NZ4kIB6tkZVnkfiY06Zdtx
zwPl+FuYI+BDbYoRLYprLDIKtNGYJ7Ez9yG8NOakISGI5ka+Lh4kFbNfNH2H6kQ6
EOB8q/UeY0w6OhToBkCYkd1K8i/wTpZ2Lc9mlLStQf0tQpWJXFMDaeVPR9vNw65l
KFfgtsY06suLVuTyHjCBGT0hj65LAoqJ7BpzC+ADI21jM2KlVXo0nA+LVc3CUVT0
DzEDHmEmmpONzOe03oPMWl6yUD5hUMNT/beZGWkbr30nutNjDfgPoYyvNr73IvPG
rXdMMG/Ijr4XJzXKZgrZYeeCyRCMI5M9NfwzNIUfmx9c2/vZt2g7vYtULGlmdF7N
z2KJKvW9MhSXOMNsvYsrwyn3G80PcBm4WOZAYE3fHwhleaxHBAgmk/6Cf8y5tnDd
V2qU0z4inpScYCDZCsldaUvML3kDjBEgMyW2yeqxMV440eG3u0NSG4QMnV4Y9e9p
ra/auOFpdgBfCbwypaV2D1poTsalPmAb5TIWurl/5VOu+OA+iQOVlt9eM8GTRoLD
cp85C6AG35lIePNnFPHw4InMcc13dKthP50Lqe0NvvNSSYXtyGCsKq5iPDyd5PrZ
OoQXVlxjvg9+dpv3fpYZl4b7t3TMw7G6pj76d1VuxiDNBkwsfotPu2iZnNB4OMzE
pkm+6QSnhvrGdsA3n/eW/H1vhluvqdjrtXX8pK0L7qXF7zFCNnep+aKjT+6YQwJP
vV8fTDhGUdw0ILLqJiipiC8mgnMQt5Plna9uwgyVhqbdzUFhjfxzX/5uqBL/qh4I
4d2+67btjXUe+/GTcpOEKoh9RJPAKXumfQj5gp0By+yeTtnwB1rsIiNItDLx+iC4
ZMiV4178N8FglNuzyQGfaNayNWUrxJM3r2MW5FXulqi41lMuG3RqUuHU+N+wvfLi
4vrN0tYJIOJxM+feZtPr4eGKgwUdaUProNGWHIs2pulgaj3ZyPyrUWLc4sAWz/Pc
XXEmjcU55F/f9DtrK2+uLfklU9jP7IMyimMfvZ2xjrJDF/TmzeYJZXkg/xVXjMvM
IITomTdtZSpxluwYKqbJBmiWSwGacopkVUu32rWwDpldsgiTJu22m2uyNqmFi6pI
RyHsuqGhHcnzuJntzeif6eMVxRTbSFu8pIgNkD1UbN+jTXHxuDmR0auONZfPLt5a
BKGG2hqiw0Hm63PlGMY6y8QNtUdKhdkg+2WX4qnu2XXRu4OyE+FHU0GWKUmtdfQL
KpnbZivMnvrS/FnsCuu7uPCVV+wXTBRXETObYT6o1QAeWcIIfp6yTA+Q5dQpZA47
Q0rkgJnmuovEKWmagop/47HgGulZ0kVtyIGWDtcFJRKTDWYL6SStKULCRZQeSGT7
NIjfR5lHCyeVaSbaASA3zoqJ2BzRZ4k8XpC628vr/ZS/n87MXfunFx+AK8O+yCm/
8D0uWzRrKE6rat1BHeXF2kbY9TRBMRETH93zEiBhb5r376BzaXCmNs3uUp8JugXI
USPtFCZTlZj++DZwWON6gVGO9XLVNPGb9RiW5caCEUjMU82hukutGto7qUNh5yco
Sq1/2GfWgKGGcubpj60ixgWwZT7f7lnXNtEdO/jEA8dbZj3oFo/Xfw2RZVzq3ffW
oU2KRg/OaUyOke4Oo1J/RdMxUszuvny5exHLY0WVgE+z9N5g2YCOM05o86Ng/SVp
eAc5PqY4ejOHX4qN7oEta1dtxiTBjEpKldUWqAB6zx3nTkDyWP6E1+T+GDXV5gN5
AmspRnaMc0yD7TkjcomQLaBKMWOPgcqGzRUYev3Em+ySoFEQfzZ1SHmKT2km9007
RHXIyEv3HuuW407oVHXxA6xM0YzOjRDJtu3iQ9Rav3gG/DwrPb5uOVnILrLQ0Us+
KK4IBEtfKA9OjnNrjo9h8/32sfFHwdOO6jNmnDo8k6tU3/8VPyXJdflh87wuF4l4
p/c/gzo1jBRfPwf8tO9GZHq4JVxxXgRYSDp39/GqFDxt+2J47ryf3mhdpoGWyF6L
QEnYyVew1jb5W+ZbY9LGJPm8OZXOcLZlhWoXg/jpPpPpNFi0C1AcBcM1g4BwH7nl
LsduJ3lCFey4BIU+h3RJOWIaQlEgzCkD4tUhRoics5ivEc4W6vm47E5EtjHuQT3Z
yaU2iYNGo66N/TwEFgDt3UnoUT0JbtE0sw7d81BBwspTRTahV+b2Rn9ktD04RQ9G
ZetKyqR/ZaKb0TQqpjQ3AHhhoDjMKjd5QElgtIW4KXbH0MU/WVdEaHE2LrpUzzjF
lGy3oAuLKjAN7MqoMKjmO1jiK6pt+/uy6sI39K+l3ZowaD/Xg1oN5F9blcnC5gAb
p1Xyl4LPOqi81ExObltmjj1OEQFcbWQybXkrX2H7l/STvDgsPQfL7hI0MxO/qLKq
0DGao0dJRxPtLXrxOcC31DSJCWgPdCyXGa5LW2IiPwy0X/71fNqq91MkzV9LOuqf
YRBP1uFMGOWAugIaiR6rwgZgcztj9+JCDeXExhYR5IwxrQx4TWjLgMr+bi0y1LzF
8P2JW5DMkg8AA2YXYhjy9j6t5oGnlYAXQsf0ijF5LvOk9EE2ytxOSTvjz2Jghmy9
hCgvzDXbNeIFYGutb1WZkYRVe5rO/AFyqyzfE5dTQBUXTCoqdFJ2sEolnVsgT9op
7NU+kNd3AfgW6Z8Swf1rw36ztjwBQCU+d5DU3IYU8H2E+rt4LvihZNmoEFgTLrZE
jWrmnBvntHbexfJkKaIPlZV7J7VG7MJ2oxM12LY4euzAOEAxDgXCdy5DtbJqSwWj
YZ8LueRuPOwW1KyIEeswvzQof4o7gcOw4m9SBioqQG9dUjGkhoVZW85sgsO86tLf
TrPhstNLRJ2w9hSpoG8oFr/jQ+eHGC7Ztylxy612O2MkjxOGb1xApRJFXqF1G5UM
bsv0AWWT28JeKE9DR79T60RWAg1wWiJHOJPZS3JxVXeBYwZd33fhYG+AOW02/a/Y
FcuOcC6QZ2PMpFVz0eXIqXa1AhQLw09phG9Yx0xDJCItKGoEzofV49TvPA1aN3vD
LFf09cCqBV0nzn/q/kNJuyd60EJmb7zSUmZ0zsOkAv2Z8y95XR2XXNbiimFDlglU
q1HR8sLKIo9pSzKON/qLsWpLZ2JGqzBhBdjyHK+1y3GaBePjS+C6R3frBdjodkC9
BgqiZFx7oBFtb2OqhQaBqbGvo2jNdxXi4OLqozOkpsTdFn6nLEzgm9TjpOkZ9vwo
KuHx2B4Sj+nXHXIrSEBCJpuDbpd3yqx0wUXvABVB8yatagS1Lu/nGQ9FqxEby7lm
pUPjzVlBogJDV4+5mTQfNWlgcIm7RmP4vK1giDqFxPfg1VmYg8SjbVYmA0QyW7UB
uqcVwHd7ERBN8P2XBtLuL7cUcjaqIhq6+hHJunqat8yvLFUbtAoyjNArGQKkR9Rw
cTxQMzun7QHnrSKfeHupPwrYgw8RrinwechZw9PB+vfKWb9ikwyftwPHL1SkegLt
AIt5x/PXxCQ0E0fG6csImercpntjRluAReCAeIq6y/nUGwssS9+4K2svbieQpaJ+
wWghhfaHaOSbXccoCkXGsSZ4VEubmxrG8dv9WKh7iYpSLUjVrCgdRN74Q09qggSv
jCXzEboOtWw3HjbLA1N1tyx8QnVihdQX/JRH2sn/9hokBUSeeyqpTnoPQXEXcMZw
BZDn/aDrgrCPWK8GMfzwJlVTwL9zxD4j74TxP1lcMAAU0m9rHA7hhvU8+AASEUHf
Zj77krskKwHr10SH0nJ4Bx4hj4wsfBA5jFH6JoimSFNNKkMyb6USHkqSUbmO+W+G
fVoXIfCZPwgVVB3k5JTYsgf9IOXGaxWLxRsHV1/o85i2bdRbo9QnuMQ6mlQyvORc
Et0J9Gm3ip/F3ammz5BzbSXgB6ZOs0MMa9fGTnekF0TFfed8NootMw7CzGTUX4s9
KvV0Iu3vMKh4uVcBWTdIMQah5abudbjPHKD4iZ3vlx4I40TMRfupjW49GyuSk6Ce
uZQ8JPA0JE+UwK3ISN6qrkqiwHtakjYHGT3A3bL1MxbbnLdFH3qdZ7i+RcHF9928
tjGz9dpQAMmgjaggnTeA1FAUU5omfX1VbTW1AfasI1MEG/ukfk7aa1aQXOiAP+BQ
bteTf16TUHFy8jSvNkCWmhQk1AjxILoGqNLR+2LZw8jdh6f4Nkc5JHqRZOw8oeZT
kktUHLRoG0GBMeocLa0dBIOuWmjnlaIzYnWWg1WwOYS2BDxBKMzxDFRcs7HAeMg3
0XEJn6t9d2C5yyTvvgsV0GiPnMe3iS3JxUWvXQnigRfYapqSzWVSK3Czd4orwRJA
Y2adgJt54yFkccOLlSbKaU47E/5ftCDagCT8Ga/lE+irYrTjLOQnzAS89LCpYvWa
hXtJ/MKSe+nDR8zrWloOq77Q7tGmaUqcAUl6wi72SqqZbmtZ7bajQyt+giuxQ2tn
F4ECruWvGPf12n5lb/B2Y7fPdrPKAkJtUw6sa5eqHaA6cS14SUYheKYyKACVRdmr
IPGsSnqqKfp4NT2NiCr46PGDVJkh9Q+mjM/XM2zsoQqIvHFUgg/OoGwlPjEv3IPY
jd/SrDE4/AQZwX9eH7IfmYxo3J/E7odMuV5+aa9fe3Dcyh/nyNDPapn55YekQHsY
XLjQe4Gi5Dtxzj61mCkXqQUqf9nTFnAfDxcyfG7wkpcRcgHAJwYbCT5juY1AaVR+
mHNnjGEWpv4XDkvM22ysD0APMDBWg1XksGDn6hFgyXfViN1reT4UDwu/vMEGbEyo
lSaj32yud4ihFN75gv2cC2PQzynRBni2GRceUDS4awaWHolLJ+gMnMXlsOTOlHRF
r26dppuM5KeHNY8N7L9dOxcxkzYixrDR5G0jf60JApIqYdTJRp1Uld7cg5BkuAk0
VOlFbFueIkNLmIlw7nibtrlTpV7geXJsdxqMP93W2TB33sydEanf8uDRSjR0P2kF
xZhrR4X7kTzygL3nby1RiWH7nGYIHspz6dTchxRVj7hJ/0u1/4ZcNPi1EgJ7jCV7
Hd9JCY23/p8gCWm5afUawBFhNO4vp4skp2X51vEae+aT6sJpL9IhrFbPBW+8l6/Q
hNpBJDLZ0JNyioHptSzLl6zMT7jTsodId9cF0ibzWo1Mcr6zk6xlyz9/67cVqjnT
NNaLEmnE1TTzBK4yNhKXEFdd/0mWPPcAr4oI4bwws1lkzJwztBQVQMGszIKusw2X
Jzf30rOKV+L77MTiN7VAcjQB70mAUdg0S/KtAgl0Yq8tX6+k9uNgPE47MO5rWju1
PQzoyOyEIpPUaPQYA5DG//J1qQqkvFqFWkDZJOE+EQz2pWbNsag53qVK78izck2c
15ENwDGmpjdJLQN4+6X7QyvLWaDFl9BKi/LoyPg7iRCU8txeoyaLPAqs/pURo3W8
x2zgioGbbkNNltn7cSczj3aN1pNmDKGUXtmPPwQShj7y65yJE7XAzOcnyRgCWELN
br3fnRbzk8DA86+99gr4nld625tgf93pVfysH9CCTcXNRD+StQwPyh2Y1ahtbtEo
Q57IZIvQsxeMz7Gx+aTPprXr2o/ItdiJtEiQ369Nwofi1daOVXC/GTF0gyzUkWWe
0y+pMCS4MP/vtOuMDE/0nxJjJxfAca6CxMzqhatKc1I8oz5qdP6Qj8EBuBu2kVMk
IPozou0syQWFA0hIfKohtQ4lCn5u2QpJPYKSJernMWU6rojYQL2XVE3xZKq3G0g1
yZGYZaP3OISyD+udLlPdHaEnlVgNVukMHo2Qiav4cS3z3ML5Ia7oBjTXrqR2hpqq
yzsq615WmCP2v+9JLiiP3KCjmQKtotAO6rbijb4MBbDVzNWUJXig1gnwKlpkdsYy
9MP8brRR2Zt6+J2UGUPhrdK+pzJ2NWeSLrib8G0+MylOCt7Kt4IcF0cBGPrpvpWn
3SiK9MVlaQem1GyOMl8db0fCulrgabL0nsKIfYyo7UjRN2Xf7djcXkQk/oyaQsVX
M/qO3OEs/iRr4Rx/vFSWRTLxxPvikz1JvcUS/JBVk6y++cbCa+IHMG4M4eEopqxm
61YrNkgzxy3frqRydm39Vx7wUGGLoVY5RYhpGp8Rxdf4KjfMmmnXgXV1aV0qNXmZ
KzFRLKOCCq1SBQhIweclzj3n8y+SC4/QCfoTq/za1B2uPvyQinFsbTzhfeNYSuzI
Oh8H/NBmoWQy25mdNnvWB85whAGS2+LYY5f4iFk/BZ1qYv9JLYo0uDguNH/t6MBf
7Xa+E53SoDXfbac5C88LNsdCR0nv5Vx+DQUNHD5VQdQ7oIyWOgg6e97giSJg239N
rXIa4AJKjMCP2AeeCWhyOE5zns6jCAMoSIYIUsNIeK2rVx9KNvVOGmZ8eP765t0i
GqBfbX1AjFNvr1Ee27vJdGfym5dLpdWOMTV3goLbSp1GBminQn8mSe3aUn3c+QUR
wuVj3gd64ZSQTC/ltCneIcWvFmtqp4BZ8fG+uVZkaAqohi54QfktQVf2ZnjZb8GQ
Y8343AQZDxSdAluWKfC9zrbRZIDjmM3+0gOZV5q/UMqmH8bv01Tz3sFEo53vPJFJ
ZrhyisyiYMHeBssuvvKaMW8Sns/wI91INEGGdStYtbS+P4zRX0A3zZIiZjQBbq0S
Gm1XlbAAc9oCDgNDQywue2GFbUTIg4vGGQuoKyJ1lx5w3FdPwftEJk+ZZiCR7MPl
xNBq/aCz52metC1SpDDYZzU7NZ2BZEr2SaQng5TxWlNfKIYsLK0B9Oqc9at8YIOj
T00+8DqRVB4Ofz9+YazR8VJfWcHVXfRA64VP5DlHZJw4u+GZ8QMCROMesvtt2y1v
eg0frYD04jK4/ABAsZRORtrl6wr7j2WAaLNwKtdeHF27sKQrseRSeYeTRqVuc1ux
ccn/vIo2OI+SnhYkPaUnMHg38ynR13DDHSBJI28au56gpAhMUNwyHILPnKvze/OB
V41etNJbCp/C08D8qMYZCSdYnLkbGAmWjyqTSGYXcEkFhBwfpMpz8DV8L2C3LSHY
KnGay0ns82QEOln2LBK1X740zofNR5oJyRhmU6/s11HxJUF7IMJ6VYx387ikaKpV
K2I/kvovknoerF0hJL3LLwFh07PZ9DAiwIw2dp7rFni8ycdNssqDX1k/cF60iYVS
NLB3EQUFzXrFMqyxEQ2KuJ281yeYvSgBiDsM4oq0tkp/PWWZ7ZxixsgCX6+b8t6h
rOwR6GIR6QcxEM7lIVW2FVbjrFGmIi1XG7ZIuxkf79gwWJ2ohb85NZqmgTM1CelH
opUrk6tALBhUc3C4qAZqOEpwTr4SXEuqbHg/04yTobfK5knAN7tvBI6Cf1mwXiio
mir5ylXQFCJwdQQvGFstKiPdmWw21MADJffSdXgkeGF4+0W8cNs1mw0Pz5kckk6c
eiLfuag/pL4UmwXpUUIGSsVL93kka2zolBMQYllh5mxknUCdldiTH/IV7nZSYeSy
Sk839ZIZi8oFAJ6Wq9VN0lCHSLLe0ce6SSXiJkvo5abXIomx3VuVvUDiMp8p4mO+
8ThrhcsJ7+nzYDkoN96ZAC8WeObBQ/RzwIDOkRcKI5ewP323U+lXX/kHgnzNDzPd
pyMcEx1wCD5r2n3nt7yi8Rln/kN6dr0iUmUI1VsXU4XKbQAP2txiFl4u4yTe1Vbe
CDIIO3gjPRqxfEm068pbGw4YzcjjETwaYBhPUBnjH9IK+8h95sSIy3ZBgDDSn8Qn
jeDVNGBikZxy8pw1iyrJJ3+vVIYPFWQodFUC+9r65XbDJsufuzY9MZ7JmoQN+qIw
hWIdxCqP2vOHmqseW2SlQywu3hKiUkuTHMzjnVgafau6CVsIgGVIPZ535Ihn3IaI
ZOqeT0UhtZJvwJWbsvLGtp+etZLs3nnEqmbkAFSarpfXrlJDgFVB4S3/K3AmuzUf
0iJ5xlWQHAAwzi+ZTRyQmKN8erj/h9QYBBONHSR4NML7HcCR4A+E+jtEjEIi9Ayx
a2ltvAMfR1kHJCwZWMdnSIBCjlyO9df8AS6oCkKj4eE5+qH58nYrEtoC3sE1nvbR
s4i0lv4QUr7OtkGxE7F0hIxmUyyJTtiNDzN1RGduUi++3euv0KmNgsmvSfiJCIOw
hCO/ZDbTQWybosAhrbjJFrRUWbyeGORwR80ntFsn8PDrnuCwz+vjaWha7CMDqHLW
VCsdMVR5phAyvYWwT5FymVdGTe4OkHaNwTVMIHREDuxQqGpu5oa6iShLRVvDCOzh
sIqipAdMw0RXOzWud3ctXbi82WFwThjkuCz4diwzbIH4g0V2s3MSZJZmC1MV2JtT
GRWQjETmBeZpJN5cg8OVkzo5aeFaIbPq2YF3pk7RjcHfDfPU7MlH08YHVqkhKQbN
7O+FwZDv59PyP66F/jgPKNu6eHYASS1J2JNXZknpL3/cDc8QpNPQG518KUsDjajk
OUQs54kqjAa5NQAnJHi+T1FH4uDeEXIZlodbqjb21EMuB50yOWISWDt1230rB+o7
B792eOkdpXumI/sFw5VUm9rAqE6oDjE6256nUi6PQ5VIPWqt1QdvMuv4weR/z2N4
X0e5PH/zD7XtwjEuj2iYyZdRm2+2Y8kULxgS0sj/eaY55y3PqBhryEjGLPV44TSO
FiVOTecFYcKbNbl08+xGGGQjkf6HFrZM7yPmSVxeVsVzNSG5Vj363dgpHsXt7r9m
AhDxQeaV3ZZThI3VgY5hHruZq5yf3LBtOH/ywmDTXI7FbU+G7yW0SVt0EFHOuvKW
QAq+VdmHTx2ef1ar7Mbde8j3kStytHDgMg76VNIa+g8TuN5kC8nsa0Kb1RSSXhwL
cYPP08RWtlcxH71QdtkfLjmal9S/2TxObfXMeVcQiDAdI9cvFiRcx7HKnguGgLm8
fUL2a4AkIh4Iw/1EFdplVTnqOIFKQfO4Bsng/Y3kT0UAHe0aFGOfBR6vkvpJtBTr
a7I5u5nN8tGjLboGsJHmOR5P0TuUMl0o/KO4ak/vNlVSMhFJsBFOOdw4DrOTQQLm
ZItqWtzLnpWafnaEgY+2dnHjRHMp3+bbSQ+wYxv8vkYUTCnvsE1BpzmDPwBaqxJ9
tDmSOuUtCwPl0OkZV8OdorQ0lvjocb5whvoAhpuNkp1Bxq/CVoVFkEE5RzbtMiip
4SljafYb0pQQd+thnQuiyCA2qTSBmK1iA7Hp3rx+h47EHmDlTpxZ7oRbI1Qvumh5
IzzeBUVe2Vnu2vDhd2F5twgpwAdVSNURv5CLnUunktpT3X56u7FjtwbRxdaLVMF6
yKziveuE9od6bKJ2yWWmaNXEexL3SzcyFPXsDZFfuGBnu/xj9mdIthhi96pAeGMY
rpVaDyy+BiUJ2oAgOJRuxR/Q4HA8nfcU58QVdd5KmLXaCJygYnwjiI1lqLl2VtCm
zN1CrYcPJ2ZS105cMr+i+EexdbW1DXW8+km2pa2teb7AHe/Ewd2qQ4/aNnEUaU7j
EL1WL29YcjDswO2UrcjjnFq8Ifn8fMyN17F+gmTPGuxanR51DSpaoEM0t09J+bp7
Cbl7mHl+Z2feillCZm6WAiHmM6fpzI3LCYli12ioA2HZDduEM4P35/NH3JukuldO
4ToD0lJTD8Q6JGjY4PV+sU9qZFEwONq25+rQ1BgJ3gfaonp3LyJsVi8tRAEDzKMM
5ToF5x+FKfRKO2PGL9lfTbaz+3yzZbBHWALjTsxXLMIQQn978BnOmlJHEQPlMgNR
ddBJ5QwYhppJVujN68rUG8XFc9diF/ybq2lGkMXoxTRQiOLCtf3URw6DgrD3yW1C
EYYKv8disKk6hI+1LdyoFhiiWG6lHkWV5WkLVvtwbvn85mSWTZYH9PnsBRhCcvot
Hbr5wEvplN7eywN5eO7KhUqgvE9GnPuGD1uWri9VX4bjqXVCrUlrBHOSTE6qisXk
JGtj5AS2DQ+FvsSzIgVPVogKX2ONFVGLnWjNSatrpY95FdKnYB1C7ndVqxkkGshA
3fRjuCJDZ9Dtqvzi2il7+RPziPGZFWWhNoacdR9VrKgK8+t77s23SPlyCAKQhBJY
EC7js829Gjvl0tIUNDt+zae3bqNhFgqmgRaWi3w+mpwVnHLexTqN6DEIC1KXImoL
JoCzmTKx+oeJl50c9cm8ngUsw3iEbLthC/zYGx9dNjF42A8LPF86dGRz9+ScrIra
XXkMNp0wOYhHPDvJwkz+YfiXi/efXITfT0igJcbSMSmGnt8e1GvM/PjMohHf41XS
JweKTOJ4CtZLlXV9oDe5gipQnjKNCG7G06Sc4p5MFiLYWEvWf/92zoUrXvOORAnc
2zTFmZY3RuEB1iNz1YZpssJ/sag0G08mln6jSh/U1t26DO7mqWGFKkH/WkzmW4W/
VlNT5Z7RObSv4kGprsQxO09B8s0fc0r+EjXCJigrmVHlfgR8hHXphuQ+pYjpfR75
ToC3Q8OYbY8+PyCS5PC8YRoGYR+D75Nqzdr9pjst1V/S+ChubFZbE73F2VM2Rju2
/nMam8G27KoXWlx1QMuHRtlEE31TV+JgSH6QflKYRSvxInVKWPbWbUGbGzVzBmGS
ye439HQnLOruBUHMPmkNNKWhgH9WFXZshuSYYVWAxHjEKxTd19Fz9tT0nceosIbi
HAImgAXxkWxNUDxQqzvqc2iME6EO0qdOGriTsV2OpfJA+sBg3cpWyZ2vqgpc15XH
rUs8kM4TpPJCxvDqlayuyNyAjBv6MhqYScLtReuvGy0Z7DUa+OwQxrY17u+Z/Esg
G7SaA0fEiZvSoWxhgHS6y3+2LWEp6uLFlzKGira9hh6eiknLpFjXjQgK1uadaFm8
3ukyrUEQXZ14Q8WXHGB8pJsN52yTMNRUj6DeJxQVGzlO1LHNxJ/hkbpGon0PJOmB
TFu3NMMyhqFIcwZtMenu8E6IJuF3QDX6sd0F/p7xPwZ84xf6mkaF5WNiItvGBsOT
RwgFEFZ6FC7NoEAvTHD4xFy+OHQHeBeeVfZrhmAKaybGHGYzEryTA5CwI0nlqybp
J6kGjPfSbFyy2JMj1gWV8kYXXarWVg3QOHFt6QjD2fuER7DjXBWRWKrwU9+sxiLo
URZ3ZtHAqlLZYcIDMS6eXJadoXaw/5kPVMRcU7sGBFnp6K1VwAvtXNgn+UaaZq3b
2hpNx3AwXaz4e+1RlkKIaBAt2iYLFfHlnG69PNdTAhP1k/60DTtWvpmjW79niTcM
Jy+77avL0f0LAU3kg1NyJxlmdrGXf8FbiN9GYD0kQMDfpHxgaOLsoBI9qmVEDCaf
szYSKMadn4mpqnFM2QOnXgtUk7RN6Fh0qZorhlquZAun6+FHS8LCdnN/EttBQ1iq
ci6XOc55m/V6yLyPcTWWC4nAAI5thp/ENaDLgBzrRp1HTgmA+mlesKvX6Qd2LLnQ
4lyPlugag4Ou8iQSe9cx6H04k96PlCYXxaxvqTJQk8MQ3lsCvgcXo6AEq99oS9xo
40HCFoIGLqIm5JFAyxxQptujqOkLZx9vm3FdGyVD0eDGhiBdhJSeawJCQKLIYo6/
f2Tbe4H/BnPFNL3CyV1oHWxunYJBgHdz9wIOLebMUNQH/1L0mxE3OiDO8ggJOeXu
70wvyYcgtvXDq4IAymieEqh9E9zn6fmT0eTuImQ0ZBRvjhnR71lbXfMmV69p9Tza
NHlSqI22ADtY98Jzb6hN+DOSdj5A3lvb6kSaN4BIcaYfOCdoOUDkBUOkBoro4BJd
G/ApYsRXWDueQh4Che/lo6JkckzwItt9dBJ/kGrsaB5leye8EcI5EhxH3Qj+K0ud
28gZI3H7JYFh3shfUtqTHC5Oco9HwTBAF6qCTieJgKxz2FkDWVE60ND63O7NDHVt
s4PbQaTFKwT1IxEwL7CRPwqEGp0KR7G0ezNd2QrA1s5AaIhxZcp5Zg/v00VsGzrE
ZS6if+FxHH/mkeS0MG4WBRQJfOaB8r99b/pU1c+agx2CqFpzt3fXcAisnyT1Uhf6
GZCmBDcpDZCkx/cNrw9vHFtGHHCVZZY+T19DrBYOFnjOrYegO8keQh11FSEjYcO8
OqD60eie/IaBDbKWzCiLvL10r3qZ1nZEWk+tlZ06VNCIkqapYH5vs1JzpIKOb/Rt
Ixb0ieNG5CVLAg8+fQmwMg51NqVXJ+9HeIJxYfTWT/lsChRdklB/fzva3IWuCdf9
06Rn9Pg2+vx/fnthXMn5n+z5IQAFkfVxQz4o792WCViZhP5g5yG6SzZ8V3jzr1sh
aKZOFeLbUx8M0ttYnF1Bz3e0YU9lXeo1eRsj+NIZbk4CvfiF8WzdUnpnIbnNFZZC
fmLXVM9HvIugIiZxnZWlozd9FEruCR1RO+SHXfwgZ4r199588w2RE5AKEGVgEwr6
cSke4u0UTR0YfH5pktBa7a9iz8nv9bdqPgGbaZc+9F9Pwub49SxCxRu4y2DS0z15
/Ov3iMAGSLhGkv2qjurCY5ZLpaAEwuv1wMN7kG0LjVyWkGm59aJKT0BQKTGHPH14
mgv7V1oB1P5beHB4elnVD5zjVm9dScZ2uoeWxcgoobZYavmmPVPVrGhqZRbaujjk
hCFaYNe3n78cKlyS2o/93NsFj2zTQDOCa1l/X5LwaKpx+Z8Cg2AuHrIZC+FckMbI
krY9ht8dTn2Lc+6n2yLuYKEhbuJpq8u8dXeIzPufOfBT0w6LS8E15HqiHsuC7hwE
sms4vHnX5Wtp6wOQJM2Eil9DOT6urR8aCo0SFXOmY/+Wyat3EEiGUPZIjwUBy+kC
BMyjjhyDhBZRnXDEy+OdRthvdgEylLfadBNnjBgDzjEiWO7CrmARySqQfxrx/0Er
eiKIbRNRSTYh/Hp1NgMAwgNjZXl88NE2G9MNkHMXeoPjSgmEJDtjnbf91ubz0An1
kjLTZygeH7S0BpiRy1bIfwuzgNpFcFms0VDcTAO9QPfvzhp/dC0DbIGvETCLq2Jt
IeCjbl2VDeUXHyuuRN/wUeHPr6CJfrFcXtUcqNaze9k8tbjqrGtBgDnZpC0fkub2
I2AdOwHYv4f9WRz5pawRZciFuLrLbWzAQpCRENx+u0aVM9G7UDjtvvs8FM+fzwdO
+NAaPHgIqIAYZwUfW3JRlRWNsKEHKVeL4ownvuqfgcYDSbWAkW1EezLYw3GArGvx
13iTpf5B+rk66ozfinWlSbLtOfFQ6BpcSQqnv0HCAwWv9KcoI+6ImQ2jr2SRM5Lr
5G4Q2Utf+1qHNMrJFVjIWobs7+xlfscaJk9IKBKFnzfWJn40hcxXJ/2D9AcY4UQP
v0bwm91bxRG7gwAeGUL5O2ng4dF9z5rrQ6ue9qpUVLi2Ej4khmPnSIalLjczKzMq
0zsGlNwI5kZMozVz2UQHVnvbl5PvAw+K7XUJU8jjO+2D3cQTBAT9+gRjcWGbzmiK
0Qg4yky7zPc3IF4OGH3F47xFlvxIGm82IcLv4SghXQIzwIQhcEMR3VPvzOlnLZc1
rtqr9xXy2/f4ZZxQM/Cn27Ic099+Gb4KQrAWJSjepW3Rqsjp4s/osgTeLPQsVNGZ
YX2wffmJZgbgS6Xiv2/kTdA3uursJaEqHditXID+VkdagsodlM+PzP97yEMZjY3z
o2nYbn/HMJt3OApN2F3cmi8pM4tzKXsAXWGUE8tSAIhDS/YnY+x9Ia06HN/L6Awl
dDj33CAKwOuWvl+S2XWoF1VjMlV765zHv5M1B7ud5I/ibdpQ3Ot5O39h7OxaY2oF
MCClPPJlAjwQPIgc6W1JNbmYNTgdS1d2f+a7CUOKJEDB6x6GsjXFqM1I+7KGpm3f
rWdm3eLIoQKmx0vAXncW4YgbPr2eoZNCKHdhGc6JbLq5rOlUGai03rsfqgnz5G6j
XDMHEWmC02sW8R/q6deTnoP3GeEd3iFmYSOOG+B5nsMWGZFgt2QlJ4qMdsHKzwDA
go+BUV7rxGTlh3i/TF+Ic+1wsoi9rNvsqttGoPu5eLeGgi2dy1P2duU6pQav5XEE
KyPAMGl9/9aNdxIq+GUZmWbH5esX6vVr25eJ9ITchiwTss2MYNRQ/5zUlSGycHFI
hqJaUp3To3UQpUnxVH0y/me+P3ATufSbCnM5o4zqA6pgkc+6+fXRlEFoQmqlO6xU
B6IlNfF16Q20XZaBXeCE3g3lAMZkis7w3zQwEuMkVvm/DLi47MxMkZvLqeRbjGnp
YNkw8MFczfhJdl2c4UlU1YOX5HGWL8PIwpu7tRanaLH5KLTw1SLlyvPpaqrveTcM
qy2hY4iHJvQhellFFftUYp79STO4Q6JQhtq7Mgip6rDveTHNilcfqs0zxjhSf+1l
Z8Sdsk0t9hE0+n7O81SI/Dz6Zj0z15ulJrS162uWpb4p/74Vq3dACFfYC4Ct0ie6
xUuWBR9KJeRm9AkgehNtv5Eybx3RkE9YjVlQGK2K6mzJ5cZKL/nEnQuB74HhrbcM
pNiv8CY4TYltmAh3d5AAFmmCz5DxG5qXNO4fwLfd1AmP/PUoTaT7VVrLaJ6C1A4l
5e8BjhYRixDby2tihXNGi5eIbakYjmE0l29fBqBRPS8kbUf7vUkm9J6WdgBJrgoo
hFespPHISSlBvIJjJALdatlR2cxpYXE0rvOSkuahB01nN7k3+ME22PTjn/gp5T2w
gM63vwgCsn5fRwgZBz+a8qdQmCutubiMGti7UxlTZ9wXYoCFgMppV6aDXw1jx9U0
xsb0lAHXGyHmBCfHMRxEqP+w25C/80OqnuMgzl1VqTwXydYr69MuwiQyLM0AlS30
UKleDlOZ23zxLcd9Q8B1TmUJHmH+yNzWg0/ZL62+4T65dvE29aGoPglvq/e0h6eS
zEl7fiLbrVUoG/yuidGKUQCBQT2Oew9m+/8D/v63zOidHG4oSQSjzZU4eZhUfcCn
bapHFWoVTpw+SmKSHyWuASNoWDCMFcJIU2+p2RWIyDNf5ak/s3Po/HE4WF6XDzZM
ObeRyViyJgv1l+LFnN/TxjYpVETV2Yb9shZ2TcUlCw6FU1jUKKzP6t8LJyJtC3xn
Vlbo9l/X2KyxbanA/agGibyRsaPvjJ+1SbzBMnsfuaoX/ti1hi/ynP3WWh2UPsJl
d3sLSDuvLfGzQ/7nLlNFD9DOGDFLEO1PFhrPs6UMkesR/AxQrUPqMlIhgkkD/c2O
0j/l006aEbigovbQv9A2qJIcv+xpePpjBoVumfqal84oXoH1u4rVtgHlyzD+0vnl
GuZFi93k94i7D3pHEmtzdXfDf7Q/dZDl1S9RgLm1G9NokxUS/MjYlsHeK+MIzMw1
9pSqj0UzB+4peJTc0Xifx0byabbsuw3Opcql+W7AgMNm6Yw+p53b4DMGySomMX7s
3p34pI6dt1KiPWg+qAzMinD+0gLyabkT64MrSdJUWbEmCmZgrz73c2oTV5i/HtHy
InIkImPNobkdIed0hKURbU+BUY6maWax+CFGZCgj5oMzISL6A16jyzNTlaAmIkDs
WRlm40rpHcYKvS/AkQS7Ew4M7NAVEmkQrSVxDfwlhrty5f9n88ChAJCF2EX7rc6g
YEp/eB26A5ycaeq2TD8jh+Ix2IzW4kLfmU1ep5Kvr0vujRcKJsPS8VBaIkoGj7K6
ibBgY5hJF4lsuL+Kpy7EiR9ffrJoWXnNvNkvCIYvyq821z1nvu41SObUe+LEYxVp
tOaoj5KcwTTSWEDKrXwuVMOhknvZgcEdkadxs+82Cpc2s/M2qJkmQvOly/a18hrd
3qywqvvKCDU4798gtq3fvAnik7YFyK9B+qiElMxS+IV/vpktN5U6SKXoR2FCG4tn
iOke2UhfpstOiX0vzC/UdqEplfM3uPGe2ffgw1OvFYak/8V10NK+nWQHgJf015ug
IgW+68/37OV+1xwqD/XJfAL4012MM/l+np/Yu7jvCeVttiBZ/SDx9ICtdnhBdn/2
StqsJGD9mdQmLPFfSMwQaKtWLnOIgIYDddzEVVsPftwcVFJqcz5a3hP9JTTfRIf6
k4/j2RfacHebGGKisRj/JAsO1982kRgqBn1hnaWEDoUo0YujFVZbzviFH/X33nWZ
KYkDWrxjQoRYXL9S4sYEJ8L1oyCi+smMhj9HO6TM6zja9dQKcp7sSdd4lpBLsP8R
0DUv8HrW1fK8fgK7k/Dt38dD80t+9FksYXWKm0H+VVleNxl3y6GEo1CiWg99H/8d
v7WRZHQDSFIYZTiU9JsJoliChBRKCjM8yR1qr16xigKoKKf37eYTr5SWeU+YO75i
OL8rVYiLMYRhU5F0Wy7gf/P/JhbUlSW0/CrvW59LiMiahuHySEVa8NztwIUv7L1z
KDvIu9jborKNgwJcEt/+JZCLL+nu4XTwh9kq/3DVxFnFpk3emDBxMl0MvI3K+qxw
PIUnarQVu8BNi/M/f+jwMZ0wzs4ysT9nwIJJ5EkmdW3fBOpWhgIe7wy/6Bcn4S1I
Jbh2YCywW1XBRdsm30HtvbEL0FUSe0t+JhdTpAEcnsOJK6PfHBsqy/WgrCew8GQY
OOvrffBOaCCpf1dOp6rmNEQBtAdNeCwsD8vqt30AdnJ8n/oi0Iasoypi7wOofj2C
UcuzihFP5dQyP8uT11EBbgJHxs1wkyuo/okzrFvS2tvpYJwOv1UguY5dWQyXiD3q
37mwzGd9vHdQiwlIC8LAfKlteejLTzm6B/9gBbKa8TQVxNdJdnph6SNu5T/22+Vi
+C9gm7et9Tc/T/NhzkUvUhKS/wBxFhwgBHyoeokiVYjfY31GPKldKwGFQpbpqTGR
Gz5mT+y5fcQjZtUst2fx0deM0jiCq14TAr1qEDShaN0v8pAlcBHf5voffrYmYfM9
Ixdbpd1n2EL3JB9o5Ogyirg7hWkmsidphuN/JWoO7v4fETry3uc0Es0Hu580Ghvg
cS8Yqqq3zptRfEUpFIUrJVgTdeZYDtRewuUhMBc9/4TGlloe/D45R+gQnMnvB4cw
xM8BEsnnnDiTtgr4VGwY8Ro35VURtXnVwOUmdoNXNCMn69OVCgYrVxkivd9rJu7C
vczs2IwPN24nA2tyUCKM7NptivUoZIjjgRDENMA/H/h+nKCfYJWrG9TtzYGDmzzS
18IMRnKCMCNe18GcgUYBD6U1HVsNa/ZCgD8JUnmQrHa8ewHkV4ew8n9CWwSRBdFa
khe4PuFkGt1VZ7aQG6SZiMkGX5QCG2nshT4A/rrswY4VUIrTyt/zrPBYif3t/wh1
dWLCIDS9W47f2RL2aZyAJ5wFu5T3nM34jat5hWALQkQCQ35A/ahlHPTia/mOkM5/
WyBfxxPBbR6VwyK402wO1DdGJdBRS7/30ZfYOsG0vx838bEoSV/+Ktt7VCBatArW
8E1owseh+dLi0wWPp1jodt2YMiVuyCAkl/mSRkzIxWbM0SbwtXDj2mK9w10HZijS
vqTt7OgO9OIT5Gy6/lXzEkMCm+Frk4b6x1qMOB7B9/PwDO5lYoe2+JflbSXVqkr3
8LadWXryP0L3VtjNQn3cQvOilNMif1PpPxvuyAJPJdZMVov9i7feSMa+L0UzTpdh
prhThal/al3HzRU7AlQ4aXYaxvi5l/daSfWTffj2VivPlhnpVwTnqDdEwaGkPoFH
ahUeG2snUPPBCiLqP7A+hD2wFuUEdDO48Pa2qHO01ZkZwHS5Eckyqjye8SUocHVR
rD36e9/S+n2m1yhjt+chimKRo1sCJpmdxwgmWExoJM4LRFq1gyZ6+F0Tfiz0vKzX
Eb2SHq89e0roF9nU696fIa+XoBrDfNhTw3hHFbmwvT4+jlbh2JBbpGlN7kqiAmHy
QM4PEknj68fQxU06w2b4AfD33Q1ELBEoIwKVrNJGIbKlcEPxi7erUEThzLkOS4Hs
7r3Wk94PTIDNDdraN0kAcpXfRTTYjkwvBL0Up23ooLic+mW7q6fuzU5X57B4MV6g
c4a3S3K4pJPHIR+K3YjqHWPHGLGAqScJT1k0s6efBDjgA4PODB1CwXqECva17OZb
9vPrgE5AGBZSUWmmHMI9u+jHQ7sdtTdHO3f2brYG60lqDNsBbli4ne9tdL9kpQAj
ryqL2I0OUzLEa3tVV3yOUQsvW//uRcR0DhwCPjH7sRWjXZhLInOf260ynE5bgb9h
lgcuk5dN6IyHjbUb8ERymB52PAlvtv0RTvO17yAEwkMA4JEeQxENNnBdJcbuIAY9
lAF/PLg4TeHXZgTOAI9R6kXom7tFGO9IaFucgeAx7zgCuetYco2120y6IROIFfRy
+C3GhMwwRU7vQtvOwstgbfEiASd9y7SV63pQihnEcCWuZNXtOHZDLlwaZRpPqu5J
hu275iff2+bcqh/ZW+euukHAnR2ghGikPBu9RbqvBDIyxZQH312pTIY5KAkT/GWg
s7K5avvt/ODe7ZB/+twPXaqJn2mnj0U1MmTL8sqGQ47GojewvqIdxG9qQh6inHrL
ewPQQm6IM0SHU4scoL8Mk4rcnhFTqnYGpaUr0zCv+URdXizB7QAnQJcWg6zJ+Icb
/3oAIQCGvOQcZPc5o7VOerv9mT5gTPk2kK3rpl3KfQzZcDiY/urd3gY0h3fKbPFX
8jjJWcZjQsjHB021ewDoUAN6U4t7ACgqzNCdJmk/qK8mU7wr+GmHqfCLF1qvGwTn
z91QiKg3zpjznKLOefIJVk+QIRPI1DNDHgzt/+C2cVmYmn8o80t+QWwSlgeSo5dI
Jix5DANHvHNATLu2YWNHYvOFc9Zht8IFYrNyZKB3WbZCKMitZX/k9oKe6RqBH7P4
Sysuo7kHIJALRH6lJrdo7nqH4kR9szRihhFxCodpGQ819v6u/ZxX7n2WBlp3ppbt
8b4FqP2HoFQKiTw2QqO+xoLDsvuDypGwI/qsrxg2C71b/l9DHmjE2a7bonlZu0xH
QHd9FUahbQtikWvan03qMhGCuzi0oSJLhrn2CLJOOcocB6rrKZjoVSOtSVtHyvz9
RzlLNLv1mo2HXvn//FXD3tnNsGlN8iRnDG0pjEchpOjR/fZw0SCwtFMk/TxvCZsc
LJHrXjivd48UqUIk/Eal5N+NJqDC2VPpJN6sWfF85rhvGLUmIt3gzAbptxl3GJO5
B5V2QCfN75VfRAk+TPkAcba6xghS2tXCQJREAlhLUyDY0JK9j7HHaADOGeMwEo4n
O9cXopCamjntP7v/cdwXHB4D0rSX1I2euIgFc+cTr7pRnGDRbGgb2ZA5k1naDBsB
HixUmAYRNdX1tPxNDxHIDq0bZ8nyGcHdFi9MqgpmyC00X/ri9nbddkh8TgNXlgXh
58UeuoNXHRJ1rUPPK7QKqy7vrOUHw2P4vyQCyMYoiDpE2xd0FallTUDsk2T02ITV
0RfrBfA2+76uv3MOSFEehGsfNa3lS+SfJWXdpLmZ4i36laQawfTat6wBa6kSvFbd
9OVdSIqwVRAET5xhWw7s5deVsxt8y90JriR2kumJgRvrc3XdT3NBOLkKe5h54BRu
/u0BapnNS+74hO5KawYCry80WyG55P0biS/I2m+j3I1pcDJ8NkElMCMV+sVUAq+1
DuNPkRszr0nYOga+GlLwrO2GupggOiPBFT82erov0nrvh3zF96bPxaQJCVma0G/z
eLTTBY1s/TIgJwf9kUBBqrRLJ179YrVK8iR8AzQWv3hMQMf3koaz2QCDRawMhO68
CKzXid25BwxT4XOjwG04zpziziinqWxlFr9MwCWoqnPcp3MoVDACXpcdxmV+4IzE
Kho1xqljiVCzKwCL3RTo1UmuepeEplqe9Cb7k5D+ibf8iDfWzRxq44q0dF8fAnTc
4d8nkh/rxpKsCWcwJgzf0Qa0PMp+VHdMXfHU+vuSlsvssbaLa3vEYbhRdScwUEMb
U1mlxtnbFXPPsWQTBkeNCnq3whJGVjqCRsRWQSfCNwGLuLQPcm4rSpgKD21SjjJQ
HL7kNJXkS4iX0+VB3N3bttjQi7JVMEsphpkG8o2OjS1H3gCJ2/C1t2ZE8WyGKACn
6VvBIDDZ6WNJ6KU8f7zARG4dENsrt/jok/ggQEa0OdG7ZfFe0weMCTub4RNeE//l
ILcjlhP4LFTVSG4tJgUsgjGOnooHVlj4bAI3mUCzrJ+sf8W1h8u1nzHDnUKrv9X9
nVI2N5f46+3PoYMLM5r/ag3LDx3i7G+nPgsrjj0DmQZ0qRrku95PQG5rdL7QRD47
LwTEmX7T6brqqmcMWyrS57t6DgbJLAZpeuNHT5MPkijMYUo4A+3PPrlAOzpx0/Nk
YiDk8YjjyF3VwjkPiMXwpwfWjJKBCbhKSgJHB4eU8L9YrAwqEp2SDmTTYMpAwxlX
8CXh04jfDqZdyJ+fWMf4rJI4UQqKnJNTTB9jOTDIaKRUga/CKhc4RuKa2wv2NwGi
pRmwbbXS2d3ClZdWOoqGINHSiTNaJXdAFD54tplyQFydHnvUPlG66V7QFQNv02Je
6JslfMiwtwN/uESC+WzF7EqdqqWYMh4sZ2xRRIuu922HLkWlrPWxH0Ws1feNnyw4
XGJvtvQNdn+O2NxCMbDzw7UnQHxD14edebqGt4AC7qyN+bkNdua9mdnCQTHPfVDa
7Xp2qnjnGDgTRnnrKBDLgqZIfyV9XhvZHk3n00y/GtBI+XxcIpNK6YVQrHj5m0dP
zUb7xhZeRUo3Jh51p1GJG74VGK8/te3bldBRWK/gp6ZkJJ93bAd9IEe3UbEogAyb
E7ex4GodMaoiaSNl6kRzkvFRxq1yKYdMkro1NQ/eHSzYhFZS+ZIh4UWBTJ7m/EE9
KvqZZkw4SnHDwHh5m1w8Y6g86cV9r6dMh4rHD7Nc+91RXq/u/uTf2KA2/lbsuJGJ
jixfFPbRiEOThgNtZKpf2IKjeniLnu2I5zxDu72Tm1r2wR3mWUYkSGdXPQWwifqu
1zyvBONKq2BbhGvSHjVmQ60IOsD47hKp7jpoecPgSzHKkOwrkTwidGAxvSvZGRIa
WCLE8WU+v8fbecdIaAaKqsthX23JmuNlyRed1T5ly59Ecwf4HT99fw5zQgpHsGar
wK9eDFHK3PpvnNQwNyTBieDJugIKtLA1q0oMekrAjqrEts5M1RxL+hgcwQ2JMSwq
yelwDZLy7eYzxa9JKqafw1DOeVZRtr8Zd/e6xvv3BuZVlZZmaT5l2DQU7FkmkP4d
WPGli+JxCP49jB049sRiII7ogZEobqVtDQKNPqoqfuyTf8NBIU5ttwzGtlRQYAq5
zJ4GAkUcwtZeqStij+BLHdMOfL3o5TQirIZsZFu40BFDpJUz5pmdVAMfGbiwzOVC
BivK4XmnULAD4RKiK6HvgBPmYxxF6QRAOKsy8VVsNwRxEF5C1BVSvH0PVs0BiJyp
mr1MsEZsTY6kqkH+NOKcGUgQsCM5k4Z6EpiLhgDgw1IdcJmy+mmm8p/o3bUZJj5p
dyTmj9A4+4nJcjv2T0pPr2gpEEHdMK9aYnGQLKMeYFDvuUoINvnAs9vmJ5TouTPP
Rv6Zv7c1QGSm2yupe9NGZ8aL9BTS4DZwfRYDq7hku7RorJ/ya3/BBOj91T4qUcb5
4DA/RoRgBjKIAoEf+GPg0+Xq6DrW15+b+9WAHmqfdTEmNpUIZT98iTo1M8Uag9Vg
ZRhBRPjuhMNVIOadJTuIIaLyC0NLdRKpr5ZEzKl6r5iJnQP6akC+cUsflpRIwIA/
Z2re352uWhrZUKqSvYPXfYMdGpihA5Y79M4jg7qsmdNwvPOszjwB6FnDU6Kg9z7T
OPzF0KBmdGILt7dkXzwXvAwc1xGk+IlUsSg9zTbNOvkPe3Psw1aWudj53OZwU5Ff
aknbSHdqlhQMJu1XUmxe7vkNkkbrO8SxhHLFyiuZ89oDyglpICrvaIa9O/6wo6RP
SUrLr+XgHPWfgBqP/iB/dQRE2ujXl5zj92OTjGA8LnqP0sxSg7jmd7Q1UoAb1Bo7
pxqo4bcSEIgQ8gAncLCURtPpy2baYteOLUB8hhfVWJo1Wfx7ElW08+omlEan8qYN
RE30+JiQOAGsCCyDeVe8M8E46UbX3pvJO5GnFn2U7YRaGq4l9ufYipYB4L7ndqYO
ymDAnCOy/II5n2OarShwVRdp0rhnX7BRpgl1XRkcVyJSyiAvTlskkOdAfuXFs4Eu
ae7gk+zsozu7HiS+GPggKTIhbwPVoVBdDIrtQDHorlLDgX4/mfuarTeIOn815XNE
OVOCflCSc07OEM0mp2aCzogWkrHSP+tFU6iN5Vxm6whtzOqZvoJ+n4roIxBf+GPg
qMv9hcDa/nxKBE5DWRAR6ZuO8CZmcfCbquyXIXUSjpMCCvwRg68Ujsj+drXLa9w6
lD/NdB2PhjHT6MELEW6eJtVID9iZUOeEkcLdGY9cw8aAz602M2rdHe2FgqNbm/6j
vtxx73PDu9x6rdQ5+kcP3ubmo6s0l7+eMAWMAUuEVBtQZ5DHD7OSztnLMhO0q70g
y5DwV5OOX/1WaxGNwdhBhhuZllGDxGMGGg/XlwoeKI4yJ8AoDU4y1us2FxcdLZw8
uzv4qKMnyGUz1tH6jf0+8nyQ8efr6LNRu/7LwKas5SvwmzuATQKN2JSpH8UgALvT
n8/AX5aiOL5d8LDjtBViClKdIk22gLzD1idcWBJ0AFu0FzQOI67jeovRfVZNhMUH
DTsrtDT1PWgKfvbfMATn2wm+q7zMVT616gmvKh4LNqxzvZpXG3uE8eTdSN9LUdmZ
PinovBBiWwRXbi/RX5Z+Gsjr3HWopxMFYfli6KesfD7vseq3iSZmsMvu0+mvzgR5
firFkekWvIuH4NYkmE95xe/qu5O2x6OLSOJg/riIU0UBSEm3IiyeIohhO2tHqvjf
IL3xyp+GPjZtMKW1qw8b0U+fY9uIwi5cfJU2OlnjaHEWAkRu4cWI4CaaFr+OdkxL
NjM+ziYzkh4mlaQXDg5FM5qhlzlRe97ez0g0BzlYh4BEFJ4GbHvAoj/paDt164dB
wlwB7TtKt2rgKlZg6RiVVyTbe2tpCJLrsupHzaex/Olb7rHW0zqljd4a5Y0qCZHN
h5gwhQoH7UlKzHQubkkjjpnHAYlvF4k5IG74EkL+0sUr1ZmbWoeHy1B/GyP/jLcz
v+OiJvUqh1QFzGKc1hBZY7ePETcnIjBZTwKxEuWvlokVXCUY7Wz4OE3/bKrbv6GH
JCoUCV4T15bvr83sirfUFWurlLLQGXms7P5g6J0bURMbu7GyA3AWOl3tYVBShJmn
Bw8KX2hkTqqsMD6gdaK9mEKt2o9rd9TONFNpupH9RpGabhMHKzYEbIVDLftohdfT
Qg71a7mBzRItZrtBhrK1W+gCym4hvGAY44dEhh+ptsVFNlV2fKDXKUFysGGsZyI+
TCplSgxl37755+WddhmqOEISO+A10O8zVaRotdCGmEiYFf+k+l9Rpuck2xGQ6gvy
JWY6ihOahWTykeXxbEDI2zZS6qov5nN2iDUImmkKAIQ86FBN9I79W324QE6LKelP
cMKMeHFygn9OVBqilF11bgMEjY87dUmJQckP1I/YAvKrsAwRN2yuejgunvy9HCe9
xgH5iq1jO2WiLz5Sr2prxJTR5YLKDihWq8V59bzHzBO32EQwjyCaNIRc1GdtAARG
Y0ArFf1ZwuX0N+lwPQo3+8s/E1JSdUGo5SsIPgnEBcCvjVbG5/FlguRpNx5nR+6w
G1Y3Or+HmBAF1sHujIAVtr1jMUJZiK3p9GhfT0/A044YYhmVkm2Ag4gsXk5hld+V
HMDRTN6KvGjoGEVMH9P5oOnd/ORWZXEaM6xQ5TQ+o1V/tZZtF+okxOri5gw9MQHi
GJ9rUIZG++hT2IMirhtjM78pV+DT3Xcd++pjE3lyC8/c3bts9SQO8cyFFkb7oUPn
ITsFPN5LGO8Wti8TAhWvHIMtvgFqElOuTXSzO/sWhZWz3wNscooC6huf+ExMlaRp
L8OLzpE/O6LJaq4bgDNe5A000U0Ckm/MoSwpn4QRB71wnyn9fg7OHhbMxSxeHZ6C
4jkt/R588XKxJ1po9JiprU1tWVBIhMWmLNy40ARHC5OuApytejiCh271g6FcegUC
lfm6i0kVf62/LK4500xu9GiUIxamQoVWTUyRrJHTv+d0bKgQJxPfaHfGUMOcpMJ8
4ps+uaBt/zhFwxL3XVAg9QWxrsj9gO0H3xC1VEv6EAIfuBF+C7UTZANSQxpigF5/
2ktvX1/R0K9RM2ZnjnJK0xjHiwBNACu65hIvKCD/KfiEcLj6ERlE8+8yh8GnjLt8
Kk4F1qwP97E9fb6rOZKBR1SAY7OY4c7sfvgCOd3P4sliYMS7AHJoQUBzgD54QXnR
slemqTmHZCoDFhYKz0+v22n4iGReI4MAtCQBrApAr+oeEhKNwNFuUiY/S8a8qQEO
9ciTaNiK7z+PdsXANUFKS4m6O+LwIUtlyrXcnww/cLXWXd0pDvw3vGcjvaU+C+OR
apMf1evd/PmbMX7XoRV7EqJExK696lQcesqS/UQzOtarX6i+Vt3cNILWpRhcw35M
nmTg2xN8DDXPQhsSkz82YDPF0Z8onCdLkPt7lmWmDhoMv/eQ3Rm1nx0BP9mbNhOH
k+E0qcNfBVtPd/jYsW4pu2DAnKUM05Br23LZ8s2ZVQY4nyzVLeqUCnigowgt2yrh
UURySj21HvCHDx9e/5QSeXYGIYD7bQMHpAabw7DEno3Hmyx+rZ32bV0sa05lbrAO
Y/Lm/vXmuY2QM2AuOmLS6vY/8zVMHwf6sRcxgY7oSUpKWPE/xjg1eKnaWRbjAbT0
pGs7gXimGb+h9QRB2FkWIkQXjPPAGNpLD52XuvUApfoqPZh75rsckUxr4UUeI1Aj
DJivJnoCjl8PjY42AAt7EX6D2CbSq4JxKP4+CX7APomOnxJ0Xt+i2XFbFufN3BH8
MfRooxwbATn3C8VSCFIcCS689vUlRiCxHv8DCIh0t2rkIkziyRKYkKFArPEPPy4w
abz2XuA0eiGFTvIt9VJUdGuNVbDML2cvbLZJHA/RvEfL6hs4a9QgkdGSE5s49Xj3
QlJEoo0hbtAxbzT+nIF2aGMQpRfftVHAablulswL5dF1zvksSQg9ZFU1zxg8rJY2
W69JW2023I9fVxYPt2sToS+H8WUzaVkdVIufXzK80gr00gSYKzwTgsNhOkz3Zq+o
LjbjDlNTXyLoGJ6R2asJsWTIIjDS8so/nGcmGibafbXYYbO8xKf3aPBi2WgN/0sE
usLAgI6mScuOMwH9M6/6S6jkVV8QHPa/q5YkLnKR+PQKmdjFStcO0wPfoOKuBQRm
46k2/RJfBo2pnkN8jAEaIXAQj4n2hIHnz5TImj0YaaXOD5qEDrow38BFkaIGe6Wl
uWwjVBoHV3O+YeAcBtmHM5SifhNSiLUe4zvEGoltE30SS8d8hGVoxOfQFy7L4leq
TQnIThvbR6FLEcggg1BscMn6evqdXiTr47CnnK09g8ULHbWkYju9s/dnenRZcY1V
dajhubegVA+x2NLB+sa8emzrqRIIBkWGEOyzbObANTDgCY5hdmPcBGHsC5ZGxjG6
+BoR3VDEWVfRV3xFOgz55pkTvumsFkP4KTJ+wdP4d31wakmw7sQjqmKlSmkRHuvr
H1ouDczuxrAqf95D4C+VMhShf5ak0OBoENHMY0aJ7wnuB1tiJOta3r8yDdkOeY0x
YSAQowKU3jdYg0lTnxvtjqWOUmBAPVfowCEhApFZGZME/+WM3v86W4/TkOgcvmLT
6bj619JAnw+GfSwNx7jMM0B5PJpBMeNLsLgPySt8LUn9GOgN3oy12bCr7aOuGvE+
Wbl0Ze1BQhuzlx+hgGDtSy3KYH4YvMpfeZKd6LQJamBpKzX8cMcj/60JMrqrxecY
iRnaaGN/QNev25dZC1OLS5sTXMk3NYYAAUoI7pVgqyuakPIXoxtcJ3Qa0BGdOl46
nr6CoPzZUAwK4ZgYw/H8WX2+/mj3m4A+PiA8/Yjjjf0CjDhqF1YF9KPcGXNHTGv8
aH8DbpgR9auAR3k1E3DeLfniZB413mBou/VZ8FjoWwNyDAgbmz8JlocY7Hi9C+QI
HsFCPjjHhrtyCJixi58hv6hUq9ipJuBeGd+He6R8lGjJXTYRchjHSy0uSwNlfwUD
cJCT9FuGRYwtTc1rYkIFS5XLhDcKhmNeaRDygjaSaotrB7ukzK8JldK0VxrYyFp/
30Q6nNfa0nIwJaeddjwaCGjglNVdUCsq817PT+8FqFkuMKjv4i8WVr3NseyGh1+6
zxwwWnlW6CM2wXjyU8iuWit3eBmXnRlTn9LM2G0Tim1xu7pVWu0R/ZraORsGxMi/
wYLOPO+0i8G1tESkT/xd9hcarnbG0xVLJ0Pk0rqrwTMJAiCfITg1/4DPCQCLzIyd
/RPbo15428BTUuMMuCZUEdUQ5CbaLeJAn8ASqGchRUEJa65evAJY6+cjPTbXea2h
KnALk7hKK5pOuJAPbOGpyffBTWLCWboDyp/Ez9NF/70R8a6iwnH96jOxQMZOwxYy
OJXsFO10P1s7Gv83PqYYgecWrMFUU/k0apEdUSh9+Xw0DtDOZLFtYHA5Xb14s+TZ
iQgDesLQAaNKffY38TPVdq/MfaEqTZ3avm+NMw3lGCjHvUgevcZAd7Q8eow1WYp8
ad+ley+w9ETEqA3u0WueM3jlqVzravTmes/QJY/Z8lxZOcToifJowKNxsQULpEBb
IRig/LEXutX77qONmprehgKkFS8FZaQT4CRhrDpYgr9o5jK3Iu9zpHmv2ZgyAkF/
8zJn3CamTqii147zRSIxRv3ga7zMcs+QXaRAKUS9XPqFmd3qxxCboL+sNw3jGReF
Kr4fl6cDNwTFtaXXT9cAcoBmQe/BUIs5SBbZDc6yrDaJpEDDMyzXDFQr1CYHmW1U
JO32STvmD5hE8sm5u7Bh11kuJxUUeJEhvdpaVaqcgMmrPHbNqtAKQy6jTcoC/YSH
ppLFfY4/+aIpExZLZAVb2bdsGp94Z9Cm4L11WNntIH2FllE4JnzePjS8I2jDAL43
9a+ntRgadUXCwGk1Ofz0ZnxwcQXsjPTI+xVPdD+w7Y2X9LAPda7LhA7VogrYIGR+
SJLQQD+ICkUGzy7lDYP02U8Ls0UrUYZm7TrRlBplG34HSn7GFxHLSgdV+uhiUIFb
+qxF5oxyN9HGDVz2g34EmTPCLZYZKVBjsKMqy8vNBQDpqbJHfHbQbyg6bVBngB27
Z2JTtNWUvHPlt7URD4bifG+LzsXQ3krZ+wtdFtoi+CEN15+tcsJz9zXwF4wryrKO
Uxlz/sEky9Os9r6C+XujoTuhsTprZIXv5/IPWqTfT2Xgt3lMbiueTIDrZBCu6dNz
T0vhGnfzmXjlW2wFqKtL5wRGnpII++1aeTYvfH2xnKsWoZJppxm2WOJIhc2OGZyZ
5JFC6NiiwXZJ8X82BaJH3zW/sjzwXHHdLN8JEwZuJ/yZ+M3ggtQ/sxyziUJmrSaq
rKBp8j9gmVC1sUJGP5G8oltfWv8kYkxphHqytr/H9dM19YMsff3v8b42QUp5ogOY
mOF5rRokdFXBRin3CJRSLqzsGa7JMIH1X96qYyxgKCD8MAfAIfLWIvK/d8jSJxHH
0Q7qdBkzBHlIaChyhLAZF0NhE5/FSzvMFojDZPSOOCgGxPCCltalVrpnHnhcRj9r
+lN8YtBQq4nbGzn/mI41Nm82bQyNZs0wqMG5nLJxT+i+4wMTjqix4Xmm2uhG6512
kQ5x5rHo3jR7ifM++uf7dowipqhsH165W5HztkdArZ46NzcCA14Z3MBGnBW7nx8h
o5HmSXAuEN3sFePqppCo4HpRPZgJp2xxNjHQOQ7bg4gVW+oxpsjGlTG1RFk7pUxL
/kwmsS3V3phBcVMGUJz92etfukh2RakovFBXKuQkn8OMW7yU2NZCSmb713BOgMIe
iAMyYpw753/EOT0JJStC7c5A1OuHK5ql3iwragnin0u6wdigmt5JoGOVwArEQT9c
5J0Vh88lPFwIaYMOSJJeLQ0awpYqM5mhOfTZW+O2z8eyBFUR4bP/siuzTY/zG40Q
qzK72yzoon4gOt5xFsnc03bmiDbP+R+aXh4EtM/bRpRwqWeAOROPUiDOLjE5vkRD
kEh4T6Wyiqil5VXORDL71vATBIEweu3cPFO9RF4/X8O5wThHqgTsXbb3xyxpzMiL
K1me/hOr683e5k4KyhqP2gLHIYkORW6BZl2CS5aWCc9WRlpmPSx1Lzmm2YJPSZIJ
Dq79fen3XOfSQrk2RdTQWgwHvAsC3xyZPgs434eMUfMNUvjn9lL/Cj/EMKSsHgvs
iEKpCtiDzgo43VLCHFW4DzklhKxtGdtns1+v0sJnrm2zFmqjdEmGbZKRqs5U985D
BxCPU6j8t91zwYZavNgBI+x8FCRZa4aNQeFOgHckyi3fX3S7B8sQDPrAPNneX4WX
5b/U71UEzRr+wxMh1LXRmqwQZsvQ+wD2vCbRWIU6bMXakh3K67Zyl0Q4N+brkjxz
XCd+pFejBacRdz6lromwB5gTghn1jNYBWA0rcrAm+yz0DP4XSpSvvY0mQb8iNJ7a
y4/njWnlrEVlZiDNSuDKUZ6n+D80Eq1sxS61FJfYMIHouBaROUOzc18AR0rdF50L
PT2uyACW5Q1IdqYX5sXJUj4ER/1MTEfUcTB/3DnJoSYOjr4BPW/alPnKgEXFJF7W
Hf5dQcl8ogYViAfX+vpn8ZxSOPVmIlbLx275mzYBhLNL+nIrgpqJYM8sQf5C4Mj4
d5GWVqRULUti8Zh/xSaGVVrdWJ5CVeigHEMfCK2ykiVUtJ8/e59uJZ1dS8W2bKtS
CGJVP8f92r32M44fw4WWhfYkYxSos+etff0+EPwXqvroQilZ+NMGem9saxlPJto4
nof/SopgV9WCA2n6l++cXv0aJ4C5lcZknM9zhdnqBCIi9RVUR7xZ8yFe1UprPKSn
SmxONJQfod03WFgDFld3e62SJ0cyaAS8w9WFUHEH47fsXrPLxUk5/NzymRz9nNL7
DtO1+0vVQgDvEz5ZGUaN69iCjfQ+TsDrFeBgQwW0/aoTJkQw6nAOJ71SUPuegOhV
dIlisL9RVEGN+ER9aVMJghDa6bWZJkaC15HvIDYzpweKmUdgPSMovS2DuPbwbquC
WMQygqT/LGNJ09mWd0/P04qtia9Ix21bXa1/oiiSq51FbhRS7A+b/kESkHD8NJIW
U58CfKkxNpBhLo1cVK8ehK70GClrkvxhIwy7o0se/gztA7Nw9SgDtbmPs5B7/Voe
mHogKvjWYyI0GFJCYow4EKajS4BWAPc6cmONfjQcuRhInrUSqKWUVTQu3Wp5fyuS
PZB5w39TlD6qzqSVAqEsgqXyHsU+R2qr9aTBNK2Pv9g9d2QRFU/buTlOm/9fO/lf
nfyV/oMP3SfVYw1nkVZyluwZlvybSzE2h9OHdKcRpYrW0XfEj9rN50v3Cd5pLT4S
B+IoDDmSooos4f7i8LoFos5VG9/yE6wJ3hdORECtieK2F6f3z3oijl6rtp1RFBz9
qoRWADeiwnixXiaw8b5YVR8Z631e/4ONhuknG4A0NTM395CuWfMcHLCooxKCewn/
xVJofx1yGF331pzJa3yjJM6vdu4//U2iw0GZcImyqcGYzzVTSL1FrrMCckb8Jsns
J2lYRM09eSyuUZ62NKqphblOpxuDH2Y2egwIuDspKyj2wJIa7ODICoHBGy+12LV4
40KajCvtjkey4g1PjoBpZfWjIeLG/+pFWV0ScLxypl7OLVKUJ/M7Fs2qpQkO9Wke
l6LzAyikAQ/TrkKrlBVjpLROiCfLWzU5fwWwAEKMXQRtEIp964XGylws2QTXukkH
mWMqsIsZbgZ3lkFsb/Qyypedauxq2JWpdtiDbiqonmszrChHPQSYitRfF2eVQT33
Sra/RxuOrvBygkWa8RYt0vQFgjaoxKPdHUnSC1JfVOnvsOnsMfGWLfmnIg4p8oEz
Dhg+ieMlCmT7zzfV5fLtUY2PLayLAhhu+noQzmhCdoNlNavzhAQdoDFqw7v3rPm6
s+Gh9kExcGgMHAX9Cg8LiSc62C7v95zO2hOqaVZIxQ3DHOIvDDTuZdFNrwgv6HjU
WQ1Pr4v68lYgLxhd9i89eT52+DSscSWim5kDX8kP56EkbJ92In0gqo0pd0u2n0WH
41QAsvj2NyXY2GD04IZecpPrtms0RDhXILYAbQrQruIKQdb41EBhm6tpc1TZ7N4b
ZS03PfG7J/TaCu2MXx++nmkZ6WVyUczPLgS2T4aBUmKvbqDvl4vxtVCcZLQH43j4
W6j3y+LKFid69wXQvzPqekrCDgB8r84KUNzJO6t5r4Eq2RwF3kj/KcHO9LVZaze8
D8kERVEFIFh2JOtcn2EsdQ6eEi3rYEulow8ObgrLxSYYysf0frKaVQVTN9ApIi+8
gfOMMjybOH3jpbsBt28cc35uM79K/KC2yF2k3OJULTb9U9n/A8NUQd5tJtBcgHJT
PWnryzRtQUwHJk1sk9b5P98ZoCE/QFBXrQzhttC7irTBD0I9mwIapon3atkICdzO
rFviYz9HuSAr4zBKQgPN+1ZI5YL8Is5RBcwY4RIBkSDU15J3AVDFvRK2J67dLF0o
Ha0Gu7gu1Dgz2uOu/ullBNHLCCatnH+XlhmYLzIblfXytImQJB2O1x0/3WSQbFsd
HGv1uJVYrICtMb7ZRQK5JFvmFiU4UL7LdVpqrigFdUr78diPkZEh/i/zWo6b6Jkd
AuQp+umqiov9uysWE03K2//+xxfPpmuPEJV8WfLxawYKxmsw5Bsor1Dsrv1rCJGz
ypI7HcmhKESlmPnUSwk5RJucHBjzGpgzZe+ZO+XTeX9s6mj22lYHAxQYAM1zTzys
1TZmubk6W49MFF/S4ZiglUfPuzh7bDqPWLnIpq0QdSDdfPGOgB4ml/gUpwWagtVu
rnOdGYlVlrEYslQg2yWF+2mudq4+g2KedOBj/bX4vMZOByOowjLDkcRmsYa21vPD
mDxfSA8Vn4Gy+aWQ7EjobUbgHewGRLHaUwZY+VYJ3w/vBOaagyrPbBAjUG8gU0mm
Hvs/DPagv2ivNB67o8gkfW8FmayLGZB0UE6i/a/KcnffFezfYP+ubz5bIwYGDeN7
TYo92Y/FrLnRhuvMV5m3JxF5dLVBqEGuX2IVko2ED+hXlN9xabiGjVpqdAGnHBfN
6nZr/7HrcNKcHp0zbJjBLMMcirur/OTtO/UqGm1Kkd34G0pxXrkeI8cduRlZWN6J
BHtviQHrz4u0M95kyZBOKMGFogU3xok7eooqSDXFX5eVQTf6IzS9jkuEmeZXR8Il
S0kB84bq5F/Pqdsf9mzHXFo8VLYweeZnVXyh9eVnmHFKR6nm/fp4Xg3ftfIdaKWz
RtI2y5XrdmHbc6JQsvvZlbsZcfVG4s3/zCgTNZJ4XnzfRBvj6Py0/CIWdKsWZm4/
3Pa0WfvVzPJTbRHiVA2QaOVeUIsCik9F75g6xaHrnqKdb9pbgGH3qfEuxS+1GkDn
E1eEjuDRQkbiepNcydY0mjY5GLE/Ec5AOnzK03dp+oSZqFC/j3clqSMtyd4sPANm
3oruUoPEMtaV8yalzPxBZBCGaEJhBRzAwm73+HXoPmRdSJYiiFQAdaoQZlJWVWaT
LvJKz3krUSw0n/RHwYE9Sm5RdpYUndqGtlEucTUVdz/tUad7OgCtMOTGNiyynG8x
B5WlJaSsHJKgUbSp1H7CPlS6Fq4hR7ouCrotBCXOOIAlgjcZS5W6/soP47VNswz3
n6+NB3rk5rlC5l2+/jIwCQuBCFCraA2mi64FQxHts9Yl87FQoZYHBK4bKhUIyAOM
IdpVWp7hweGjzG7AKmjNud0ih6s8+RxDWfr4zp3msA31Cx5loEfXL86H5Y/9irQl
NESLO/4MrsCh56WJu9iRbV4c1Tzl7tFovM1UMIxQQS20xbjGaPAkVofaGToFAXd2
hOfmU9e8yOW3S7yxfxGXa0YElUV9tfbq/O4Os/Mq66Occfx0V9d03l6w3lCW4fSz
zy7+qq9I2D8d67LbuPyvViBTK9jrhXSLbDpgdcAAEFj2kt3TJnCo3J5Qz4knl3pW
AvRaRHuxBIpiFIgeU7vLgjkgTPWrCaL+Z223pehG5KZBGG1/Xyva69198FryVzM4
NRXROF32d37HrEfaKpnoaBLNtj6XB7XlCH8TMH+WH7P76tWipIdWQSDe2wuNHE2Z
j7l9kBuKYpDVelkTjQBlaA/xYIhPPI0O9/8CZTH4xGfocGbQNodApP0y0r4jbU8v
UznD9b+MrHorkgemHb15oMZ+A551hCjQNvc06w85GnGIG5P4Hidqvz/KTs+kTBT4
Ic8BHWobsVKm6qxmyi3YlUUDQx2Y2UMGy7m40J0luohRUslixMAugqUECWPf0epi
pRvfIPu61xApY5/LA7712e/YxV0aILL0+G17I2YUvGXozXlRUgstBjnm1rSfaJEE
Td9pcfAvxi83x5iQZNdhddu2ozoGwAgYxDkgm8Jovg3joCR1ZsCEzHm0FpYrQ77R
+y3GUYbN+/uOefgHPyryNxV8hcUiCqrPMufi6TAgMUILvaYlS6HlPGZp60hsPXW3
1QVE71Lgjp9xenpk52Pj1vklK0AadGZ9GZ6YmE3eoLpeN/fqJ4ejHqXFYlhC5qq5
6NET1GX6tylyZCywywhYRSL0Q7rFhsqLJswBAASIeqNqHMw+rHMjT2cEFNHDHcpJ
tT2vgRU90w+Awy84ObwcEcM2MMpsNKVToUk1dgqycW8ajQZ50rwMYrIxdnjHgjQP
VIVjxwpskz2FpqXrvlxNpVJwGzeb5eNff0Bhxdg9A1s02TXtxIE/sA8+KPiB1SPi
9LV5ROsAjsUvp3v5fUy6MBqlLRN6lv9+ZaclkGBx/i1s2R2MDuITK1dDuucwQ5df
XHDx6yz7j7joYv9lCmC/VXUyfioLg3pqyUz7bkLh5KBpxwcYBJTgPsQRyK9gBmUQ
ezF2norGQ7Isf5u0ujXEfbGYwEAQHFEMNyrxiONmJqRQ+yXsEpqT9G2SsDP/KUYx
X1HtUILFEMVV5uXP5OmL41oMffuP1csJkNnpmIrZtiNuHskCEBjFrg/zzKoKNk2Z
p0SFB+tbcpm237SnOOkimwbVUpApaGV6kVkiRp+LNnElWbD8BwYTAe00p1t31pbM
v65Hb2wu8JbALvvH8JQC2udUN157qqaQQGbPUkNwSJxWmwjQgkM7oNbrjxqH01qX
oDoIpCTVZG7zh7Iep5Kovooy+POKt4CmQICbu1CkNwmp97wsuaVwYlskxJYys2Nm
CRVffQAWeN5/aka/6cDOZfYrtB2xonnYIKM50IQ3XCd7772wsKD/wZrStbhAGamz
FHN+Usl63up2N9cmF/BWMK9lv9yWMt/45iaRjHh7C6AutxRGUf69WHZtXTqVMTld
D9dlFbvlB7QGLRAsU1i7D4GXRvVSsqANwkRNDwsqrY6z3nnR53GdKvrAAlbGccsT
g4qAjTmqly5d7XKBaTnVoEyqcF+47pKOE3MxXz8U0DGZasjzj3NgVBORkzdC63dG
314emQaWPY2MgHDTIOgR/Ca3E+IKE9NHrnAWM0+LLPeLSOJyC2Xm4fO+5PUCtOO2
i4o02FHhjU1Ha0UrnLSIH5fbLYR1wKICCMma7WRYbxmAoUbsF+Q4H0zMH7p8ynsh
bzz+LdgjjAMe8YQSMFCShiGhrPRG/A9VhMS7c13r/i3cYldM7lzWH//Iy+ogLm99
ihW7QxACwAMbYcfNqWXuz2kXnIJ05V4CwpbcOiJsbkuB6S4YmlPz7ISd+wWMA8sX
/GmYLHS3QsZq8pY15uNvSyyAHaWTApuEz5zxUXKrqXqVATWnkRc8kBCBCj/Q0JeA
he+7944m3QQLCfvD4PeOuZMEptwdpohJLNFf4UeVOUKJNR7a/ZFeKb5iJdbVti0w
gS1GXoigLqvy0X1Jy+JGBV72oN7IalSSmlT6z8dr6mEx4myYLW6DPwcdBzY6VXbF
X/R/o+Msy5Wsb0tde3q+FLHnvAIwa2IaumQBkf3j45J18k78m7xRZI9KH8WRH8RO
+9Nz3zIkSLYU/ksnOB3yxKbPDo4cr9J+PyhKwQnhgU8DHvK7QbsSB+L4q7t7xibS
ILFgLGfYKXaE9LovoBG6BfupnH3GufBgD4QxSBWqEmZX9nyCat+LST7hZbzamdRh
+OzDtpV+Ckw7lWFxlHCoBi6QKIP/MeIRVSX8Y+eri4ymOihzzwvQk+jeKRQRunQy
388KLxHBOkbKBejVK/7CmS+3DJJbrmBFCzqKWLn88U3okVsKurzfOlniBxoU15uJ
BY8g763ki3MdDT7ulgm9HlFgd5iM9CoNMLRSCsn5sQXNAAabodnp+qKHn0+pmqx4
k+6T7Jd01JB4m2tSesJW/OR4Ok5PFRZtZbRhMteDqNdiOFPSafWU2RMRHbGa/boP
EelMi9TQU4Qskf0LbqMFywGgHLlMIBDAVSv/aU/OVMyaTDj2xZqr8555+Z+EnD0s
AeXS5b6xmjZPd5fWepKSFzKJx1y/sm7eUI7IVpVyMfj7c2BXg5dRKFxUrfiHsF8C
pd1rdYW4HsLwDGSDRZFouQccrh2WlKcWpXP3nHMd1ZSdq+U+TwX58Q9T8APyED/g
vvSARjHapXY5i4Pfzg7sPqnSGyK7ksT+IHErUSRAtnxYn3Q5DP+usl3YnEiXuGOE
N8clFbDVBawSDrR3sj38pp0ZIkgfT4gmm4DEMwFebWEtJUVw2V8AZUsjWp+hU45t
m0cOGxiU1Pv6cP7G5kodge4NAmsMi6gAby2rhqk654jUn86AwW6thLRycQj+LLSl
NHJN41or7h7Yqjzp9K27vjSIDuQda6ap0mrFZJY8+lCW5V8UatqSHPVurN43o2bo
UN82WJWOm4RHAeClR8oBX4GfR2P0FxzgoyLlLb1KoSfISoDn6g8o+8ah5z4O4pLL
p+5gmaaRfWMe6l7i1jCDLULJu+S72pTWVmv/yXyaoWxxIZKyoPRYJU3xA03vxtjc
+1cikuIqEJ/yi3s7WIUi4EfsYoyL6Ihwl5vONlGyRuz07kMcEQoz541CSX99CGN3
+f8qcISb4oXTLrJjNjCVo2xIVO0aE4L97EJB40V2RtDmty0fpw4fHKjdtlfOQqHB
tc2dPcyKLi4qS1L8bzKK11A6zFXemt46QVLkvIwcxdb+6cXDF3wVvHwXQKjo9ylz
UmT5bUcd9mvuEwsgMyCJb3aRhr2KlRceuVpsQZWh+mVYwM5IJnJojocOHOruaIAJ
uOsVXRhWp7PqKRuhoN5JyxJPZqW0gQeaOb4vTIAa3udYbSBOq+X/f3+B869bpJhc
GS/krrzmys+dCLWWQpu+n+v8paKZlYRfA2cKQr9/FFDg5D+5NNJB66Lm1i42gIEy
dQfqwCj1FAgLBdjSkmOkVtdg4x7j+kpWU5yknsGWOlsPUUBx2weZKzU6ERGZQ0jZ
uc+e2TQBfmCw4ZC9z5RNtoX3aLlRpKakQ9I29Fqci2vdECe2dJh4O6huACSohxsJ
hMLV+bCwaiVC7jQXgIHMNeV2YjMqfpCJTIzlWvcTV9qnZZ++hZGMyff0clFGe3v6
tNXezmP285OVKJb6rN/GkVRSdNC7cF7KfrimvcCsEwEI1Qmg0Iss1h56l44VR6WI
/F8oEWWsTsf8Od1eDZN1lzuYwD+AR9HBtwcQagpuAwOFtTGJ58MC8ebV/f7T5mqc
qwEElDG0Deomi+X3XR+ZC+OmrJBFb5eGUd2NXJURfNuo+ie/F2WVuAIKtIPmW06K
Sh4MBL8wElzi/271UBkFIz+cAWi/1MtX2fO5s5uTdo47XjzV/D4dJ1NtuPlntbtj
f8kkm5F6ZRdiMy8fZGPs4iIdljwyT3YpIahI78MVYo42JFHQwJAbuL108qR6T0iT
RiP0nJMgzYgJxofAJQy9JhkwIlxI6/0j41BGkXjpSWS7Ujx3iv5fQyfQ8LQ/vmRi
UFt5gZD+RXPWmqTZOKGNVdfB7f1sqZgo4S4ABoG1jDJCsK3Awhtvq/KLCOHH+3GU
f5tMAUjMNaTFbMGMdTilW+tplH+o743TsEwaw2pulaCIKJMTJuWbgYlGYBWx/41V
FHwSorbzaqLnjKi9O2wKonVFIWe93UpFp2+fLFb1CUxU42xdmKsRYl1zXE3HTK9N
Xj9H19RDxQpg9os6OBAoOl/bZWQFM4FVub0LOsmAMjYoNqayq5W4hhRMNG+JWcBF
d1ZVKi4Q6R/LX20DDnzr9zI73r+03iz05sSZxYtcdUJgXNRaoiNwEacVIb9inx5V
arMWENnoUi5ACJDBXaTuzOIanwx18nxbBsBeLt98avALVoZRi3KzfEdtNDULy7QC
9tK+8XPCN2cGor1Sqcr1H97z3+JBzPoxRr/Hg8w7PplyhulPgnL75NgSTWf9Hime
EILY5ugJYTh+CnE6xwl2Wtc7kdmOv9xFN8t3hqSDyhd6fbC7kjktFRJWwCUNqoEm
gmbu6USxz3Enss8dIdu6+yemp2cDkNs6cvfaSxS/oH5WcAYtfic5OOF8uNcXoQr8
ER/43co7zP004boc+AnyRUgwh2DjDR/DImnDoMBISgJ+s6nDdAuB21QRpIXOk4TG
GNm8fRUxMvMLbYupz+D6Wnyh/6zweN+60vMEqraG6FekmomGVO+3JGrdanh32GMl
ANtfdGHHNky5ybRb5ZwdareYgM83jOd75tcqod/hvW/nkGnAl5aAm5+D+pe7vqKh
G8jgoabxiOh2hlba8FqG9Cj/smmfyEeocpOvoaaSk4LA7EnVDLsd+iIe3k79N/7v
eYlv4VkCp+ZAJ/znE+hkHiSYexnYbwjWFJCZVFuUeKx4MXsbD+Yo8m+ONKGS421U
bmGfUzOAIATle7R6w2M0vODFoiSLPe/WjD9LETKk4h7YQ2JEtUGB1NYXAjsGVXHo
dXgQajuklf0gPdbrxxEMXt5nWUFi2GMrw5WKK+eJ0/RzS8x7A3hIQO+s02Sm2rkt
obC35GwOCQgotQTlsTfRLvUKKLCRDOlUn/0ImV9bcRj6bEHWhwxCFofxg85pLYP6
2E3QgUWr2+mYdOD2od4qrcxN4sa8uc39eya5mgu2LY/MG5cX9Eht7Fg1/F8D2GvB
8rxrP3bBrbCYxaqO65/QUitVEhoYnd5nRk8gFxEzO1DM3EYop4dG/YYMF+BjpS+5
4hPVrgtLn+rc9QVWwRxY5Iw9SHYq8bkDD6WwORqO0cZD1JJ+l+ncg6P/erTD0iWD
QOYtEXv1LbSjIqcDtBb/LMnChWRdFSKyFLYjeOB9IdZScevR6i01FS/WYxgAJ2nD
ov8fTpx9rnVOlDGHgE965qbIG5Qzp44X0qD6cV+xUIeiClEtnz5re9/QZpvMNab9
QVAC4L3hRekR+49JLPfP72IDj9DYrtNu3ldBJrTApjbbS3moCgDjHURStbuUvyrs
fbRQHftPbbkxNIYJFdwgjh2BZOnvA42599iDnUwtVFKesfsVF+aRt2RQuvyrpLwh
ofcWzH4cBdLHdv+QU6gaUb4xGK5EdM+KA2QLwxMwXMbt4GQoBV2FY9FK6T08IoPM
yDHEz4OO0uTrICY4LrMX4vaQ/sVjoU+ykgl+ocrzezTW4AwNNWlwsI6v4zO1obk4
KqpOCMN5F5mSpHx1N8N2mRF4s7jAes7VJgWtRY2kUV5G3/C1lT4UN9ZXOFryp1jx
wrRFcBC+vxd755ciTQ8riHaDxTdb3nAYwDMQqehk4IdhXM+qcnYHaT3w8FitjxNb
JErCs6l1uRHxrtga82WW8roonPRKmCzgiz3UNimlLkcQ/w7JzCtwQeHDNoLTMgQc
8hKc1rL2sXqh1oIyQB1WbVZVayiolA6TXMSY/7HoQ6ggCX36zuZghps2AKtTDkDq
zfm4mj6YW2MwKYul/mEXDlZTsAEYmkKVsNBOhF+Cvj3oqjnJkFiJvnLTiOwCTd9+
ZNETrPihyMUinuerFR3n/Dkir4joIfSjgj6f7Ix/FoZxAMih3K5+9TIF1gxyAUad
LlsxqTa6s+Oq+xoUcglNU42nrkz1m+Wwj7WMV2QVsIoEww+gJ9N88NkgvGB9613n
MgMcYanN5Mqdwgl07OVYph+ODE+VmmwP/TSkck8g2By952Bhi7crbUJ1Y2gXroDS
48Q4j0epwvLWYXcoxnUOXNw3EhYkPjWI52a5jskn3qdWqevPCdwMhT7pemx9ebLy
zU1nWY5XVC99TH5oUGuq0c1vQPk0R15xwwmDuwOAUGW4Tr+TFbOpnDNhlVt05KZp
gRBpfocFQt4GBpD941SjL2O1SLWC2q672Y03Z+v74W0zwYIbNGrJbBL9GwxVzk9p
f02dCGhsdQ6hKBldMZ80gNacviTVnM6dMYKFqQMXt2/zLLT/nGDezVe16F83jeqC
By52HRGNN4U6t9ip25bNSLyMnDhiT0DVGv7jChmic7x1GphzQ1NqcgpxCVshW7s4
OqMQ2PsR4JYUOlV7TPTPlnrOB/XmfRyK+AyjKbljxaGTam4I3p5x40hatdQ5HTWH
jGZlpsLIhfLhTxb+T4v1skFb+rRUZyBw9SuA2seDV51REFnkCZNgfBq4rjIHjSNR
iyUwT+apOJggAdG+AF18qzmi4uyMQl4YwH4u1cAHQTxSJJNbZPlz/dV6zb4A4Y+8
krXVS9HxGixMR6yfn8JKVYZbak+ZU0qmKy+ZDZnhtdJRNclV/nXxjP6KK0jg/vBM
44UwhcPpjfTjsCMHWf8iHU8vL7txaRrDipg1iLBhq5poHfFwA5nBwwnKyHNisJgV
dLEtzP61eAT/SnSrTqXYWwC+TIvdtBPw/qqGH1YCWCDFZuTD6HlYSdKYFrzVy2Ng
tMD05ti/sLkvu+mATgvjJ/lnsrjSeJImcPfRvhjZ5ugGBHynEZXSqyiEqoENLbaR
77VxAyA0/m7K5F1CfthcE8AiVWSWSfP5rvAqQ6/D6XpBzhNukRHlryShXwzJbPUB
LLuNO7TrAvxqS8z6wEgTlBr4wWjXZaRoEsv4dQbrUZtJbzFnPfS1JMJ4OF73Z4wS
dVJFHpjSJ3CE/2HT7tPxB/HCXI/CQBQWYjmHH0mn54cQ70NXzAJBBXrHGpIrAZvU
/xfgmUqLT5LmwKdLsl+IBV9ovUpNNxvk98O214Rxhct0mkAGEcfuiW+hRK8XvXqf
FBHM5uV/BrzFFT5aJyM8uPwqtJpaKMD8JkI1a47yjHMbsrG6zmwwmWxc8VGkckf0
z2QxwAWg2w+nbCjWo1Qw7me4BRVubnVupjvFZH33p7b6uWDB8JrIYBJJG1w8RcPS
wMhBtY0lF+Ao9LsBNq75cpZe3GY8D1Ru+mgS4iR9jF9Idlz8doY6H5DJn43dnWyj
0zmOI0/sPcbozCF+o3GAuE23yLktVRTPgEDVcD2Zu6RftkDtszTZTQayC8TJ3VrB
G7ZurltLQc2wZaT9MnEZCjIPR45bJwWE3ILSMYIKYTXfpsX5AbHBaPhH6U0raOad
Gu6HwQyMg9SbFYrnwOp+3LB3OnoUD9zSk+0XCe4o8WCv10M5kKL5cpUBsGM0WNpy
VBFBs/aT2JrJFmL/xhIpna3S3InsTrNesq8CDOk0RLI0ZnQEAEV6D63xuNasSxmU
PtnbdeWcMgqul1RqczSkqid9U4xVDHK/hzLg7qlQk55wn8azVr5C5lga+D8RJOQE
eYXUNcLIOpJg9w2uaNp4lt9Dw4vNg9wxBmEa51E4xbwRfLhGgOsngmpiBd1h3M1r
6Y1RYye2sJI891mH7FUnF6HZ9488LqZmgu4KRXHig62D3xUK6eLzboj6OTZ9e71N
GamTNs0fT9Ml2qL2zOiwlsfirGWmAbhb52WZqZw67qj2xWn6Mo+m376U4o0aVj+C
zegXH0MI+AON4kBHIMOOB8UN2XtZ7JtuRlblNvI0Hqg/Dt8mmrVkEzrXyTIpcXMD
euZKGZeAVyO+bc9lKmXDa0ZUl7Y9tplzJsW1JDL8jix3qnDbEW4Yblh7UiDuboNJ
WBiaHljdLb51QNR6p3viHGcLtKRHSaV9VuqDvnOZd4g0f5b5kjxRiCMHoImmp4aU
v4Ww2cjIQsimbeOZfMtRiA+38tgdW0FXCtZsFq7UOi5oxWay60tG36cpSvToz4eK
MPxIGRfTq/+Ecz0zehvG9kX4PgV86D4HlpQSNBkePCxGNll2rp3HIwCpfhLAYcEc
Uh38u5bHTLG9y0yzquFNQw/wZg49UeVutL/GTrvC82ycWZInI1RqSg8zBevnKtGy
VmfwQ6Is6+qL4Igckzj5OmRGkKly52fLfAHiTF1pJ7CcmLA44TlGwx0u09mn27LT
UQHlyb7gcG5tLqvEQ432peMV/L6alssS+MmD879kfri+PHGAIM/jFO6t/BojlHlK
3cgU4dGsTw4RQDwpTw7m9HRaYNWyzqTV8/1n1jB2n5zMhmCFwA3EMlcPAQv5msTF
dAis2VAKfHIEJc6cKhXLfZ57jz09BSgjW+lOmJO5XNhwr+2FiYDhLbdzg8dvmLeM
a1Vx9nMHzciEnOH7GgK4tHm86Cf6u9b8zvXUt7fsmMARlSjWEvcCd5P3YhkV0PhL
hKPdmq8KBRzGX1ADr8081cnEsIVT9oVHEKqtq401djoJ/ZbNzR2X9O9eRv+RNlwk
koWeh4gWNQU/92MEr56yUYAz6WLEXeGzWuzNA6oUOwWOWKOvg2nSC7pvPR1i+18V
ulVJSXX7TTKudFYB6zKq8ujPuG7b01K7mvl805YtNPqemYgEBAzf8Nl7kJL7Qa0F
dFBh2AYx7fGz6TT26rA3jghcVSKM9bySwB/sIeItqvRL57sZVIthIcHHew3bl2zk
iLPns8+R3ZvN6N4AHTxelDD618MU6nh2QyihmgBu8xf0tdCDjjNT9u9CxzU+tNC7
BeGBI4LVavRPRzb5UZWJv2q3FTMdniVumFmdW3WRwgV0YmBxoSF7rscC5ZCJ0MBC
5AgFVnuaUDMlnDn11jJ5F9BRmDVlwLCzNbX4I8pqAClm+6h/h4eGis/qNmSs9HKG
Qk/IldEVe0w7E/WyBfLWEBpksfiFHDfqgWFCI00hJEOq5THoAWr2JDXr+ktBmE1X
pYfVPqZVsPhsT/z5OGJRDFrIUL82e+y7ucO+puSwNvb+nEfC3twEd6t3ZUh4c3Sr
L3N2J7LHpRYZQO4y0VlSczsb3VUzLJbgVHpd1AGwHxE99T/JZBjWmTwjTrFDO2k9
qTeMGuhB0VFCTaxdxoZJfVMOxFBNq+MARLnuLnjzFLTo2RtX5R9mZeVUD4BQquAt
SUtsdpAdmY1evoaKGdZ61Kyk5ckkfINY4eBHlvUSaRdD768TfYMDx+AVHUCtBdSl
meu4wCzHnpUk9z0HapuOkesAApX/GhSIMf/wgBQ3ZIwboOJO8G6jlpP73TR91Uld
7JIjXMiFvldLFR8daiINsTlKurlfsgJrDP/pHKkBe0hU0xjFGhM7qtT6I9xNIVni
FHg4ObrGVYNpvPydZW8q+5dCmWF8cl5TRQX0aqPXeapRxQ208fgse8EptGAzhTMb
m4SiHpigJbKp126PCic6VCqCB0q705CnUeHCt7mQrC7UD1E52LWdr0X+jM+CxElK
fjfi2SxRMVMzTIMs3GmKGhRgMoJ3hPp6U3XBDeAjS/FetcYgW4nBOo0JC7txx1si
YaBsNIr7kq8qfo5GCh8XPA8RlVpATYasWKK8kJS2tw3rq+mn9X9ZTFaE39aqCL8i
T/7F68qCLUSwcKK/Zqe8O0PrSoDWHwvzgpFDWI52KcSlNQbd1ZvQVX7QqSJv//OI
d1BL4pJRJW9si2FCq4uUdE+uBY1oq/LqXH0n5Quj9bi+6+krGiCM4leSM5B3+l0J
9X++0hJEY9Jvuu0rV9PL+aW3NALepkzTmQCSMiIec74PkFRw3awGBbfOit1Kte8C
scHOEpRWAuV5Ws4khV5/os86WJl7txMryd3rYqjlXJgvrFNXgLrZVjByg8rorTNG
CjBZNDOL/MX3smBHfk26a0g4BObOD6bR9uc4KxhSjfCH3BCvgzUSDvyPu7AfIP2h
pFf91xj4IcKIDKAouF0Q95hDFCwIS62zRjoxqkuILV9hliYkUAnB9YEpXSUTnS4s
GyTPsqcZ6kRJJEHb9a+m0aMgv6n1Ovok40fjlsaQRnCtuB2dfoJW//OAD6RY7sSa
AkP1aiiU9f3R0TpWx9AB2H4/H2zCQ2NF/OyZKhoM33a2cLoLv+V3e14Wx3IpZMBn
QJ5CsFX/Wcz+c7mJqIr7zL1hP0HbHDeoOukcIiOC8ZSRwkk1uvh5Rn6mRFCutLA0
Wy96iHtvfT8vJSOPbZy3VnpWH5MTxAW0Xw3kPgF0OwaiEY989LgDowyNWUxBqrYx
Nb0qpIJNkhq1HVIFN1L1mY4j8qoRvKw1FeBxEoNsYXRmppP0lBLsxdgrxPKoIBtH
0rd8MIFXven0MBRDXRxPMKeTj+bjOrrb/JToPoDKYfuskKfRIL5SHhz8Gcpt+YK7
eWy6HqXh6dLVpS8fhSPT7Yf342MvJou2jO8fzRF6bqlI624rGv7VGCOSLkaldc1E
mYBVBF3LSxQAVZdjX3VZi4SNEAQwEMYJAgUhiVqJOpur5XMsqBClUPb99Lfb2/aI
I8dm0eVnzk4r2dXgfIB2eVoZt7I9l1P9CPyfawq6CfQQWc81RANN75TyqoLNWn7n
FHLeJds6UOaGedhvq/aMkOdGetKSngPxuKSmCFu+u2zgYIAcW6Ghk4oTj68wx27E
Y6Qr8G9ZIl3J/3xfoHlS6FH8MdCcYo8rl0DpzjDvuoFStcgiePNeiS5Uxjpy/T+U
UI5DwcvQvVoiO4EMcPwYQ5msGVGLrmU6g8j/zBPaIK9I7y4JBU5u/Fwmba6Hml66
m2/tbb5qhm5gNJwtTOGrCMoE4EDHhc5z5Ud8GxvqxEIWlKqB9ONdTp3qUwC/qFwN
Z3w+ns0IWVRORDny1iurSdWhjRKoxus7K7j2mbi5nf1OaEz4NUtkX+J1M13rJawf
d5IC09/Q3BvUvXgyYrfKn7u7BK3VYu5HZds773ASS70kOvlXyMMAht8mhESsCe1U
+HSIPTDdLo3wo+C6c59uwgwiy6fQyXEwESfsrvqJm2o3Xu2ihxV8drowF+yZ/OH8
0W037SjJKJfrwivXUoWMeIvCe+5jF/jP1mY9NhrNocnzyfXbwCAtomQiecsYpS7H
AOvx+mL9UAxJtGAAJCeas6i2GFM11Wj1IIBF+NP9+g6inlghQWTJAzx6hjjXOaMO
IMv2nU//NlSXnLLXRa+HlHwbT6wFPsL+2lVjJ3x7u12biOnhv7TC5dWcCGYlkz7f
MSNYUK4mqksBaLlxeOgxZ8zuA4HZZC40UFaC37mF+q0Dr9krkq7EVBiueDLNl2u3
n1dptmn69XUq8FFLoYfCkvXmU9QKOFHV66eJEMK1h4K1QrF7fJuIT+eB0iZYElEM
N+4Lyd0CvU1vj9CXtJcHUPa1MA0UJD9EfdZpUXQmlI52rJ1uavlmwaPvPjmp2pqw
XxJMQ88qwDM3hroJg+WeViEk5BwlrErgl4ePWLFA+zKG3BSZ/Kn2Uaz6o/+0rM4q
GcRRVYTKcgXzxXNQUdjEaeQRSqmENfm+DbAX+s27wyLYH91XilgHOOco99mCX6Jj
LFhSe87K5ae9GXMclqrYCCB/AdsZ789l50oqarVMF2dLAAW0UnWt2wwxsiKYWOoI
1hw2R/McgngREPjFJBrvxMt63/SxtexL1QgylSUQzGVQAuDTiEJo51ezekQad5oH
j0KSpzU4xMJ8u8UGSKma2D4gpxoGLnb9pZ0pQcr10JreTYG6TmbVjGKDbGkuVp6M
WLO2KiaHyZSAoyocSXAGS1dT5uZ1DXyWqKNQBkdZzPSo6L3U2TPt/dr4rbOhGKeQ
fOG4e/cbI9+ryAhG8RjF0XVfcv/b5scYl4RM8klSNpx22TMorhVGYzHJMzAYRjkk
lXtmz6VpRHuzRAAbCMabu+EwqVN2nqb118esnWkqjNDynFpIOCCJtG+/hWacLBh5
WA/xRTs1QmFQ9DCEFqv3VjWjNsLjJjGnbUKiFOXPkMAKiIhZ6v5nKyxmyCE2OKGo
OEP28G4k/93y3pDov5bCaZIzgHcMfZaNSVwjgBIbv86IIKZt6RqZMcQA7wMUtWeS
dxDn6NG5WXiZQopE5QOUgbuWRqIgEDn9FfDNxaNL7eyU0QNRtRkYFEFWg38+B5iT
bWYswEm0DSHjjoIa5CjzriphN3HXXDk4fmvqyskDzXpnIN4r+3NaiR6f+sU7S4N6
cthNpt7WO0CCavM8u3CVwVSKpF3o3F0/ZHKI3gmxdpMls7/C3voH86StyKdDKlm6
BvQO3+wWShaIuJ1kCbN6jjmKW+WsoFB0Lj8VbJI7+sQMxmOws/KVtZmrhnxvBk8v
s2gKi5RfY1o8KYaw+xxMzswABkq2Vsg5tmDsNNn2hzgcXbCUFfmGeRqCH1rt3Fnt
9sPv5SEU1D09b2vfiNSPCfqR43T0Eku7fwoAuogormpQNJoKK0NLXQalgIzVkHc3
EduJYKFNSyNRPktKR0jsGtYxESXRn12ZsajG0PxFIy78HLzNnUKnTq5ISq5VfvHF
/xbF4IOusUy/smaiHhbTXczN2w5MV+AO/oYIqy2V2zG08YcC48jiakym7pgYA205
qRYPXmGze5K1wtDJ053PfF/I3OfRdQEc6BiJxhXH58bmq88KyQ/LrUJE/ssyQKsq
rxZdxKu2WHb0eMAJabRO15dRVkdgDmYBKd2d6bDGsQtZl+T2KrlFTebPTkGN5sY2
aqflyDsDpY/aPjHBfNdHSOyaxCg1cVKIcLlGI/hihB4OYxQBKaHryerBTzyNELXx
vJ9r4fPK62yPuJVW4psbia1nvOH0UlBejaOAhPWC2VQyqbO7F+su9NERMjKiOfJi
0meJsSpbR/dQolYBzpyEnmgqwJCTMZ2wX0T+21bEuacfu/sh2w8awQayW2clowQA
OdrscQLXUekmO72eOotbrwpUdP108aoW8SSFBQ8sVN+s0S4rJPhXoNWN1j91bRDe
OPGDCgi08FVjeZLrj4+4IPOiVZxZ5vzkJ89gUbwzkjtrqLK75wROJr5ryIo/X+A7
Vn7w0aSSDBIQMORtKKAQ8SiD1Xr5lLsfC1Od/DFDeJftK9U8Upb3ZXnKrbLx5yes
bQvLnBt70o2k+LsaGp9olRp/9w2dCpsDknoBMJeuEh2pliA8NypFgFv+ro1GCBTL
AxKN4s65/PAG3Vf4aqKrWMl1n8GnT+mGst6f2T2qyk4eIoUSjMQWrKVVqDAydXc2
UVEqEcPq+l01eGeJDdVLHaO3E1fyYhrhcjh338Yb7KbqpNJ46ULZCl3nJwTEiOl2
dCJoi+fbPdqpuXRNB5iS/dEzSeLNLLv/bqJF/b2wmtOs5Tg+AT249jxh9fxOd5Y3
U7DF4stBBrp4QCbuJCIYodkud7G43YO6Ff1F+4s329Knhncn51Q52n8xzWKaBPrf
eqt122IgzgN+aHT+2XkWzoQhIDkTByed5/fwLnHfhmAET9aysM1g2bK7kzde1vMN
IuDgNlQQ1LzZeo/Q4LrcqaKvtPLGuwUFr1gmt/OS2ncnYcheuPwQIzAcEqwkGd1F
sgBFeWSn8aysaCpC1SIvNCH2XygjKRlffNnfG3c3rqdyfKSS4yhBZO3/GjMumdU7
TG4dW+6vTZiky3yjBxx71FNEwcO2EQz+eFHYqw8Sd42RdWpasGDU6GPVM3CdU+mG
3fq2E+vxlUnytbCqWbRMr43ow61M3cNF1Qu3kGtSYk6CPBXNj0Sev/Fo/9tDOsux
2X8LOHjZZmEULGVC8qyEcYDYvJS5rY2oXYHU0LYJmOUogg+9C/ziRjFwjFjtyDhF
G8D4svIY4/Q+dWTVHbkNhP1Kt5sxLvmwGhL6d3rkOcYV8/AoHJX3cJxrhvCez+Ud
NdN7WlZ1rfv/b0v7YScbWkc4ETyf6lMHE/1nxKmeBStb071JJLUqNboPore3L3WG
AFf+nJSJek5tZbQn1QqhyFjrr7T+W5i9ZvJ9NbvlkNmaZuVdqBx8/U+Be+jhf2Ni
ycWuqcnlps+CB1YF8CBlC0FvRiZZkfo+fxIfoB132jek3X0YnZAaH2Cbb0DDikHf
tvVVqi2Y7XK2CUVjnq2ev6amFdvA3YPqCHzcivU7qU2LK5To7LOGteIMerLAzrJB
Jdl61I4WzIkq9I1kDNwn9B8nTgUy4G73ZjN4sNiBlEKwIxLU2YLXNVPH13G82IPk
m0J5FVmcAWRGnlTQxwxpksiytbof3vryP006J8kVWhuVCKHN9m0lGoWku2d2kL3b
GfvxZ5jd9ZHyAjC3yyCGf3tU1Pt2efSS5vnoNwaPLQeTs2TqHQWlO+30dKO0FcTY
SHc1RsNP4x1bzbkztuZ3IvFcK7cXRfU86A0EEKYujlqGBEqQNnWk5STUbhH0jazP
37ZGvw0dSLbUKUHTu/4gqyksYTlgOJYeW6zK5yq7Vp+cA86u49VAww3OLO0b3c70
/mNKK0ycQVjfRVsZm2qw3ug9BV6TMbdvKGNfL8gDyk6ZTbHEodNN/bE8J2V/pv3f
ACrBjT/yE4VWC6lNvUXWa2VrQd6+yh+RetbcseVUDVbiWpVXLXbpO+DCHTqv7rIT
FefHqysqTh+1VGBcj/tXPKC1gPtX+xuPrHaLCiNPsYYFWBx15Lwi3OjixkjjbP1l
fRiGri6nB1KWu7GeXcXLHl3U+UJSX4l5X06UH71h2jnW7lUVFPrQZ49HjnzKH3mX
9BbrStli9pVlj0KZint8xvfWeXf4U0X0E/QyeEMTAxpyCzFNfZnoG9JhNcDVy7gy
F2iCoAGfO+/SRecWekZXyGi+AOLllQkPn4NNQ9SKHd1EVtrQP1YLjxRBzii+cOCe
9TggPRzRdYa8IIQ9F68dMp9z1MPIRPKzt5Vla2fuAon01aVQziymq70ciYX4lpsE
gfU/lyNCxGk8HyCtKzdNag+OpsEjZoVJzrrRReCpp9yX5TEhrdsJ8I/RDhmO7ip3
f6I/3xhQmwslQbOfANn9Q5T/inBRR0YsGOVXDaIePdxj7xvZPS+6P4L1EJOMqR8b
B7uoOMN+H+gF/Nhyq1bH7RsFxCeVDYVEnmz3sE53wkenBQQl77N1W9xGWcwrIoK9
3iNbYaYjv9qmv1+sx9c1N2NOmJpHd071Bz5RGHRbSUqsDF4CZFldK6LIZvsYThbC
cEwsVLNlra0QGevp+pqw4Szi7cmiyujdb/osNJ0YJ6upWQf9F8m9MlFPTm21NUPw
SSGVAGMM4r9HaHb5qwiSKAnxXoo1KNKD0xVvTgbDlO3ErlX/lcoyXZH6KIj+4RmB
iv/tlWv+dVjzeD71KZlpyIk2KZ92314LVsoffy+lDgZm/lDbbm8KqDtFJCWQVrVJ
WZt8Yz7dvCCPvCP90oiYLKJpsw9WulmjKjLQsOaMle2nXtEFIFG4s4o3vlD6p2Y6
DR9LRDFnE98+cxTJKozcWs3iko9l8W8BOhoceshQlGFhVSkMKMbMKpmxbERQNWTJ
q9eTjES8eUPL/6siIgTAhpgR0jtJoAM7tRkc8QjBNMRxG/v7N6451WlhQOuK26VW
w6xaRNxSuxDSPlpFYV1s3uQuP5r0C3IAF7IZ+h45UsXOLbzu928s3idB1WtVZlNB
73ooUcWqQWHx33X9wXfWsxp8psxI6R3+j4VayN341Yas+WP2wSTjuQW6xcvY4z26
UoK6ddQNEMIBbzSHNrojF4G7rdCFN2zASeA/Kv02WdowiuyvHSLM/eUma36//3Ha
a8wwAxd7NYLBHCPpehjknvzBXqBgwzMu/TcyxFdFLysaAPHdtnN1DCtGxL5AdrNi
6XYDau7AGzvW62M5MgsasX+OStar1Mr+y9Bucjkt9URZBRegBH1HfjjUxIV6g3O8
8KYk6IFJUX0+8rcvJZqz6djvyI8PJXeTeWaHH8dis33wMO2q2/XkUmcyVYdL9BmU
XHMxmZwgrN1HVGQ4YuXU4yA/iGrB53KZeo6C1zbDlOORXC9vlKEwGINIXclpDATj
sqrZ8cxgzTJldIpf6QABaNIrTH5VCnsH1tlMXXMqblhe6xNP3wUDv6onuTZTaV58
hivQEWsHuo9fMXCYGlRFlAqwQgr3KkkRXO2EevJpcpUv9jfYH4HOeSVC/U1NlqBZ
tWxra69GOahYY48YUcpxpgeWW9ja02IBm3a2i5Ajbq/O75zPr3DG0WSqtELl/rgc
WgidHA2pEq6g1FGxzrlu/nV1KiPTX30doXFsTuANWnNSu9j69Q22uVblDioHdokE
g3ZOibIp8cK5CS+MRWVQ2rzIAJoLWH0Q3C6TDK0jSTab5X1IZI/8gguFxgJRTWcw
aCdSEmok4rrzrZQHNrMPxB2ez+gVIHsOcoKtZio2QmpXaE8iTlCKUHTgctMOINII
XjHSquNa81GQ0ZgQUdSGvY9bOo6opNe7wjE8auXrSWj4wa0ize86NEHv5/PX6Yqf
nLjvVmw78a0Z0HRfU67VlXXAnrYYntolwUa/BYIQdr5LpHJdFYOtqfOdbCDZbYYU
AB9fe4QFHi1OMo9y15ZOqmyyr7/3znM4cyukKP9tZbU3oN5U84RCWtmuL+rUGfx5
9AuzU4wnabf0cmrf3PLGGNzrP++QBpVIEFaH9Q2susrsKu4JtnU0oK4sxPqEAazA
A2ooSfNI0CcUWF0fWCJ1iCLTUlYorK5Hg8pyZZ99GgABEn0P/LVporOZL16OlT8d
ozxQppNSQ41fTRCD2Vf6G18NcMjI5Ce9qehb8B6LMN5oweBS//yad8bniYeYHt93
uvI7/UwbCCoefCseQhTb4U3tgF54YTxmAfUNy7JamPN/6mnYq+CxIiz/1mcRKOdv
BqyM89CLyk/sXxTZNKiQ9kWDWRFkmqzY++w9k52SWDvvW3SpLmU21TOHvdQLQ1vs
jpMdLK62kuUUEIGn8GpDBnpdAYtSMKzoulXnik6uUp+6Kzn49WBQTLyLSzW64xtN
c1XyKFeq57qxySOP1x9PFJsqzKhuMoeX8mCmkYYH4TAza6+8kkG4d5NxnBoloPYd
WoFkHvOij2QhwQSTsypjIonYk8rk/Wn+olLf0liyYCeAXkYPov0moHzyXyzWXJPP
WRgI7njYMOwE5hp9NEAEw2agV8pTXj/tkxVLdaDf/Xj8HIle0BHGJi1tcdVpaOuP
9dJ7Myjc1d7okdcgWnWDy+eARd4Pv5orFOkRuCEqZP3Xq0NogykEUcxsh/An/DWP
lcl+JEXIBEhyyROPKOF3XyU7PoHfj0QHiAa4HNWL/YxACiePjH/kVPb0VMnaTZ+p
oZeKrf68r8DwP2RgKserreYzCCvkdEN9Bv30UrYKLk6KWbGgGwgt1JFREfgroYxV
FsJ7AKOR2+M55MR8JmVrQYMSZZqOusvxEwk8LEyTIHnCSj8K/u1yqHqoUxCw0usE
Jkr/tWMC5bx/rkMIQEkeqeVII9uRIDgCp7cb6MYdZnnrFHlVHc3LoQX1HWmxMQnV
1MIuuq9CeyxQOY6eltIsaxWKIFX4Bv1VxSWOvY9i8w0C5NtPemZSECDHxSPkBibL
27RiPAeM/HVAaw4I4i4rQkXK/6FHC0q1YnQieAtersoY7uo4P9rBbPe8+qB/oRO5
QhiCXNJLvzC7zq8roouZn/5fW7F/q68rmnnAtf/npbSIiIQuXA08O/ZPmi924i6o
VQX7Pg1aJ7Smx8uuDLIf5ox6/DzU/Kk0TqlJfNxIVaaD8S9f1DZFe6F55mC3MpQi
hZ5CcI1rjfCdQxBnBep3ldB+XjNL1L/lA4uAjUWOgPgS71/oekcw3OXsYPJIGydM
e69z9vPj5EC7aloVb1QmahTOpnjHhBl0DjXHjRxFGiIwHSpaPZOeVGFSbJFT0qY0
oKf6Ima8PDddprc5TMR/rY4dnjy2TN6YAn114KR1O7SIIpDoWHgV8kXKteBMPoLL
hfBughMKKrFKL89q1oivddc6Lgo37f/6AKmQjeJnWqx5n73qAzHCJWBnzy/lqJs9
NKDz2LhLc/hpIZ0MgI20mUU4rRHEF8IgIO8PxxH8NwXPn04q9ewga5KISgneeSsg
Sz8+AF9D8rai1Q/CFZptd50R1cgZqo/0U5JVpJK9IKtUylo2hcFHKsvo796FDepz
hFwCAlQIweg5JXBXMq6Ag1a+p5rH26vx/pFsAqGdcj9bKRdXUGXW3e6yOxcvyY9+
X3FTp/2ZvWTmv5FDaFTzLGZvGdYUS1upT+0b7xExkbUVTTflukBUqBIVkqKYJjKO
nr051xemt25WD6F1O91vDB4lKw5JZghfJyWRoro+i2aG3wCj8R3TBqgyR/nVvAzf
/oNiU0944vwENgrzDjl16gAsRrFkA+SxItkgbkFiOBEs67sc7MNkdi36M6GNNLmi
gjGvkOaP22sx3kMZ60GGwI2AL0Usajg3H06YxuSOfBmk0BsaVGRoP1AD9YV427o8
vF71Q1+UXNMfEeb3PX1LC+Py+UnjNPPOzcI1iab8I2zaH6gzntRs6ewPps4+OaUE
eXBLD83kS9NdezedbMy5FCFVBpHJOzdhiQgSEWQm5my0Guil7jXLir2JLxFIaLAW
mArlaEMDc9X2iZJoC7W3tm5RmtdsUCQRc/oawLbN/HIhq/L3mgS6uXjaMee+R2fi
9hvYvsq6LC+GXDJbZf4fNIj9cdipXtjUGXG3oc4O2Ml93Njc39b6+7i/yMbbZV9D
xq6SUkMwiAb5k6s+IiWuHo6cFjeEEKH9R4WRGXmSvBUxvlOEiSRzttVZL7ty+Haq
AFX3U65jaVidSW6ErFMFBFUjeb2OmgXZC5bXWLvvpZ7duddFGuE/mB+wFc+wnc0K
QOmO41C3/buf08C4qFR9BjVZdi6XVO8PP2eaCLHlDJnD7eBrXwlqX0R1kj/5+DfH
0u4utHSuxD3coaRSwWuLnFWRfkJVfLcGPgaNADWuouW9K5oxrDvtaqLGij6+quEA
bN/nCpPAqcK7uZld2PA62zpsUnQo90sRwTrqQiTxbxt6cMOqycm1s5eh5350t4wl
Jv45IZ/alxco8F4jEj1MBRGzi8c0d/m/XbwdRkExiPfrg8aOyMlBVJuP9dwRNOBJ
k5BvibR+o5Wxn5IIK5KWpfzo5zbsQdbFfP96I58Rk6sbdhQGl9/UzLGauZmKR/po
ri83Y9JWqqAsvOOzwDVFgLk5M5h7p891ncEEYF7FpdsQY6XCRD2g6pYybDicbxiw
yMDkheLb3VsU01Zwt8K4onTDqc9vW1zhGxxmME81Mq0A08gjJUnBWcL8W2IGEtJi
M9sLzZDr31t7iTmrtbDCt8CNV1TTrkvFAjmddXnimRDi+9E4MQKB/yfZQlUOcrim
GpxrxXh9z6ILsR9BXGlnxs/8jLyrThiuMEmIA6RXwXwvHWH87Gy/rZRTjlstdJGd
a+C9B3owOO1U6BAi48nC4Hjpz1dqsqutFekhkuyHD9aKDGEISyBsXZDxZUYXGRre
19iRdXVIYPwYzXF3vcXrIv+0FYIxNsLs+TM1FYGRjVHvZP3Cexn/DZEOBgBucpO+
DUA1rRMEJTDqHPlsSsH7lNAK9AIN67qcTup94fzPuflcv5SBdKb6E8KbVnmWo/sK
/1QmAtFwLZKfwwujL244JvUelDXtMV+uPoy16kIOys92FgAjPj9AXcN0QY+O+7vH
KhO/irnk4zjtE8tnToRU44weu2Q2woW5iu243r4tiymV34teoh0uL90pRc7Hlz3j
JJYOCXKjy8HranuL/8IRhekoqKYdtJZS2aVgJQAPZK0G407r1ChCXpg5EW0wqQXS
CANNhTIa4UeACvFt+KF6B4WjlQK8cjpKZsxFVr9m6heMmflJRfozW46wHKDxPnXI
oAoD9EVNHnBqoITk8uQxOy1YFgATBB0CrXymatoHxkmHaWR1vzoq3eP92QAdwmWd
ggaxhgu3OiQoI25TgYlMtqBPdv74AfAets9Y0ZHm/on9BNWs8M8PM+ffa65s2oVI
wY4x1KRF22xPjKCgcXTmwjQntg8+0d6binvqlUkTsondZanbI6p6Z5fruxUK6S8a
wC0R9fnjLQoHn+krvqoNd7B0kMDksZt0YyxP1Ql1/IyeO/CgYUAGZFrelyZ3pUv+
BREyiLXPtjY5X1hjIzpksmpMncywwgtDwuEDQRK7D0lAjXBW7CxkYImSdaq/x5r7
+GnKGIPxUc/t63TLC2GLTBOvXgQBlgU0hRg44EoZEDJuiZut7U9/tVq8XUZdkWPD
axhBQPF6D+L/pn0/axGbS4nP5+7u9Xz6Ge0BJkx4Mg1xfV4WEp8E+D6aD7Em2n6T
Tu3gM47G+4ifX+x4INx+isekDzRDRyNFnqYICOzxHrnHRSCfoDUU9CIVbPhgNRo+
LfDSrwchFSHjsy3ri0SWZ3RlKo+Wu8M1AA4gmkb/Kv9g+s1cCM7j7JAAqxvIgAIH
uu2VpWP/FbiYB3LD6TlZ8hAHTy3cY5jj9Wwo0Wb7YA+k03lern5BWivdx+74Mgfi
SfJ+LzCj7PRJcFPyszAJN1x7vhadhlWJR+GET1BCptnlkfw1EonK/RAFYMtggcc9
wMBATIGdAMJUzavrvBbM79EydB6ZGPJCx/jZRdgC6MTqR4LIocgYLg72A4vGHZTn
auuauR049D4Smu58aG2ddGbC/rfxz2+gDgxqUerukj521FkdVMeP/yBfCHyYWJvO
4pJpkCyDoc5uKRKZN0JDut0+4jwfArEkewNKzhpOaywzzuD9qf8Jo8HM/v7Swocf
b75lX2uOAe7FpghHFbNatwArpsIhPsHjh8noCobuZoWk+Wt49PuvgjjUxyHrCpTR
xDDvOuA+pR9opBBhkcpkkPPPl1SbyfifrFJOyYOrXbCPWztoIVhP6Zclg2/Rea0F
0fxF3lWQW2/mMzDKUqmEQzSdF83YSqDcYBZPjZXL3Dh8k6xabw4/6pISlBihtary
cjUvcst0QYKpowW8vEOg0vOnJM3Am7GKteGymUOcy6Hrv3bnlFG799m1dgBYU/RU
Y72Mi8JcOh9gxqyn1lM/VgEsYRv6aMMoE4WV57Rai+wTs5/dsbV0mPmaRR1ZFq27
yX+bR7zP93DfQ1sdgdSnTWz/RGbmkUzJLlZ+cQCD9JkMAnLeKapz6cssAqDsNO4w
A/ts6BlFrsSZ0ac7p3k68dfTuas3hSas1jduN+NDzPjs58ern9/LkVnOKHfzCiyY
ZxQLXp4bpSda6dYoyCObia46juH6e50arj15G03XJy477qWWAMdliP1OmfxC0kT2
xcB+nxw4YJYkxY2Kb/p3vISArBiiS/mc00WXrgwq3o0+QKgnLTeb50rY57r1T6D+
ZtJSnExa4alpV35Y+EfFXP7vhLgo6vd/WHnKplxEtxSQIFOldyzTHGmdGU8h+MdG
N1XCyA/+EaSNNJlWFv6PHP4qi8l4mF3jP9F/1SrNijCqHyXdxpY/En9rKPe4oVJB
JlUOywnSD53giXgVXS7z3OdJwnSFrv9VVgb38ODWLn7GLTYFiy2WiBbx1qZWGvvH
J3ZpQygN9x/c6bkfI2ryyVSZYgVl3WB6JS4ddoYYt1n9v+41+igi4bVPCfeoQiQg
Ou4L/zSlYM5zf50vwzZtRqYO9bglO+1SlFyAiXGDdgKZX2g+Q2b8FQv2BdolXQrn
tXPeTGwYTQDTUVCt1w4Rog9nuin6U5Y+q0KOZbePEU++n3PZWS6zFlupwPRArHK5
y3iGT1a5CsEXjwbXRewVdPx+zSxkNtQddghY+rBA5tX9j9IQoC/wq5JqDbyQ3Kxx
Cty5uR2fcDVMtQDEoQagE1V3d1nx0A/4Vo7AaZivrCq/KIgAM4jeYQD1varjf4H+
mchwu8sfhZEj6mWsg/wEFBMu9H1sym8OxdtJgrXB3sPjvg3w0K3MUgSRXsJb3lcF
V8YB7YWkCVUZ27Tn3TKmwHZFR5FaTQsbFV97Ggyna/R+RZoTzcsXS3j5L7jZsq7d
nxVWuBXBH/9/WL1sEL7MMFINMKCF6Bt+grWuKU2jFMO8EDkNZiqAR1ry1UGAG+M2
hvkYMd0qvaKprg88+aZh8I+zMR357bw3KdyW33FA56ayLRpyYlkRD1iuwJ2Gx3x2
2IuXDE/EJzy0B0d4vc9GfiiRqQzeAtseSPuQQLwLCBUlrjsrtLgQpLykYnpRpeRe
bbBFw5DKtdpUOQeWABMkvYtgZI/FhEPNPeJf+dIXfoSD1KG3piSKBlTPslPXZPbt
TK9os4LM/nOC0lasQD93OIunxBNoOgwDvhYyGJ2tLh6f28UzFR3xkzgJ3tRGNppy
UJ1itEkA2AL57R6rKaE+6unQ8TEsKGVHe+wxPjAACPxeurajZ7sLfvZiVN5kt3fN
OeIVoaLT433EAIQGZPZubgGGq4Bzg9VWR8+M0PsqZ62gbKo1kZLji/MH7ZX4zu0l
Afy1DL7uCPeoqZWi5KZZNz5rLM0253EEW+4XppFs0GM/P3HWhA5nFEL4swUmP+jc
g/3uSAZcmRks9ATAr9fZ9Z31261/jghtk4K6ZfGFxXzUs7nLocK7uZFE7mf1imXg
hdv1aO+AtRfX5hG1KSvTDJOls51LNZ/tnJNWrZiUc20QtR9qq0fmkX1Z7S0TlE6s
gUgeCOKuUeHvSIIsJexygilYGuRLJUAsZfoSe/8/VP0LLjXh6CtGMlUVJFJZ465f
FGvRZDWRd5Yp23zBeM0faAZTz6paRUjNccK1jSgsP3AG4KCzJUV+R77t/fLES4s8
UstlXvwHDNEjHSuTuLllGW9B/x94qq9tTN5uE41j3SRMvy4Bn8sBdLTSsM6ppfcA
36eUcyhhF8zIdCISI6qk76FvSF/2UHRsSb6L75eMxWEvWU+KkQ4QvRulHQDwEu82
8bwR9KCzt0GrG4Cq0nBKNZDzOQN9nJ2o7I8SlLi2IcssKRtd8Oq0hosEwjxiPeMh
QGqNHrNzbAUbKllzBBycqABchzeBntZsmfepIsUR/eCbj3KpcW8Mj7+pZ0fO3UUW
kxkQ2Uao7dH6+OykqVHIcvynvHmK7FmjX6QuWNVXTjlWuUMa1kEI6W/MamWLSD57
8oYv999kBQnhTzUdgbW5D0d7wctnQIQrBRC5f/Vb6EBBY843D59Cgne8oCOMEjS+
gEIN+T0cadfQDt0nYZx75lRrKLGyFvKGAnhGi75YWmc5OMRzFW0z+PLu/cYIkGQr
ZIRHcJy35mkNXTi47l48cYGMzTt1AhqXdguY2Ku9bwAhckcqIZp/bCMLq0nNkVya
Zxe+/AXQLyAerzKfmaULJ5rXf3juedI3hnc+CzRInw5ZIN/e5yI22D8Dt6LLA3vm
nMkj415iz/gjXWmiZtOygGtqDP8CDceRbw4EKozbkHMIZjKigw/xdTQ3E9KDXpQR
rCRx4wg3eNLDRPxLdVha6bo3uhEKlIrd17jzlYw6gge3/11IyZ48FM18clzIo3+a
RAqNf8AKA5F+lsjJTAxt4KBd1Piv6Ncrfq1iXGtYsw1vl4hpMOR/AQyAjakPVeO+
K8B7EYLURHo28/uioCOyPQHMtFD5E49EJ0pLIG6iAf3u/E2LsPCY1RMkNIXyzwyc
rtCPEdUetFPOB+haFmQ2QXOEmtVXJGlJhw28K+78sjLBlJJ2Vab/tX1yUfTLhzTL
WVdhvlWSU8gbTuCxAx+Ds3o46gGrKDKVXiwH9Amw6GnuNfZuwjnt2yfCgEiK2tiF
0KR/Dk5zBo65J7IqgRuI4dZ2y390ppMnqjQhmVf6tGDOVR1QkW6XSx7bsOrMAjrV
i553QxFwa8TfD/mS2Di7DJ5Kl0/BFzj7Lhjk6r4oEfahNePGJofeVgPWp6msTS8E
v8S/cj9BQhyIDl42WPg5a+AGHT7HdBJmgP0SiOU0FQCjux3/IXFfHRIyzYEOfy+t
6wn7YRbzSpeykXMsgSS4cCjpdTswX4sCb1mMXTduKji8XkIlh72lLCmczZfVsk5r
dQUM04oIirFU96MQVmnfTPg9l0BlxuHs/FcBbh6HN3+nQM5G4/YCYm58DY1b1+WO
TkLCXTGkhK/DJ98eoCJrw+B/eRSzFpVOsYbFG8/f1dn9c5WG3s0VXgMEaKCDfAJy
7Me4op41dstwD3UbK3iSaO6jAUMGSu7JWDUGvqAtNl9E/stOPfk/2VGAbeLqo74M
XTY4A/7AxVPQ7FRusoF48zoUsv1u+7fn5KIlHMkyc2WM22qY6BmMTn2YH/MiGY4M
Cy7bJV/vk2lGcRbpOIA4gpvn7nmghkNBVTokxOpTxlCJvx3sBD/I05koEQz7x4M8
BT8K2MT8cLyaSDr2uYC+nlMD3s0aXuMqbzGBPD+KV0WBGB0q4+NW6bIGCzpW14R5
YcC9bc6kTCWSIc9C7T1CkHgNLP8t+o0AYvGLjXXAjHPka1HNocuQVqkQsIkeCmQ6
t829dRzyBBb1+RPHSmUcXd4DI0UrqwAgkTZcn/AkH82OZRnqseOBgjVcbFAczbNV
nw7+Q6NRU0xzoMmc/ELzjF79R/ZwgUBnG40sFeXCOwqxEzbpQQpJS0KSJw2/LQEr
3Bnfr/i+qrncjcJa0wE/kDHjfa12Mnv5EBuX8ykfgLqrFdg+J2qn78tnMMlWSb2p
EQpE9JmBC5YAw2CLy0adgl6CK502lqLEuXNZ4I99cTCRVzBnfwkETAAns8xk6HdF
3EohHbxdUcS96g29FIDtcrLK7CElrCyCtV2hlZOomoOsxLU3xwXtqc+F1m1gNM7J
LRf4z2QjJGtrIeEWKsEf2pE6Q/JHXTscjShaZfeRqslIet80JiPQKhb/2u4ZjqmA
MuclK6LBYOyWKRR+8hourjzas69WpUwYUcw+KQUiaYClDCLlA9Dk0JuTrc0Pxkmi
+tlc4Iq7Sf3FT3YGwULIGRvqC1+JTzpBy0fy8NSzu6ooqF/RTynfgo1+xXKMiF5V
Rf0iNDWKk7+wU2P7v18Kd4AkC2hBd7lQjfsrJDj73DPewdTMQOBNzsXV6NAWXqxk
sPKQUfxqd2BVcP+0IEMYLNcy+16yIkiHv1ijM8rMS2N1BZkecFQIqWRqYxMv4kbE
lZIw8UMIVxqrC8HQBoB56q9rfvDfV+nB35wT4/BPA+rCACaW/iDMk7brN1fG89Uq
LTezAgOd6YjyMkmSgNGnoJyM24kz60oOQIez0BvGyxXeNypqQUIj1WhBwS+RkGAZ
7kSTaEUEGndsGSfU+z1SifuX0I3UEFabtLjz7gE3TkdRPHz/z4T9Fhw//Pk//RF8
efD+CNZ26t3QD7deJkElbmY4UBnaeIai5jHGuuNE2AFAEDrAPWet76maAxjC2dHG
yHVqkfxZVfT2yefM1i1chTWzKfYaB6363OeZetYnEBqnmhwKZVCwoG6nwUsnEK/a
rwppccenKH+wLa+o+n0UUnzuLph4nq2xxGdwqNhNCiW5ez/dKMZl5VylA0iPTtXA
J0xVVGqcSJ1o3KXzQbDAzVW0y/TWeZEKXxlgzx7SA+dkVBn4QDe8zjlSAZSqocEE
RtN655z9i6J4eGNKcmCHfoxk4xO0uomtbtdxBTn4MB+f4MPbDPn35OsJiCU7LcV2
UksHq0KAHOybJRZ8v6Qd6dUtIMywrU7+LGi1bF4rK/zM3mr+nFQbRVfTPosbhZIw
A0aL2dCKGWxaZrIgvPSlTUnCz5V7iVN+6cbs1jNfsZXlwISKggxOmJ8jC5T4c4aY
sWz/Ok/4au1cv0uPPAPn9yxbkKZSeNw6Cvo8B8EzP9BJcThpG1eT9LwQP/8TxXmv
Y+EnSXs795Gqalw+FpkrHMaFUoTYUmNX9lotfvSPhkuTiFLd4TS9ZMNjm0bqO/xj
zfu8Uomblq0MvjzflFSy4/E/i6LZnNF6zUlLoo/xYOqx+d/+B8/+GWFzO5+7kUtv
6wOoOxF4s+5Bv1lRn/+Qucr7isSiAYSznqUGSaP66C5YNHSlUShzqpJ1Hbdpb6va
1L2pYlL+MJ6VQ1hoCUb8R8XbrX/ZB2eeo740VusyyfeYgV/bhJfmp3VHizzgUKD3
zfRlRyhq1Jt+o8vR0HGAW9zbOUbTmBPTjJlzXETXpBHzVyPhxY41SmB/Z9RLLsgb
wIRWHkTIk8jA8LlFNTZRGCymVm/gwdwGNnYaBfnBrIYcBrKld2WMRApDdkkZJtFj
EXBmBqE6qrZEXIxXXEeL+N+EtQ31ygCADyDbzNM77L5CbukdOfLOnpkMTz7FVrNu
T1FtkviPTQl2bX8mDQkGc77IB1Hjn1wsGSXwr/dMe87eEB4wyJjV0H9aztnvdQ0w
PEPCR5qNbHlgyPJvP5fWVrssYLfj4K2LAYPXukF1FRFUL2cMSNHlAJN4yh7Jzm2r
WbwRDvRG7MwBRQ0qpEGFDEZGhbYMWRweRik0r6WgdKsreC53hC+DG3UxpKRchkd3
+EDBdbSZq9m+vuXPfuGribZ6ZDH7pvKZapDHKYOPsk4G2u6rlCbQ0DW+4fEzc+lk
JZrvcql9PGTxT6Tc3Ho9y1QzXk2UKqIO7d0Uf3mjDeggw5plXsfm8UQMBmx+KJtK
jCC2RVEKul+C1OuiC4QWVs6Jg/cnEsSy/0+g8LK+CQFlOHITELVJbdn0lrEyAIK+
QQDlaWkcM8057KJd/D0GCZnGv1DbwONZfhfB1pbCX8dffyVE/6PoCpvcWpMH20eL
j8HP4yPaHTA6DSOhIbYjDgX3tjv5M0GM/gXssWqaWQZxgh6bvnSoPhzKxQqL67/o
isYhJcNzo6G4Px7Z5wqDX6X1sK44uFu/z9JFS+xXdAzRbnr24OaOBpgk+3L0KPO8
BDFr8Frsy7y4lXRFF/jfLUTQwN0wl7YZuJiNqFam+4Vjbj13veR/EQdmNOpTtVxe
+bKrrxl4XkCFU9aoc6YpehXv+S9wTEnerp5QGY+5c2BFk/EWVfO/TGaYg9KYXn0F
vhViZRdD1jc9dk46rlV7xXlm9cfmoUpo6j5d4MeDpirJBjHDD8RRnoEfRMKAAsE1
tIT0ZWusoZ14yoIlKGQ8PIgzKEzHKEGEIO1ulMgdhnD9ezOTUglT6m/OOOzjv0I3
lvqnXxWEuO/DGe2qS8l2BKAUSWwprvGLMNE7ZXiDhpXyBbj5r6+Do684PmoIZIf3
VUhr0Pvk/nBsjZ4xO7TAndoNHWkibQPzB4yaVN0PyaAUAU9dWOZJ0GzA+fFhn411
G/rPTokNCAZTlSVoM842YGLw4kb24L1tPLKFGo/jp0hffg8lqIoBPZvZxJ9l76ym
MEtcMHyquGkhggZmJNVTUSkrybHonFefPY0wEd0ivmHDia5Dc4FBXAinygbPR3yk
mVAoTktNlM20kucM4uPiD+UloZc3CmYc1J7qhpgXPjZ6qLIgSvtdUZvg2sFueiQK
crMX5K/FnjwLkr+ilul5jH85ebKL+nOWxVQkp3hfz/SbGX6uW2KdRpr/ngsHNPuX
ZSkRlk3T30mCKZvaSaob9KRX4uZ7sLA6+3d4zO+RiClKW5H5KoFNWbowlFWl6nED
n6mldnZt8KSwfj3WTAgrh3ccsY08w7KbViZnb8DwLto9Llki/jvMJ0V4CSsqRdR9
/miP4eXEH6zTsw9JbOp5uX0LmjHM6FYxhyQhf+qnQ2ZZZLjX15S7qu9VMGBOFasn
veYajElkU9Z8D2+VCwsxYujsNeHXxt2tjxu1KOwDb1iPXd1pEwYi/2w9UgOIrBkf
Fk0MivskP/YIGONdAbYZ/zdttPqdDodx7FZByldQiVmeThVD6wPLBkljSjEpvbfL
JQ9JJUkF0NST3BbXCJc5UcBFMIOFI3T8QCiFWIMI+WjZD/hmm9X/RFXd4MQGP7Xc
dQfqI60f8R6iEiaY4ZccTf4C7VpLpgD4F6YR2QIK1S6YHlkpZcUmRdQcFQwo1hLN
F6FmZYNoWZ+yH/RQlTYVj7tM74iiBuOqMNr7tmUGUuvVyMs83yoE7tW71dKxn6A6
1+kAnNpFBsyOspK0EynkR18/OOGwEi1cOLOGubUP/FnCB7yOwd1TSa9CJyMRkJC2
0uoD8PLHFgsRlBAd4WIK9BoMeZKsYg2dccEA/OKWQQ2YLL2HpgsKlsCxV+q2v3p1
AHXfUaLH0nmTbiVG2GQCIt5tqkK8n3ePsNLdZmxaw7Lc/tBePaYNl1rgMM/7quyI
hH+A/TMQ0csS5efgPmR1TncKHzOKWFDRceKFpLxAwBG4jO+rdCyaOpp5i41KUr39
GO8fiqG4YXYHZpwRgjzcHkRmpJR2Dhiip0neBKCAUAZi8cZGFv/xCe6yqwZBozyz
NO297GV8SOkum5odC+BQq04VebM6Ji7y9Caq11t5sbY5Ayz8G+TBlQB4XznZm29p
5piO9KWymk4NAj5+dGi2ogTzfICV38+VMp/Cv1RlfyCEDpAanXyR2qImxd26HI0O
EAJW2lDyetdo1qrUA4DQrbaTyap2qb/5dYikVk/gcwnJ7sdRSVvlu50+5Ztg+JwO
nRagBfldpzUpVCOoJQsm7sn4DdEypikvrtENKYiSFuUo+Ir1kOB9kZqrzIyXnP1n
rUDfq91iEc0InZk7T9NrJWjXuXa/Bkh04GxmckeeDjm2qdmbXC0gzq9naCfe6mgt
XCT2YYl7qMhrE0Rvg9W4m9VK0x9pGYdIlxIwC4sc3+Qot7WL7ZiuaVB9EtAtW6Cx
2ek0r+pZw/4XHVN1ae8TQ92BBCab4p3fQPYSfKbv/r62pbooSnKHdWdh6HzkwZhK
eCdkiEYj0GSxb7A2Yr3ZxErLJdTxQ+je6fune5jy1C0gm0aTWy9y4k0d1KTaohv6
KseWlroOI28O1JeyY+RBl8cT6WfhsnIVNYLArqQCFzkq8vZ2Qb5POACazNFM3eyO
jGcI6/Cvb4lZsB2ZK9yOMJsd1wocWs70LsjnmroJfmfCSZwuNhKNeKQqdnW0oIwE
RAJPSeNN3uPIQ9v4OKd47Jg/IhL5z2Dpk6PO3B6/0ooF+D7hnyrKXXu3x/wpo2Cw
vXtSbf5nlunDtnKh2QnSo/Nix0yCu2dWBMcqTB+j8IMsU9ChdMAjxXEo4QTLwNcF
OTu+kisVyNfuQB08dyJwP/6ER/gVVSTuyb7YItNX2scTvk8eVBJUEfQhw6sWUM4l
eW23ddQnp/+UISIhMznvB5eDaehCWYudl8Kl/DCGGR1UQx772yRhlT81iZJlIkbf
vijNnTgptOpEbmwMZ06NBhGB+e7FGnrXnwdwevSdqHMJM5jrcwuXRI1JLGabYFvl
NmHr5su85ZhtVFIZ38S0ca6+kycjIlFQaMzWOAJrncIdMzRseN0iUNwJIBkEexsV
e3mJULRXEP/+LlrRYcRYbvnaqDdkeqTi22/fqw7OXQekrceXXCkHlRk7/Yf8JpKi
436FCggcer+xJ9n7KqaQovC2O4EIhueqThU/biQ4mFNH2BzxOnBXa4jMlXYgoRwt
dRPd0P0qhcv42SEZwbQorvKkAfkpERpiW/38dmwZsClLvvVn9u1vqwYWpFnQm5FC
eWb7DV+/V8O0ybJH1H8quPT4RPzaQL4jDmqo2Wtd/0F415Ii8IYEYHGemUhL3x1l
S2HZ9BukT4ncG2hDBZxTyM/6ruFIyzQjFD7zFVO5Xjc+vhKecKCsbgcqXS0Q2FAk
WTof9UvdlJJUO5/Yz6mKi9Sapaty9w6L/E0ISIRzSleEZl5xDsaZ4RQn9mtV+2wG
yNujlGXtF/SOIRudtpmvpFrZTMVYR5WwDocWncUtudGeCgZ/htqFHQpX/i/ua0MU
qRwRNxu6oca2ys3DH4KjVrF1Zdzmq+ulLKyY5lRFd5ZIWvXEhZ+ewAul0kmnqFPw
CPMUDnZGkotmGtgqtrXjkFI70K1FQmjvkG+JuMk4VPrv9H7fqgBi0+cXbFILyGds
bGO7Hlj+O1U1ZN2PZBxlyslmKgpZ+IR22RP3/EOK4BXCoXM6t43ORWFsscrFiFqS
s8Oz6NDTWb5TElRiLRXJlpbbLTAvoY0oyhmtF8Xne9NNE2R6oJ9XYFNGO9IPjrji
atyKOcMqWwAzgC0DOuwTL3X227IMnQWrMVtZWzSG+V4FwMcmSUSZo2YEe7j7HGc9
kCWbEYwOTDnJvfbOV3EZm+KGLxKvIB/ghKynPSvC2tC4ZAo+Qo4BgH+yeEzg80X9
8bekGmz3royGbQzmS/TtUjXh8UaIyb6tPKIcL91hNl0kb8GTzZqYHmg21/j/qB3f
3CcQOiDbswpH1loARjt3D+XZxhmob1FcbLfonZM1HJxmtSQyVe+w7eH6dodwXvy3
81E65DxJEH7NOAqptYDwHJzoBL0FtBqjW8Lvp/pyk3tg+tPi74o3l0Yb2JI5r+IE
/FxxTHD7SM2dBrwDQkgAfMEJPmNEHxckmrJ8T3w43OJSYJie+bZ+k/4KYMXpQZ+u
MKL4KqoSFfOcLFck4tDFKcDBpF5cldol9WhQ1DGVXhhRkLMPcLrRGdTLLpcqOUfn
iYfl569EYZ2fqy7x7y8aw7m7LkdpD9gB6dvhaopU2EPmWs754mbaNq6kgcYTiwnr
arQL6ZoHM4GhihHQD0cKMhGByJYMdimzj5VI2FT28Z2XBET+H4ry+kWV2iEs2jFt
lnCCMrcKyPU3RFVUfKP9UUqzjlOeRoGqD9PTbp0Yx9GKIvbHYnXG3vOcN8Iod6Wz
0biNxcgCD/ZS91+bYSPMyTiTHC6WvJXXyvkqKmYij30lzOX2G643ZsMmJONB7Iop
E9KZjnSM7v+aENhT+rXiEKqMpyAazoe0OEKXBM+4jHkkkDJyYXgPEXLj+y/QMNtf
VSWaYhXglosrzWB2/OXaOpicLmAMeHqKpLofQVuE7jYMvv33l6PfrYEdXf/r9FQZ
jkK9/cWnAnMAg5RjhwCD454Bh4Zzx8pMea4Cv7bxqq+A61kmNRFq0Y42bVoifJZH
4TIeGVmOuvN7YVfeu79UL5yt6h4HAKyOcxo5YOgiuje5EJvhkpAYpANAmdxGMZjp
ZFow79GiyAt6c0dt82VPDbnN6CTtiHH2/3A5XWeifiq7HlDxM8tTmeTeePDP8e1T
uK9QJMwyU4WPPb+qB1oS3XyyBxZnyOzh6F3G6m8u/QeKuJWDjDkG+9Yf9cjqTKLa
LLhDzMffYTWEc03fxuBtQjzuKzyhhmywbaj67q0x4+yCRZ04rQSvoQCxHGNW+a6e
OwkinlJ4p7zbfBpgEZGSbWIbX7RhJWleGIOzPIyljcLoCFn7pJAA1gIFbDHl6Z4X
Jivg74obiJuUq1MywrQEqxs9MhiZqn2rHnycWmcAyuUJdeT36XVoF7hyZ9jtaE85
vkAaYzRX20JU/jdvjjjHovY8SBYnv0uGBPW2G+zKL4XEj8FJWTmfO5JS1TPItNze
+25NKx55cS+A9EO1YzZS/u/KPzn9eVwwpysfB8+sVa2IjghCmBBbjpoi7Wd8EcY+
JFkcCx7SmqXtr17Gq+G/LfzZsRk4BP/GFwEhHTarxZ+8hO4u77I5aLYLBDB7x4np
DaobjrTd8sU5GJU6dDwan5o7GZ9xnW2ZExU/NqY9sxcrzKgBlDE1Pj/nPA3sniyI
mme46eZHNWz6M1SLUqv+IJlGTiKBZt+Pey43FBJU/2wnZQAuOX0mP7jgByl87OpI
MQKcCiyhJ5T+MS3WykwOEX7ZxOGR64m7F+TDg7mY+L/LY2h6hF327BIIjrLEr28F
fSagdOQuSbRNt+IV5QrZGKxBIIysI6I8Bc3YUPawdXPJJUtSHQQsIX4dHHMTcRl5
FRdGi8+K4bSlhdHMofeeCJB8lFzB/0QFgOiMPy/iK6LU8Bvvcq1GrdL3Y+SNHR6K
pEVzCagIG8xhM6EPE51gJh16AIFWVNotSk9V+MYZrJlrbzVuEME5J6IwIZ+ZrRxq
HfMEv83YdZw/k7Zbf5EmnlpmKy+nzVgM17SgGHFoxy3mDf7THBY86VDnnaO9xiCA
z8MxzzScPY5Uv5QTOZ18l/Z/OPpduiEIYYJAv/ze7IJASBJX3LDZ9EreRU5JiF1V
fHoATSn78gE2ZvX4Ze6HmHcfdl696nB+GjOSaS27yaAhra4hT1d32iSlw1C5fRyD
io251HP46eqVmDgiZQ0Q7fn7EztHI1XfrsVuOFSHV6V/PP/M24jAD8Yk/YeF+02f
HZoCXitV5mZX0gnKCMTdQ+KW5AYHf1KjylWWRxE5NIZ0PV/IKcRarhu3LFE/K749
PXWO8La3sQtE92eTL1pN19HMjLM/qDeRErbJ3afgn3Nu/aM4e/t3+SJ69N8kLEDY
d/+i5tXbRKfdwT40wgc70/0QUagE/snYbf2Uw4UcJ/Hq9zVupcuLlG4Sp4+71Cgo
sndlE/lYF5uFFFWx4La4LaVbHhIA6KBWL53rKn8z11eAOstwWp5wp/EXoOG9ygEf
OnJoCHtGu9xpgsobNHJFZ/co2PS64oUwQgAQtM9HwB/LbCqYfXtjil3OtvwFwU+n
oz1bDzhUnKis5bDE750ybPi9CLMTw4B4wiE1WFYzlsehcHCEW+Wf4Sjx37/lhIGQ
6JdrCwEZhY1OMKP9DRCMLY+jkYSA90S9WBaaRsm2B4baBGi8HzlNsCW19xtVznvb
MA49c6MChcrN6iSegR9/Je5SuMWuBHnWpOCcPhCWOorEyGSLfoJDlpD01gcOgtXH
uVymtLa1NRDx2gogW+2Pmz3iJw5K7dRYQbYYLWC9Trtomfh8lK0NeBxURo65Gg/w
/aHhT9GXEzz7dPCk4DTN8KYwGcsxHCObboR1+W1a+diL8FtXL58dlgto5Np3YXyi
PPB5fJRe6K2d5VnPXXAGAU6L5qTp9v72eUmwZyIzUfTjkL+OoUq/HdsUOuETVTMO
7kB3cdgotp6EMh9o9DZG6xSWyFa87qCCUVwOQ+h51+aeFZFwXFvdDpxMztB8b9BN
H1S8Whby2nuuBJnFCv9HlKJjz9unhWemd+uaWEQq47GcidvHTZXLOI40n+wnmTqn
7vXlO2WsrlHyklkHSZgI9H3HOziCkZtLuusCsuCgQb1cxdqeTayDCX5j1C0eUFfz
3EcunBOAUje234yz8mZ8iykM4I/TOdbJU+RTT98f9uiCmjHDG7ft+m1VQ8x0ArXh
wPI/JPqACexWJe2iL9uQFE85ZfDnWElmOfSr6o5K/TJVKm5JfU7UpMuHfXQBmYNm
dB8bvvSPndFmPEDXeDjP1BV37pSpf6e/Bv4Z6oacxvgUWpOVX+wA+EZzceDMrXPh
EfteZliGL+lXDEBPoZVZPpFiCXXEKelaCafEeRn/BIlr3se1RB2QZ5LZVrx2aWaj
WQHmCFQfB15dFuF5C2QLmP3yqwVLe4pGVtkhT92cr5MAKxr/L/OB+lH3VRpha73R
YCoh3phGt4JK7IAdNlQVAgGxj09xJ7QvfgMP106ET1EcPMcArH+f6LMbPd6LZQzy
PRKxu6OSXuyhWKVD1RBREBgdrZklWh66+4ofxxKiwYvAWetzCn7OH0L2Q0Pw5cQU
W5pO2J1R2nZrs0wUdgQ3UU8/iT15gJfbFScTPZApfbFy6nfqIlLGSU4QzGXOfLDX
ciRT4RrdAApsX1nT4c3xXK7WXnrhmZVgavQc4hp3meUT9rCK2U4IwhbK8Kv+VIWE
Vccgm2HJKK0CQOTRUEoiriXQWz2jgnhCfj6IDrEGA2p67GqzWWaZbMlpmvqdZSLq
pPfTHMqclJBm7DqCv28iPRVIIZv8GlNICRqB4Proj9/ri9EmBhyXTbWjQLpYDDeC
7nVOhQu7OZiip1nHCPm2e3Jg/GnrwEi+NXtMBYabrjKENK9MUywUW3JzoFNSZDRb
XbuEDmzR95IBqT5uE2StIGmd5YkISCnyzsKM1R17UFyqtHI1kw/D16iqy/LMeo3W
Ijq5TtaQPPf2Vuxk5SbgP7yl/M13Ux5kUGvqyETGcAKFUIEDrySTD1FcH296IQbi
NoIyil0PLxrtnltRPHpQZjIDPHxlLLiXAMOKKl2T/Cvmz0oQpUXCnVrG5Yc0mxKe
QQ42lkyspgeHeCeyXUZ2IJFAobXesgx+8wYLDxVW8q9KV8cPCD5w9ir573U/XKfs
A+OW3DRJConf8RBlc0ZB6YE0alkxukfolju13a2wHG8MarIxcb0z60Hcqe1wAx90
ZikokIZ6EWZ8h7ORVjq9dbVp3B+b7yX7VVEpslNstSFl8kyRxkdgEn9ZBahwgcvZ
T7lF8hnU66OmbkNZSER3wO9e/qln5l5/GUs75HGt6pmn9GdAhdRThi1TLfTUmf5b
PErks4B+CfmTeL5ZP2vt4xmKfySkKDRd+Hv1qzJh9Q+MMkyCLT3yQfrF5JkEAc/p
/tXPcTfdT6rjLHnKNsD4+jZRW/zTjLCrWevqCKO+nPPOpM97z71j1xJZvro796Ze
tZRL5AJWQTKnb6UOOrxw3f5Pig2erscLaqVfy1NBgY8f+TkTsp27i6wZ2ZhpnZlq
CUedZ/fNRvVocAPIeoAApQV6VcwtGn1gq4SWd1VS+MyjfyxaUSzIpFmkMgO9rnPM
MhH26r1FAb3C024bAp3nP3KXVGTEajLXa8Ijyn2mStw0DeYntCzTIIRaRyDjLciF
SeO54EWhS9fWc6tHbrttUeWokn0A1C0y/0dBPhakUCPghgwY89OEBP/m5ZxIIkt/
Xc4bcAkdT6HoRoiNMBRjD0Ru3MSIfIksYLSZvBqWAYpQNdYrCz4buBz3kTVQkGF+
DLduBhM7AojMhNUgJbMxYJDlgaafc98HhVBOqmZV0oLf09ikwtL8wffSsqLSvtTc
mc1tQC02ZEWIK83DG+NppTHIcA2EA01Res1bdzmuFnzf8sSzTVhXk2h6bvLZyHVO
vo1GCMK0MXo4fJ8b3h1EbufcPPMosd4EdYaEwecgqFO30M0ZrltGasKgwS/9VqV+
q7uD7Qf4c/sL3Jf0meWg/5HKNIeMr1VWIJ3/8UekqDl0O5NV5wjJmSHIcZnQsNva
4dy0kZZ2/aj9r43Mwwit4DWuFd2xLNgFsj6cB8G2PR0yS3Ln7kGj0vy3RYT6K0dl
zCTtioU5/z/2Xh8okJcri7mzNCsWW5n9/aVZjCah3HHqIh7R3akC0QsG1GLlSXob
VAns4z+dSiwuyiR2AIBdnLas4pbAGlbCyBaMxyiKcqDh6jynfLx1hqHSxaKKIJHn
zlnZ+MIO3inCQ+TwiO6bSiqr6z3bpMpxou6m7awyZM5sF2Ed42UePQXaVOetpMkB
b5gsn/9WkO991eiw1kOuewTWNEMgcuNRn58eOMC4rxDn0ZzBTamNQnDjZpznfZ58
TmEH8tzxRfvpnHovK/k1ahix4xRW9WB1oDmvQ4WqYN1A2MB/BaNyhF9xp1NlB3ab
BMVT+SKzO694Ms3YB+Ily/LWPGKatrEyjicJmb3OPh0qZCQkLm1+uOabIdmWR/a3
lHFprTTNej1IT1UY4eFYUp9rM1B8LvkU1+FZg52c64e9n5XLC2yOLAPkec62FFXf
nVs1hjMhg03YvHtKB9UqbAjnoexqO5QIDzJKB7YlFZLVljgjGsuROq0dOvUQkG6L
s+NqF6xYlUpskkNrFr047hFZ4xQ7o7Tj2L0AE6l6Jhc42NkKazmC0iyCvMbkx8hF
zXykKrzkPZl3iII26/85HgWG8cpw7elHc7EpRy1fst93efGwvNzZfuAeceZSIsax
IVyVRPPWr2KI59ukaknUGDK3KRvgtX2Hj8BS6UZCkJ1ptzov3ZJJ0XdnISUkC/tl
0qMHX8gdEmxB0WbsOA1yhuktyYwotC2fzVyv+nADV1lXXaBGcJedZeaFJwFBTtbs
bhky+23VAGNlF+SCCcYy5zjfX3HZv5hnMgxE/m7SEG06WIp7wBp+ObdXYQ4QEt9h
RsKjMrsE5TH5QTRSaLF0dkIrnRSSZFM8fwdUExO+Zmyf+Ze0OxKraIvt1n4wTgL0
2GGxqLXrOKJuwrRytAIN7wpqnJqEM4crkzQdsPKqI6yO8mvcPTmg2aO+8o9e3Kx5
JJxOlNOrU/30ImCza7nvtyCOHoeP4x5wvi78ojO1blQRNDLlj9Gere6ILIOeT0+D
lnUeV++FoX64TTtu//mTXFhZy3nQL97zC4S/cw4ncdS3SW+XMXG6LFd8/IWFWrWP
roiUGXHPOlU82jzEhXaRB6DCsgpuKHtHKB5571fTXxnXLpflW34IpRmLYbBChHgP
sfpFeBYR1XgxcDgdYrfyvUwI9Zd/f0ZU2VXpIYCs3fcY+6WWmZGGzR7M0Bb6dt7h
64AEXDWBLgFg8A/aRr/oRUa35y6tql2jv+KEB54l2QP68BeqisjK0BDlubaJXX2+
RixcyCQ2rN5QxjpquqcBwEoEXOyHLVeXtCQnM5ygsoe4K386Lq2GrKADC0Fslvlq
/DiCqvim5JgEVIF0FXTzSzBbmyC+vfTki966EywkDM9o1nSQpHNQoDsqV+fvPwmc
tO97j7cFUvU+y22cSbjDxfLlr6x1mvDf9gmLdARZ4uItdgKrtSVDUcl7wnOsRiEv
zUjoOOT9emCxolH7iFLe4B87SJ7FprOGr2ajzUAiQbSGnC/8vEyfOExX8ra+NJF+
9K9YSisvn/xxWCna5G/o9dhoNOAhK9aVPZPKsN8RbvdKIroKenAryVuVS208A4PA
u8097tMWCtKaY+llI+JUJSqy3QX3Wu8VX0PoXhdONdQU82PerhjqVkoModyvkCIO
/gx4KOvspqgN19qxy7R0WLrOWWdVKNQ5pQYH/abphLf3GfDmyqhEgqpKVuJFsz3k
9/GmKc23AKH/RVGEPKh4VkP1H8K8PkhYnOR/px6e4ExsmXH06JBeZycpUMk8XgNE
xbENLSmE+zmdGdra+Ud8cePmOYaGGru6MxLnn3pRVUQzqUk5/B3EjPywiEzEe73B
iBx+dFvQsAsVUueJG8SZ5N5JRrrR8erSwj+JzIh0vu6+Kp+c41QMgwt3HYS/9fkA
WOz3ecr4AcoZM4z9rWi5p8x0GYLsFX9geoGTXH/UCLYemrxK7Ck8fGEYii2cvzg1
fFqhHQqgKSUkjEBlYe+AHfup1MzKFPES3oW9FEhoaw/TCyurBI1zOZDH8Tqnhlon
SouefKbPqLLhBZV/ja6kjlb4c+SLZRZk5SpXvu1kh+k4RJbkmfb3Dk2fMufWO2V6
zKAhLkzxTATDnUOroqksoBMZUCs8AhlE/QhBBQyQ5F0HCjB3F4rv1srtysY4lpoX
gwFBtI3Z9+kI5KJTLRlyaAYtY05I3QAn1EbEJQKOJVCBT9luSPHtJcNdgk56Ez5/
SqTntBLrDlFqMwBZ7/of3X1oxHC7aoxpzXqe+zc2/3Se/2R36m1lLCYcirT8eWuS
/qIO26YgyxOBz5ESVdqXTrneJTF/gP6iCwQojoa76Eu6fQlcIBvlxSXn6/FgcoPQ
LjTBZhME7IWyts5C8P0yjtxWhP499PKiZ0vyveBCNxgl5/XJz4FW/QzFQ9zkRDAC
B7ZBlkiuuBQAE5Yveh6i6pLZJYQf1pEjjxQWXe7FEexWeJ2mV36Ac9Iqt0sxdR6S
kja4CvYTUaLpvo72vDpSJ3NkItw4B3WMPqmx3ekbibFbm083ApLkQ8HHHYeyPkCy
BXM/8uixs5QVQ6jNI1Y3MbAHg8HVD3VGR3T3nNQCFHsLAMOdihzT0rYczcIxeX07
cNp5ZDxbpdPUdIJdL/+mB4uNeR5HvNKBLydf4AWCijcZYAPESMi6nKRp+8A4qVJq
KXkAL66zItm03gv1GpTlqTxW+QHxGyrYTbNvNiSOlksw9RAaQR28cL3pcTwJ48Ik
0TDzrAQUgeAniiTBQoGKs0X4ZRWKa5RdhAbryEWgdB3JFwC7wtXJIKZd9qTpBZpt
nMZlH6leQYNUbBoAK5hk75wd+AkOO9IHDjXcp2jnq4iz3JSV9hHBKn+uBkSZPbOE
0GlLsnOqHHtFUa9ozQvdbMQl5Szl9HBmFZ7YPr2KkMPOkCT8eBjDufbrFj9llRRK
ISJ7Q1wMWNJ4YQgMb0rnutihW9Hh4RE+MHNAObVPvixGALDweQ59EZfhib8cCMaI
O5s2sLp6A6Drd7Uw/twteL5W8sKGddlNx/OMhEhmrj2/UMJig7p8r0wD02w4iNYS
Lr1N3LYzKSRuQA9ZwvCIt+ZlwuKnQVGDlzaDXc5ivr8hzJRhNi5hPTlGXo6/rNa3
DPgB6wqIPms6eC4z9lRagC+o2n2QPLXyWjKrEqP4YV0Es5Yk3TUhkLz1l180snqN
XbJw+2iygJ1UJHpteLKCxs+RpFeByW67FFX58lQBOYNawzUG7HuV4X6JFFUJ7yQ9
gZH01jg1wNmgjf1PpQCbgbAK4erhYqFhefKeNXHQqDKVjUs+9GnZ1xc+q49JP/Jg
5m1YlITp+RhtnDyGZQ1KDvmzB8kMwCUtfjiA+s4kd8CSVgEQxIQqDytpxuDSDp4z
xo5cr5IIME0rel/+xx9XLMbcAxnkOmgikNQOtqprcEmjiwPfR9c51LnKn8OqKQzI
1HyY2r500Kg07z0EWF9B4jc7s2IJcaBNMGecnGmsc+A8yHMI+JSs5/DMw7zosKYw
5+6h3tLfWCjn+bgs4qkFr2Ym+idClwSxKGE7ReM4/RaTxYOXo1HDpN+/+WuTvkFi
zcmo+kBrPOkWFcLucD4ZMPbcjF41gCruBhWNW+sg2KVAQSYA0Pgaf6Th3aveFMxG
qOE2il86/YUeFa9TdKHcG7uG2V+TEOqnChl/qWRCO74lsBpaOZNqMC4RdBYO7SS1
xIPSNQfQsuUBIu78v1dPjLgM4TWQ40HA61gCilL4sTg7OdUuCYJsb+M+raq0L6VU
SK0PImjn1y/A+G8HZhExlbtNM6OmMPaUZyYivZaba7nhY+iiBCX9X1lwnhNrsFhy
Cg1h8whmKbgm0Z1UF+WE0gsmWkvTHfpb1XEtfo8jvLm/D+nsTG+wwWzpg9gpsl+5
cgujsITF6eA12txl9i+Swn7tHxoz0wEih5i36QCTQx6XBYSsWsY2N4SfEXwIbel1
gA4gldKNxTqaccPVvumEMVN2Zp0g4PXco/Xs0+IWMU/+KN9XSg80NFjSXUgPNJqg
ZfZ9+ddX3VLbkMamHEpvR2gtHZ1l/FE0pZ+bP3MRY5Uz+mp3KMuPDfUCcsYMmLr+
k/1vFbsRgNosqQCalol0xXNju9E6qFw+O4tPyodMHlBzWAOjth9Kupp6mYnmS3ZF
/ZOreqrUJuz8uwNyMk46PJOnTrGv2mVbo07OX5+BCWYjPrB5ZiolRcmNJUyrzDLN
WXz65E/4TDAYcjw9NoqiooHpOEZiaIynuiqTcRhiW8wanRz2OwB8xblsqAZ3zsNv
sKEzwbIPuF5WC9r38hzeJiw7ccCwvL7Gr3KQ/bWn5kQ7HJ7B/7YcIGOeNIv8pJam
wF0V3vnGf5PYb+BHrjFhpDM+2nkDe8Qc4qzWDXoyKXKzeD0oVPAS/bnbOeJS75VH
UKwQiEykA7+N6LGf7EWCKzL89y4TZ2FsW2ya9fp8o0Il6/Ly1L2+CAMZAP2O0CFh
2jv3MA5WsNnJrxgHN4aivWbbrU7ustroLK0Gbg/jzFfY/bzjYcGf7OA2TO0PIUbB
CE+3W2OBM/Hte15lr72h4/j8ecOGw3hkSTQb8pnvu4KGHJzU9c426L2IFV+LOzhV
xaIt8Z+T9BQgfTPhD7O6RAQzfkeIhNVSQt3eFIrl1szZaGuCfpoAXYi67VrjyhRR
/xovBTbuUpQFl5nZK4r3e7f3ZXH3wAOLf1W5OWJwEsGEEE4cqEEeISC8BLromfzy
S925E9K6OIqt1adsWgnpelzygEmgvOxx4duYtGT9yPeDqpF+KZw9+pOGfrsJdSsF
rLw9Y5CjV4hmt+JwKolNyYnZ+nJx658XAA6N/NkFUfjlW+eCipcvN6ezxq/K+VDY
wm77DFksF70UGrR32wawMtehReoW/BBtWma5qhRtcIw5gPqkQQWrQ8Xm5yDVeRC7
R9SUGi9M6sMbU17rU47N3iraonfLGLuhdR59gOHtAP5Qxg48ZztCXocZjwLcI4LK
MvsoAKIgBQ3PuseSjJHNvnBPLtPdKIwWnr1n05TGegXXcOVUFytqC7qZNrsSmnBD
W7M1rXAEsyEF+MEHw71wO9eAcuApalZXgSPGXwN8kO1cy8nyW0f9wEMitYQDNpWF
0qg0agCKju7FrrohFeCa97e45KL3LBUjlIcaT4CZnXZBtCc4qB9+h1AcF/308B77
8imjIoZDSKNCRcUXGxR+062VU9y5zvfQ+AASCs67Ijp+4gIriz8Hhv4wyF+tVEod
tiGs7EgNudHEDFO5iYlS3BAhkMKhck1X5G/MOG6aTRfpLGg3UiSCnkNdo2hO+8ck
tuODTlmeYDYyfmUqxPJHQj/Qui9k1RlX8bVOKLhDvlsZ9Tch9aEcP2eGSbLJxkRi
FJtmw4DrMXx+bOerQBNKD3TtlWmRcSHtpavk4fx7X0nOc42QXeNpP6XAdrJYR0YS
igRX6lYzw9bzusXUIUFZGx2+Jk1UT2fUJOybCwSisF+SpNe7qZ5Sm8f7vRxXmil/
XjjZ7n2IhIl+ulpH1HXENfe5QGLZfirRJ7r4F+Y+MTL23w0iKdy/eYBl+gWactRK
JUUw93K9F4ZQseOljsbicy+GD6GLbxSiHNr4pRV7eHJi6qDeaN3715QHx3uDfFJ8
VYFG+uaxj/fUEdAQC/yRsmzRzlP99BRBWTWRyB1hZ7owSEm+puC1yxe9VTr6txrt
Lygw5A+eBaotbvSK3QyJR+s9DFQzd0SEKBuZLbLVLBWrUTfrAxtmCJ8arz5VWye4
J0i4VY72bwmttK3y7f1+P/vgIMIFcobPyNsbzWh4ojXnFGCc0OMEJLdYFHoUJRHK
YidN1Zmmj2NahIi4cGCCRIrqJNOI9WNNSEvKoJUo5JrxbiUOvVdb8Y2x4crlQdqV
aRrgSyq0cbRusqdrNXDU/2MDz884K5EPBAMiHu8f13KwBk9gSlg1rQBPMN6sB/w4
4fXhDTdFnEBEmaRR9aqJZmhWjRcyoJ6SB7UWWH4ofzvlAjoYxoD8EiDF3bMH3HfM
omy/aETB4GyHrBb9tCDgDwFEYTTGvT/bpaw9lgQzdEVCunRp7XYf6aHpzCts3jP6
3a8rqlAUBStIvpSFhul2aMJhFxgnXdiFujl1l6fBvk75r8xrZQ7WoTk6/Q1nFFFF
wunjqRunwmovvuDGdGN/WL5eUeM3YF/uSO9IBKILuH6Aq7wjMJZKg8OB2iFSQDnU
mMhETGr0s0+ZSLEVCRFpRY2ulGKJ9bRhP4oUyk/tjVAaol94seARJKYQ33oTSjVl
4oEuicLd4fq6WFvEyMTzKe+CdCVaQA/ReC3x8F9Fuy9E78x6GNbDsy5U7VMAaGRT
wLxa+vkCMG3WJbJh3KS/XSHbnN217gNfrGkXF7dc9ufc2uipO74qjjNYbOmvViO9
Y/LSA8S14zG/Z033EOZ9d4g4xPTFduk3i3fV2PoE3nd9tcZDzouhOkR7DpvtqGsY
ORXYTFYAJ7aTSz7s9BbP8YUwZnMpMpbzZmnIFNDIexuoz+hmBC5yuJ556sYrrvC/
fHku5VFgGLpaDTP3MzlTAmyN1MKLV2R+nx/haJEKyEgU9wfHcjkAVjqAX3o2BNiP
X4JvH2QApXCVnHPtz8yn9Z4gQIUHzwQlsa/xs0ONviNn6I2sUNZ2QiXkekrHpcNB
lmcDNSxOfjAbwoo8y/ENRTVycfarYWxpxLvp0jzAO0z9NU2bSQ5CwBGwh9hnXGSo
hue23zqg5UCbqESCSSlWVZt++bZnhjmGdb3Uqe8k681N0tPxNLw7iEt+PJtlQUwq
QiMlv6lbnr9WKaSb0YoUDv6qXiUnrHw0PY7jViM118Zdt0Dt87wdc/9fddBnBO60
DjPlkSXhQNbpbTwAqWCT5A74UdqM7r9ejUlSFjcIP+rgC8u8W8Hm10MgevS9S5ME
i/Aen7qiC2zYtHFMj+d7gcqzIe2KS7sShQ2dATFBEM3mwOh01ymdJTiMKDPQVTjN
zqExEYyrMWQjnrKf+OXzZid8mwuvArYL4sCsUnN9JHxnyYxR4rSQVOYga77hXThi
I/U3gY2K7zGIN4fbxDgTzNdOEyFAQwP5ri3N5hoKqpi85uibkbAUFR6Aaa6J5+Nm
dsaKnGM5XGii3Ta1j9VXiU5nLzjmUXp8XUojdyCDpdbvwqIotBxYqnEU/oA4Kjbs
93uBnTMG91nMPZplJRL/SS1T9Ciluj8cgD1lLQAI7398ePRzKMuyQD/3K63Bpb8C
EO34jVrdrxyemSqapfFavtYP3Ec9H6sbwdlV1We6DYSfW4yPHkIWkfruTZx/KVE1
36/izsLSlQCKf5lcYpT33hdveXB098tJOSmdb3b+/Gitgp/Mz7oXKCOttSMWSu7V
r6XrYB1teBeBfGoW8kvpFmt/yEaYF3oWLU4wK57d1hNiobKj5Be6Sn23J6xlaw4k
EjxgMc1aG/dVWoDF+W2LMaNyAzTfBIVGL5Zc9dkvQAlQsi+N6A1eZ89y1uyCVAGa
Or7sfWBQzWD5/dlLgSTau0w/4wFsp28/deXiSIIW5EWyhMLOwMP/xUOFDaVcB5KP
Ywu9mKA8dhL71GFoHuv7QyAT+K0GbhgzekAaeqcqKK1SW7DyjrcuKIc0EsR2Bftv
n6hrgYyQ4S8KfPFn7Ei0k6Yz78I3LhhW5grJEFyJcu2iylzYeVXVOZPJ6CezsKaN
VVdFALMNzTYFPZFZXys0CFlO44P2nmWahWC2R7H5Zsbr1Yp/2M6KQRK/d46WvtnC
5+eAlEiWqgOh16qbSkcXJdwDSfFKA6HED/XMVubmDM7qDwJSipaY2Un9X/Kozb06
BmDmoPJtW0Lv4NEX08JxjsLQ0GV/YyWjM6K4V2l20m0d8OOCuIyxKv8HRCYS66Xi
R2hAgpWJr7HotnduQhj7P9PhKtx7EOESa34kDPaOQOGp4xO28mgmTR2WV0ZLFWG+
A+uF2MJAvi4/xz+aliY1ukDCVh7+vTpq1DkHoDkqsFNwcgR8T7hRsNqIjIzPnfTw
9uS+20vYXFQIIFQ38WXMq+OEtBHVMgExCoDR0Iyr2jnTpK650p66+E1FfRzTqAWw
VhziUoeGGVkFAwRTF002Y93Eu1yjFY1ZzRbsa8dZkrRB4LjfUNapram3+sbHR56t
RcFz/E1hUOV6LagNmBDDGd3I3EpcwqBV7M0O+0BrA3qxGywE0sYBNMamuO5CEkQs
eLgGYLctkNA9jjgFMR96fFk6G1JgfncqPCmo+oaevIQXYtKlHZYoq0q+SUPlwhBr
3PdWDzHIYk6GHGpswJwOd0XVM0Y/wuYdXEjkMlYk8rSVA5TsT7edUEhGoy3gqykl
LkBsiyh+wUGur9vAWwBVK/54Ff1rhM4cDqCVFngK/NoOYLDSVvROhvfyDUW8KDY8
76t5vXUCseqfBPlopog0XqGtNmMtTIhF7yW622QuG4KwyNFlAJ+mFJ9prJGdybP+
ApOw43t9FyuMavp5jBrXcWr/NpsNW1MdzxCUYLz9YtGk7LWFbODPywws7YUaQVLz
4VtO8QlrAckKo2Sji/9cTocF20BpDduPNHPLG/Jzw8ehPpCuvBjC/6/g8wVTIrYN
WLrclp196hd2EoRvjFszGur4ZQX9MDTmNp4pMML9WE4b9vw4DNIFz9Ax2yOBvFuh
V4BYaNiJ/BnCrUxiYdsJpdxjo99cETwuCGpia0YI6IdHE7PBzyLM6HyRGOK9ARIg
n8knXg6eewWMf2YeMLhHgeatOEBBTAW2iur7psAVavjVxH9ouJf6T3iFg7loIrO1
q0O/PutWr/f92KzRMIOYl7DOAKX485Y2JOJBonjC9+tkjTUh1iWn+iFSUx21y93o
dRlTphmTNyT/QtT2O7bdWI5FoaBq7BV1B0BSME2rmJxw/jfqUH1VkYVbIcfwLouG
Tdtaz/Uq06tFqrdkqY7JfxEZxd5+7S87Gxq7ay8m/2J7BerDBprTjU9lEIv7wrgo
w1M+BKA/rcFL70/3BD3ElQrG/EgoUGWxLuNp0zzGjCa+aLqGvBniKyhv7KIZFkoY
804jEUsS0epHFQCtWyHEUtx+zIuGl9YoHTOxaLc2mnEkF3XQNbsh/eBr4y2O7ncn
CxORpqfWzkT7LvkTT8WP2FbnPpwTSQN+gofb0ZvPYBIE/szDWs4iWaq7nyjtBOhc
NLW3e1B+BJkNqLgPuyP8wQl4CIR4GLD2cLCWRRoTyHchBcHnKhMQ+tE7V2gi+L9i
t088Y2JOjTx21KTlobnbn+mDGZXaoo+QwAoyKa9tvPcRZ0HVptU1Vu4rIJJqP6nk
76VRPEtwGVZCYx/7dK3GcWm6fUThQc7ZM5l0L/R9b4PrNICslG59PleBwhPYuNgt
5wCmkTRe4eERBGFzvyv4wq2WbfppzwMeNgPphfmLQPvL9/u3+74nNCW1TBVBFtc/
clPjai7ww4/0MEL/dq0RxTzf+P2/InJu33Yal3UiYjtRKJkun45JCEXjzDwmiHDj
mYHUe6ol9EwjZTp+tBdkOBI296nZxXalfmtLcQCUyNupYBnKqjTyQzXgj/qcyKqr
3I36YFttl2OaO+1bloSpLzsj5Q0N0bjEoNCvUsIUQ93wGFOqZPIWdwiV9edNYWew
dZJJ+gWXswvcLGo+ck2wp4O/jJG7gHP9xyHMUl0fQjNGtX3aLmlUjLTbthiAp5RH
syNYiLy3Kq8FXlW2sduhn8MdDBUR8YcNrfM3h3rofJFfEsLfvo3Gq013aRePov6E
UbAmQt7NbB3gZTYLbZ2B0D7JU9f7yZI6SZCaDofvEqYqWgPPQizCAdasgtTlBlIb
Gc0qKb+wP7l03VzSYOju+tR6VvU7crigZaZsLfGvuT84TT7+kdR+zNvWq1RYWm7r
y4/j4GhrvHUs2tJxD51cBi3AWVVgqK/9bV0g6J0KJca4zQ9r8WX1dvQutHhEoJtn
r7xbcCgmx1OtN300qNBqujXWpi77Jd1EovNYmLgFy6BKQhUpD5X/VkRMVgFcM9Jr
H/VGiYDrbvFIR5iXv/lvqbwanl7Xh7x/N8o5VdUiJd48p5w1z1qj4s67qE42JxKn
8kJz7jpwGkmzAORSRW+jwxmk/eLl8e3yCp6E/MuwCrp40JlUJIRRwqA0RZAD9hv1
/tEw/azPaiUGLcpPJLuekUcGeppmNx/T5Ih7roO89VuKAWN8nByJdFruxar5vmZi
6Cq0yCt+u8Nb+BY5jT43jXR7ooyBAJE3c6E/lfPUP5R4ly1SxmNE44mlnlMJcJ3z
jQGo7FrAj2u49H4i2nfZfW5kNVwoskgYP/kEuDXRTMl4iKh0jsFcjt4ALX5m3CUN
225xf0d9PvScGxW5Ce0Bk6np79lsaIhCElOBwJn6vsLuFrkMY7BhjnlUsfBlzf4D
NNRkxPXi0O5upEVzFWYH9TM5LGCLO1hckRCqdwvxgGzluoz+d8ZOWVZ4whEDPXka
eg8YK4OelH82dYUPaG415sqofQhAeWOZ2iLJ0nL/yyGCI8xO7EZjVhKF24S1EQWf
EGdm0NOULtYoQSX9YluJw6pq67Db39oVsO0gXgScmFlZecRxVSnT3drMZtoxnLDc
flsDWDA2If6CtNxdvGadOcKfaJRKeyDBJRdisz1H4AlKITFQSaAv7nBAMiL6m0UX
08MgLKP48WnHF7FBpnGSUkyRk7YIe+5+gpvTs4rASLURE6tKleJMUMoE/uQB/LJQ
BRDnkiZtaziyKBD0X/wFK8FYIJmJS1Kp1s9yO1t2DKrM+QLUSVOiydIU9RdlUB5A
saTMozHZk0tmyvPeGOLPeQSCMlFdm8tbfOKT4iLNGWVW6F93aOiLh2qE7o+P049N
CtR6WRpRWf16gWvvPfjk+sM9kfEFbSVn2M+VGk3OqkwKOCkRDezzeM45Vqbh68jv
ZYhOoMHaZT9Yb+sV+hMqnL2K7iv3ebo+Jgn/BbgKNmWMpl9mhsCFMMI+r37A8QE1
hR4Z2N/w0HIi39L5dHEsX/qC6TDtOBhfDwh6a5dmYuaVVyAob2tUBdHCg55D4XFS
qiSfuWWk2NUKY/42jcg9vgYOiTyxqVpMpuZ4Z3VoMhoGPXxZIKhZHzlQGWgFkV+v
DRLdBNsFEXcauTBXmLvcSPUTpjEUyzVmqDwXFf4+HY/vC6IzDQ2j2EON6cJitqFA
Q4MiU55koQW522VgGwqn5ucv/1nvTnKbVXF1uIp0xgBQwil2oFkMrLhlge1gtYgp
c5FCNneBLIpK5LqwuN7DPCw0HvXJ2/3ZFVXQvGKYOsiBL1CyUaTUtElgGeQZQPo/
phL6rzFJKZ+wdLnAU7ZwhaR7nMqy4NM0rEYbc+WYkLmk+5H5uIX2qeR+Ai70oOr2
1QI6KIf9ToHDt8OCtPmhdr7a3b2DB4emb3jUYkMfbL8tbJOzmQSiBI7ECa2n/qkP
XSwQky4vs4mK5DncIApCAFrv/33bXto1iqVPMtAWF0pX9aRyynZ/XrErHz1M1Lc/
sSV0gdpgh86OnVZ69+4VdTagP+zvV38eSqWnfXkk2XS4t0jX/SCxRq7xcwU3RyDR
mVYk+QYNpNO17koz2Q4RPLfHYbZ50GsNFXw/B4oRKO4SZWzJoxDDsx6kBOB+Alcy
bW/632yI9nwc/6YHj3rLGDGXlxOGQ/olsmbcLeIdcGYNlXZqEr+hjc6OmnfEs/gM
PKxPLr3ME2oVXc1ee8yU4f5xeWkB3fuBvKm0syjcnLhFfTxOy+mFvnAWMKXSzs1t
7GbqwILepVc8y+5GsGc6Y7mL18Pb2lbqPsOlIeQo93wYqiAiOgUqcg80hq1I+53Z
AHvuOBAbrX9+V68hHIJTTWIXdNY7XfzDFBUEVbR+ev4ybmyxccshqE/46VIi8nJu
I36N+UjW1hKoN+4HlIJuAI3g9xjD4RAX/fkO424E0yXEnKRJhqitYnJl7SgU+ovW
fDKlVjU+I7vZRtYww/PjK+a6gVdhXCqm443IUMwGjRpnXLpb2RjcfPYZ9+K+7ffu
xBr4BRNjQGwA8svY8AJfC0qLWewWDEMFfYDU+CXUM1yYf+oNNo2HUZbKHUWdn6yS
Qy9BDqn28OYak/q96Gjh2xz8uvrviRlZglYh36VndMteHeWK18d0UU+9w0YQItCh
+7+HwhY8xLtGjVJA5fYmE/N0qesGD8K9AgQWJtMBlEqy16qtvyWuKsvFnVV7k0ry
5PFhTKJQAl05SLcODOc0rpN6fAs4oMyxvM21n2VjTbLr3XLymEj7i5o7N3398oIL
UipxY9gj1GGth+ur+2aPdXrQ6JgXimQMQYCLwGCAZkPoyvktpy6ZBo4zJoaqsU/a
ykopCakxGAo2L1+uwaFYqAb00x1dmRYHfb+vl+etd/BGXfHWi2qTtSjuxug0je1n
HvWmoTLcctU3NiPYXM65XzeuqFStn61hLq+9J3Q271fAOWJFiOt4FqOT7lGXYX4X
PP9aNVZaFBE1fKsntVW+0XhkgZPZ9a5iONpH6MAuqJRt3CqnvFnlD9n3qzTeSWBm
UBH1Ga6VAotXMJwmrdDQcELm/7YIjYncakscGMUhRW2tXdVkw1jnifRZdmMFE3Xm
Byc8kU5FfU0sei4wg6fEhMgRdH54fw/j3PT1jem0j+0pr74GarCZtnhtNiMtfDTH
2KktS2OTT+lsRFtOwy7gyUtFm8AR0do7zjUN6+1+0rvVB8IUiNr36RdkG3bpqBEm
ARLvMqUN05uWxCm+kByE0s9txRv18INRnN8g/tg6BwqlkcQveIT9XnkCJ8bUCr6S
QOr7eWd1i8+cCgG9IYVu2EFSrXFWf1IceWC/DO/XxB87dFTe/z9UVh/ZGMg0oRT9
jFa5JIhfn/22W4SjKtjx5UDQA1pmcIva5W1WlwC5vskhB3J6ab0cQvpkb6rwFzcb
mlkh+sNwXD6s3RX8cXO/VteFH71CcyoxCN92RjTBhregcW/25kyQtV4Lk2UO18JG
c/xFb29UCP/LrfnhmBwISsFeI8rUyo/Ci4h6Lms85qhGfTnUqfW3kuvNNEjFF1C/
KIWAh/9+okxSyF8uhIwhYboViLpYPELDjV1xFRPZHL38aRPV9wBfeWhEuOkvEhlv
wTKXwQHMMN4/UVikMOIZ+9vpOhx9nQDFbB22nuY7qhcOnLLjNup5YekGhYQQrm8q
p5ZQJuBMr+XRJWMkMXCBA1f13ikExs9VFM51VFnaXe7Ui1T+Mz7/mh0WNsqD+8mE
41dCQ+o+MTH2OB8OHtMiktD6Kp6oAt5pEwB/Ay0AGzFgsfNIAUbPJWDTvUSSPZ0V
m3v+K9qspZeknKNBJnbJ4klzMl9fCZo4IhPMFmDes7q6k9TCbbxzRTpBIkpP00jz
BV+bhNCpcLmM1lTsTm8YcZrkFL/P03HvvPKK8shP+8oyNpipHMimpTQagpbFSgZC
QbwzKpXeAGjoHN6/rkLWa3US025wZI7Ry/p45x6Ssk0snNKZo1tfJl2FclQlpqZk
MAZtaH4EwiDJmqhe5QByHrfosC676g7GBKb5UP6vrH/IJLDNSOV6ln9sxXPYQCMD
hTwwNIaZEo+gVw4l6Xyft6emrLZa11BYo0HEQdTTkR+6Spe/uPS1ZXd2qCFgqQ3o
O38Ouh6aepEC1CC71x/g6i59x0EaATb/+1pK20F+t2LiuscSSKKA7DaS0AUQXXmH
0MTMGhMk+UAc9Fik7IkVGjl27abpLBg6tY4xKs1h32qWEHOT/XEe/oBlRczl23bO
1ahspuSV2sNh33wkkQVHA1Blz8UNl7b/6LU4Zl469sjsKqZKS8us7nWqpr7N1mcz
WJbf67he8/zot7OVThI1JvtGbk5cQUiXUE0jWVd/oBEOJsg4+32X/andVev5s784
tUo7rmoSxTMUycldbzIcDff98jVG2uX+HLVGwSNmN3vHePn7Iy+gIK9RGdytUDza
ksbvzHFejYkjpDjdMzX0j/pqiEkaFq/z89DM+d4cWO3nYYVUXxfZLIjhWm9DEymd
jn0bvCmov1Y3IItjW5GpXaLlSrqdXNuQNkM69EvYHsttGpEOSiBYkD5ZmejeTex+
7Q4EYHUOEho3/FPj6PrYO4COgW6mnPjBzaJ+MMvjKNiKjkNJviwtO1FOfIyHlT/T
q16n3Yr279pCnOuVNJyfCojzjeeaZlrqEMYqjhkxrV3KiymYAxg32CC91YY9Z2LD
Ms0mTF/VuX8gSp0cVoBdG4TylBKCUG33mU/qCAIklgGV72iYWOJkG4PqGOwYFpwV
Ks3TNShttoeGH6ZcO9S0A4Z8O4p96DOfuLJOKHN1W5+rfi4PKyAc4D5ZWaBCAbad
WyCpFf55wbTNKp10ZhyQ3KPJ5HLjd1xoj44/8t7AmvzkSt5LrO1NKkYWnTfyZNT4
1MqIFxD+pNrOD3f80VLwDYCE0HgL84lahsmzcpycwVyX+Sg6LrpV7K2mzrvPDnaA
s6Eu6ON8vM6t4wPb8GFvid1IbT+WAV7tkaS+AWJmvm1KQpGiBgDapAqDYOdBSRsJ
Rt+XA/AlSKG53FxONEkjoz3iuBHBzcuvZXsLw8IlvdNVamS/lqSDCdaCqwM/Gi1l
4WNw90pFAjJpSGYmEw8xqNUOGsIMrX4u1Z7FrorrNseQv7F3mXvpeRQO5F+1uDVm
Kvl3WHUp5W7ZLySfm7DkEq0MMbn0JbHwCWOr3COou8CvrrsD67kWLDQ95C9Qaozl
OwIzhdBWSjwlDUmhVMhJvffubWjN37RSOounZpy8cGYDG7Fdwrs5/Z44zGH2WSwL
UMB+IJP96ICQmDoljqf8U9fe1o/P31t/mEoseL5tvIIXL965Ji+pfRAE65Jk5j8f
cykSOkeZjvSJoW6Rz5zz1cELE5ODrMtS6TlK1v+oHw3ZbpnVYBby6MTFAh/QmEPX
wwHz0GH678ZxMgDkbywmA8BxHn6Dm4pTrCgsabCfaeeM3zYYGqPzW+Ec1S/D4Qlb
pSUbHcpfnRsMDPzXLiSaTbi7vEaFp5o+710QpSYkoOh/d+E64aBQn6B1zSjz8bsO
xViYDoLhbLidLvbmqEJGICXtFPmDgD5NjgMcmP27iITR/yW87gNVh28RTFKReiLJ
LlgAF6HwHr9vsLCyDH0h6hcNirujsh4uCkcECGtIYPLWL5C/HHNflHlWrRqgxFHm
5SXm3YyEWtoEJb6PtlaZz2ZhFwUoE50FQoHO3J8dplDtuBvjeXdJ6lLWBDcNjYfa
xtMr6Qrg6DQLxQ/ltmbX7Vvh6jOHb4Ccf1Sx4vEv8EgzsCSry7X2Lv/UUJA6GwoD
Q6C69Fl8YehXZjq9o7vriiRqk2Z+DTObswnQ/o5/D9k2NUzZKMkTfL3KR7MyFKw7
6lBTykJDprZ7eURbbSvZtdPykBeYhooW0tv2kR+3C8WaXBH0JKmAuiZcdMcdzfnl
U3HA2V5FNda0vU0ZayWtsaZ4nwDkgvjuygXFb8nWNeauem2Ueev9Sd/wK/jw8ypu
dMbCBzdY5kZm1KKsE5H1u8qWlKNA+i1wlZ+to2D1Gj9CXfC5yxbGZ6Rj4I/H9r5u
dg6AwTFocI4VM7/8XP4icXyopR5HpQudSTBoQGIAEaWnqNTmaLHYfRoVWLpxx7qR
TGHidvrZMt+WSJP9Loe9RA0+seAZBJ/UeaUhrhQcaQoAtqZexvlpHuJT561j9L1s
Ep4YGtM64aP5HAnz1nh4NgfH+h0grSrZhZ4rkvgaxiQl+vu5ePq13KEUbxXfj/6Y
ggkClT+aplHyaWbZrO8lMoC0/E/eaI9q+ZXdleG7JUv34kxMb69oJo4Zq2M2v4k9
Hn6qEWCGvGCfx7hKQN6vRwayOFaOErBtumH6qPa+lw+gqXLdEWXDv6+907aIV9rb
JA9UfoMiYiPZur6O8Vq9WwtuHkS63gcmvdWgzA04pgFyoZgeCbj7GelOqsmBhk2H
jEIZoSRz1iulVWDpyLRgy0pwmcnkuEe++EDb49UefNp1GvUmLcYHsp5C6LQiyHzX
Hd7SmSSm5CGWLf3hXqFQY75MAbmYflrjKo78dwPGWuUxWych11eUjS3elJTsOPjs
rEUA6qwwxLkXiy0R9cSuJkJEeM5HGkrGOCF2jB4kvfoUzY/pLXasaDv6a8PoD3g8
O3y9diCmBu6XopEwgRMOke7u6NxDbXB5oDpya2vwLc3oRU/dIbd+iTkUkELdeZ70
vOK4StU1fFxYzeAwgUJFSfFSiufiHgxAj73dgLwklowBy0IVZ6mr0RIlhnZR/cOl
CUmGCfo6Id5XtOGG8SdPC676ZS3DJm0k6Qmlh8sRP2xQ4yRcb5YDM4WHYjxWnXet
RCzJGng25L5/pV89MC9fw94vtff5bYAov/xPfxuBMWdcFH/B2yqcnQOwTK/EVCU8
2KIr0d+gWb00sNRn2ADdmRwHFOrzo4JseHGDx2iOCFHi9MPBMM0OHB+0jgXSC1B9
Tw/zHeqeUIrkLznfN5SiZNcE4ewaNoP5qUtIyKQu9jO7i7iQdoIsjdu+p7ONwrzF
8vCKoL0UPe71zGdYjo4oxpbT8UL2gSknNJBcpDUoScBjHlfl1HVbykt7dMKKfoNv
/IvlA7Iy0Hx9Im0bSR04K2+kUNw/tC7BDkikbaPecIZ/jmSKYK9HaGpKVUA9CLPJ
pXfJdFEk8pPIBZki2kUrFk7/yqK9AFVslxRglS9AYKPTH/pLikc1Y9/NtV4k5bHv
URmpEv0jo37qd2PYVnaqK4SC7B5OOlqY+at3eHkV3mBmPtBPbQcVH83OlQa8kgq0
DqMov7eTjSDEeMFgRvyJ2icFBKqEMFLNBkDtMG2LKdMznaiYT9cWO4GhKYaKpXX1
s7PNGGZwx56wjgqs3ihHMkUNRPsKPgdbuLopODNYWuLKafOCR3a9Q1Yrwat8Hcrr
zfYvhIaNtV1ASQv5WX9HtZ/hyBa9lERciyPdg37XR7SRZSPzsyaxdaLZyUT13Dev
Amm0oCJ/H8h+pm9WEnjFZN2HMEcXyrBQIYU9q+eQHO7Ja/XL3wJRxIZH+mEZD995
4wbvaslidnZ5zeNfd018V0Z2Xd5+WtRoSQ12pLMZlSUzaXrJUjbFXAwjXlWnRz+S
w2shUr8BcMpNwuUvzlkQS78NOS0mHj1TnwtozdIXG42pNyGZ/riVjBKjdYZtcthJ
JLkx+4yhuJn5D5nl8I+XOBwcrCFOs0HwGxEDtUtihWSufD2hhurXLKk1rEsMt+Ym
qXT3esEB3lVOJil5Mxw0uRoNlz95qqaWrgXiaIA8+6wdiTj73kzRbQma9bFgb+eL
JPKTSCb2YB/OQcNZU7BloV/LFk2rxOgaU+T4an+qSvtArRRO4EASaoH8BUpLH4XW
Be+dyQEsR+O413QpyiGkfO2IycdfjXvCy1HFcsb4QBg4IAaPFr9HbhXvj0If6czm
+dKmcvV//UnY7QiSgM7QOLLUBYJx+kyqyJUHTbGQqmNgXNozdTIhza9Dm3HonVuH
vQomL3Ecsc2ux+waoCSlMyKIXvXoWhc9O6lL7gOA4jZ6aJxqIrbFAQXOvbq0jgS+
q5Rkd99g+T8Mwdj+1o/rY4OcIXFXzg1bVaUivCmIz8r/wDPYG88UdD/M4DDTzUU/
GytM7BedDiF/pVla8s5BCGjZw26xzpIgloraZjCOFArBbaHc3+B3AKNfcCpOYXab
d+VjUNrDOZ+dLRBYn8dHZzNBlEAcaqHdkOVgP+Dwnl3MHxr+U5+0aUu71aDnj+XC
xIyK1n8whp4meZlRhBnxhDQPjXQGVXvw7YH6FRNZn/jf6MGu1rrVOaN5aDrMwBJV
PvKZxgOvDRkkmPq4bBcge2SmCehxv5FNBTfLQoq3k73L2UKtFZ31DubdB+uI6cJU
umQ7alLrDv/rGkGuemKV1yeROjXMHqEKsvr2bS8g6sM4CRwniB9XoxqzYHLBrmiP
o09ImlJ/q14CKPouO5Q+a2xB686Vip94Ox6TUHQGodUaxsGhXOgVfmeEOnG3fPbT
lLz6ugEMfUXUMfSvOMES5nxV9vJgdsPi18Bub68jcsUEufegSpMb/4z3xAi8Zw9N
HCYpBava7Aia5TlZH9spA/FajSqVi1n0vnM/qyLZdkdJ1ITjhKhgXSkvyNIOf/ZD
E9TEQUNP7gplVccDn7r4xdCDN3Di53t/i/suo4fn3f3haOwPoAQ763dMX92nnAkF
vC3z2mAjSqxAfsXWAg6XdLEaGZ8rx8PIktzER/okDUpvocfyZvlc8tYDhIEUmDtI
dCE+6hFrtkca5SGBXlQQkCoLo4YGa4610nSsGt/MD1vqaSK3SPyO5MV5LyX3OEEb
TYfwzRQ6mqp6Ztjb3G9i5IE9/8oP6ZEmWcUsy/OmTq2f+3fgHv4T3o4xQFqVn7FG
URqltQ9PLHoK1xgj9zV3M7upzaqB2YT6fOfV7SIV7lIXkklnnnNbkcSypcNupivE
9gwIXuW73Z+BRuWQQ74h7aNeSv/X6HtOpvqEXVLEhbCRhvad3lJo2nkUfRn0U82D
x7Z/kd9brQr/SMmYDZFCV3jUxn5xR3rnv4U+y4TqUAXB2fAo3/yQwb0jNalZmRxi
Ad0VhejRmRhLCizjZRLduqmdHJQ8UJlldyE8H3vXUWCVHwQCgCBKW1+XSGsEywXQ
hHQ9C8tpWnHJUf7C3SLQy7UjonJMUPpXo6u9ga1w/2LB6eZLCJYIYzy40b4149zq
TW7Fe193bhw41ldHntt9FZQ8Dmbs1v1UQr31z3fefFwE5t7YcX3LWS7EWBbH0IE1
BxLX38LnShwl6UUlktFmcEyVDH92UYNB18N8fyVgHGlOzpCCEnYRd8+iUwq0nxpn
Kj5scZj5mV4IHOod+8Ktj/+aASygmao4oiWMEQq5rqdycj2X91ZDVtkjfyF7MqNI
2roMoYlB8LPwSdBUYY9ejvf2jbBM7WKXT5rlj6kjCWFUzYT+L+2zk21mCq7NA4d1
tiTJ10lDVR857qRJ7L82cHui+AwDWk9DyMN1wI3YOAGFxp91zufv7J8OtoS9FTwB
hDlw5LAjVGy5Mf85d5F4dRHpagqEgoT520N0IJujTGZ8OPJ3DLjnzbWpvJVOACNa
xtM60teELyjStzKhOhztEtn0nt+WnksCD/ZhHNKTODiMzVE3m83yE6D9J/V94XQ1
ZMcRk+mlgynek9VCxi9/zQNPiQ+dAnI7wvQ4nEBJn3FyxQcPt/yyVHXeho1HFwUW
mJAVMuErsaKk+9tbFH7xMsAYpQDCeAwHwGCOhUwCRc2tX7ikbLbmmlsnivkbSV2f
AFIy/FYPOkDusTzCTr4ZLuCF9THRL33uJV6rPylGdXmOH2WyutrUCOFHjYvT/Dz1
8syHZhHgUi5BPqNcwnj0rlGj/mrvQvnhvyUs53KdIjIxJKGpBqURy5HAA8BVnN2v
E0kA6PqKA73xy63tlAH4br9MkoBN3kU+YoL3PrbWGb5C+JGrSpTqqrLG5l+IDQuC
zElwy7Gys6vZzjzLpGzgh61nlmfFahZAFRxGtxN+gtOmfSBLxWmhLcYx7/29do41
aGQf30R1crjAC2beYeiGxzbIFVD4ApoUCUc0scEO1JgcUunp5auvVJ0WOugz6p6U
Pr62F5y2Zbf1RKK7fmfQO7I2qOREZpBC+imy4/uQ1o7htmLSjz8mva0q6RTkXFzD
T0TwqkgfWLJCbC4jCHUEmsgHMGf3mAsKFAnYwFb2mmk5s87IG9WhGx9XizyLFPix
4sxrc5aWtSYaF7qOA4+g/luUh9XMHJ1VTLYRDMNikrvnURydt3EqgY14Xkc8DGd4
/pAjfxH2e9fRLEuDGgZZxMKh2EWNKtHoEx05b87ivJ4o20Rck7JHB3f84yjT/3bA
1hJ6uro8UyfGcU43P13m6iiad5Cjh9l7KL+6DBqW5UURtgqC3lnpD2GJFrokPP9C
ZrbGO1gzPvhGsZYWjf5opDOXDvoaJzjfo3zSlKDzqJX/IBPhLEdPW/KlEQy+c6cs
WOVzQ/J12do4vwmecMCY2QGkFNCP/gCBSbfW2E4Y0xJk9Le4mvlxMj0DHznpzDIz
JvsPkOVcK/SLcFzLHmaJZ3MnzA/AlUOVZzVKbk4qvAn2PJuPr5ribNFJTFfgfhoK
IbGHTGops3gkL0xLqigcjBM0C2MuTdWJ1fnu/xkrIpkGFmAnoXwHmKR/IF3glmsK
lVdOFSAMah8i2RRTZe3d9IwJosAuOVpVjQfMAafJAoXcHILEWlbgiWIT/2PaBezF
Diyu5cWE42Yl3GkJXO0vLg+VmnggbDuabIj8n08oi7WvnYQcX2g7nwNaT0ZXb33T
Do4YLObtHKCcvFlqFBMwf4s8IhCROJNoqEe4XFU9Js/7Qf2813WulsW6tRnFUxNg
+o0rpeKI6W0OKvaB/TT+kDylCeWIzXfHeSvx9krRabR3bTGjyS5QVg6oORrhPcp4
QNHox1atafRpVGwdl+p2/oFC3a+R3SGvDb6ODNQMroUndiWK+Sw+KaiWOa+xEOxC
qfHzfckXPxQDqiR9juETiHYS01/NLg0kzzURYKCxd7bx9EVxu0bH4+2Gwtpr/mad
7U8eHEGhGN3TXBWH0UoDZTcjXCPA0LxTUmnsVF07kEWPAsprLPkJScMCLSlWMnVI
5qi052l3Cdcn5peJokD00SJgVVbNPOlWB8SeSNfXOr+zV7SGa/zDm+CUXbDLR+Z3
dcIhzjQKcMZ7DtMRPpn/gWaUFmk3x2w7ozbMad+duyKIotpuo5Kazf5RrKBe31nx
7QQUzO1A6l+lvcPNey/e/Ep79of7jmjOrzTLAgLmJn6r3xlEmdTkg3EjmEIqcjft
WSuagr+w2PH78v7YBC7aPQ+SZckmW2qo2JHuy6iqZ2KHgGuVBc+HFxqutWgxjYBK
V8hD91sW8xRcUsUaqwx/IZLwxMEmNqUu5XUiPHLoNlTR27JLaEgU1oVi/Np7sErT
v6wZFg2nH6rD/sqYLgZOnEZu6PS1kpmfS+iI3QytdquRw5J9rqecPuB9BrEIgNT9
L4hEqeu1S1Purd9h0JGmBkKe022MxyMvRxFevqKBTytS+RmL5rq42rBhdTqNepZ6
gVdYJ7tI75G+qlR4V7MqQmH5S/dSG9M7y6mcU4l3qOdOKCy/Hu85ozZAP3idRaOy
e3fy7ELwdpcunY9TYMEfvUhiPWSDQAPvS5b7a2sX20QH5x4hlYHg6nz29QeJHiiH
aKkxSsUWpmbqSBhIngzr3HcW6Vr5TgHFXiPpjL8PzkXRCWkxhtfmy4tC7inh0kOB
uW0y2DIyfj1LoaCY+ApDipVV2lZLSvDZEihekCCj77udA0tpl1RMUJFXQ3g5/KlZ
pBIzGcdlmbaIr9TaIWCFS6m8Q/gtoYiZPyVDBd64PpHuVVAB4At8KFseYtLBTGtj
ZGICNDVVkvNdQ80upWkAzwmRNvpyKlpUjBYhE8P85AK+qprB2IWDbdEPYpx/fKcd
kc7lV/bsJP6wa2UyIFxqZceHrvAi5ssgemLMCdztedpkrSuPtwr7E5/ibqpD/uaB
gmsum8VyXQBWxZWlu5/ACSjn4Khx2xkt0dRy7g4LQgGUhHdM38f86U9jxv/pvkDw
etEP/GaHS8vkXxhgcRCLOCLl1YW3qDzl5rZU/RE1ZdOS7zoxMAe4dqWYzJkv+Iud
X6fz+BmtOfDADNB4UhnHsgkhVRp0vXcytC/TK688+OV0dvOEte6U1twuOOm2lOcZ
/IAp22d5gp010k4qvo9qufydqc+RzlHgco2K3NHC3mG6gLRdm7N/PBbm6LQvHfSg
sFTm4QwricQyHm5KvqQ9iThbP9TGh+WFFO6v6vtKlFVQnYRa1k0SpONewPNIYNU2
lSHcWUhTE4GIDjAGlmCEtJrMk/i/e0CcbIXUER/3kFmPGUHNURXZoHEGxdW5MKih
cDAsHzXQhoSYImd9lcWE1f5d6RtQJsr8hVCkrw6Ujtyy/SLNXcn1EDLmAtaSMtsg
nDKaTqgRNlRsSppxdlGvSa/WjNdZ8wCISFFQIRyWD5fr5NJhHQx0XIozXKgsU4Jm
Kd9wZ3DAsYPT3h03rKJFR3t1wjFe43G2vlR7PTeYGEa3B8Tv7xNOijfn6YzknF1X
L5Jib9AvZ81Xc/60wDvFOyYEWVp0osj42sLZt7nfwsvRUenxPxtR+PYWwkSxrBEB
RDobviP/kvNX7ljyJsjS1KjQRmubx/CqO28YaRQMKKnM6YnWu+xyvVuy1GZG8k8b
J4ql+2xEZt9+85IkMDjSzurqWXHUcajjoxPogL6smHCTOy4NpcNYHsnVpejfi5PV
49ZpdZvlx2ZYIPZqBl0YJ7GbjGYifrLRjkA4F1MHl9JVQRCRW1TE5I+zivnVZ5xp
C8IVJ/gzgiJS1L+8OBwS1hpAZk37CF+p/RSmrv9bE1wqmZ+NgG+rkSfnVXcYeUub
drap6+5NByWEDLaZCQSUSMeEtzw67kkmk1XTm4oFTvvzFzpNGCideUB5o8H36fL2
ktn6OUWpid8T1Z4Ka1qfCyZK0lf7tgdDycIRxSV9ZzTtnnCj8jYByFW+1lhHRnwM
mnbKu2Jj5VwM5S5296m+6Tv/HnZCtxgvHV1QubJ2fPrUgU8coO0OrlQayxQyI3xi
bSp7NxgFaHUeo4zBN1PhAysTG+015UZhTIUV5cVNuLffUFcYknDMCvSTq88ycs/i
F2o44MRcKkQVVu3R6xPiXaxkkKZeelTDUOnZmFdSuDglFEEL971JO0T8HS3oTbHI
0oT2YbUjH6kgdYt443JVMrktsAE0EIZy2v5ltC/XJlqPQFxPDxkf1k0vzeg757G/
Y1+EA+DKA7zC3RObERLfVqzeaJy6RzRH8eGNSyI74JrXu/x2TNtFwyj+rFXIgKOo
nvJmiyzV81Ghewi6D1s31gAXeRyHlwon7X4DSxNJxDBkF9D1xkKjw0obvACdf1L2
YcN8ASPoDLTYw+0F55BZLv0VDvykkhVQ/p4ea63aWNXBdAaThkGtbMQ/J/E0WDdm
yJWGKB7Vm0yOFSnycuRRMnevPCShgoU29oQfD45CA6JemHNAg3ye+RfBkPL9RvW6
+CqSEaRX3YNos8YpP5ZODs7teqDJRUMcf+K0/ZsN8OKq37HsdAgLxLQEIgao9u4z
jPLYEdHiZ92RrnYHpZWuYKbdJix26iuU3GKw7K/RBiAgQaHeIFHhPcdcYgDCKkvH
aKXiePf40wl+jQPDYn+v1XWnxfNIWkhxNj6o8Sx+LkiTOYBJcXoxIeGoCmB6jgeo
+pID7IQWAHickBkd4X5bdfjaPIkdsEtEpeBLqIiRnWNije0b3DxAvMKDjJq5mBkr
f5elGht0/ya4jhE11G2AmDwHjDvWgp1rCN54BrXOlXpbB8GNzoACZcxvyxjA6Gle
/pm2kHfElCmdd1+hXJsjaLmKm/EJHtZfU0LT8XzaAL5gFh6jCQjShRcPLleyPTq2
ueMvrpxvCXpHL5oe4sJlttK1jFf8VHOERwCZsJ9MzTYaHXL8VxB8ws+wpl76YQ2M
fPtIlrsQ5hOVkT9V21R2Imgh3ATPXgRAD4gXa3SZl5JIM3Kv4jbv5gm7MLqNaKjp
PB+j6hvjuju+l/CppGpZSh7HPrbE2UNmcvAQMsag57WdF3zuaELWlDBYHbzC92b4
A+D0MPk7a5JXT/dHdY1h69MrTz/eYBQgxcq9CY24aUy6sKJlwsxNgZdAWBeOPUWz
hil9odTcwCUHrflRsgp5iY09ixkJVbK564yJtitKlDtU+9gDiu0aKoWlHKDpUGKL
titygC0qk8SUrdHTyjrl1GYcZM4YKHto9EUCqaD9VnwEcDoWIzRTeeZ78xcx7g+X
RManw1H6dkjPeJlQzvJZ3cdVMqk0tIMAyX3bXN5qbzo70eI56pDr2auPZ9cvbDTw
oWF/p5qUH/Fyr4bVtvzmIy58LKJEQc3XIYu20XPS7lcb1kKEIKT1UJNXhnZ1k+LK
N8NhJrTepl22DMpp+BlmL0w1TeuAfm/5GRNJvDckbRKEhSL6LOgNVm3Ro3jE9j6w
l8BsaOs3nTXxxilRidtCLEWrtzqnKkRU+JphG/EUxkII4jMxDKQrnXL0xMzURqoU
yi0jRjy7JZR9mwKth60yCRWxaPBpITY0KN20PvxwJTOA1ZrQF8CJ5hZSKQayXE1W
Q21pvv8wNY4ptZN4um7aID2DLkxmW/TcakwJ4ArQq/ep/6n/bVZrMSQ00by06Gu2
kSNOi1n9zbc3HFu3pFbizHDl+1CJQsfQUQvTECn1+H2n5uhb8LfzQM7azd7ApMXK
8w42ISAr7j+qzkVAeXHtraPhdJxpBjoJKL+Z44sZzUKk+bW3De9TGVdVMSCu88lU
lbnLSO8VA8xtT0DHRK1wGEuJ+KgH2RgWep9W8WSFtjhb5En6tmGod1z5KEQvL84J
Na6kqe0+j6yCyLmVEpOAQwv9BUp/0UxXjb3bcaM2WnurycRz6akmmNMP94N42LsI
OJ5lEcgFAmL/O5AXGteEbE7HeuEGg01AMT4BQdwx4xXmRssJ4Uyi4IZhUR1qp+V/
XitwD0ksLyrfYLD7IuOWgSmb+aJvn8AIwZI4cbWwnmPEUUQTYDAxeWG2a7dQCehb
BkPKD6Ggu+tH/bYQ963E29PU461gnHCy+WVqWMPalxAJkRz+/EiOdN4W/XJkKSfR
xsWc+oQmr/0jhPHct04X08VC3fel+sjTAROz/DbdDeBCDaDD4GFjFNjZAOCP1zcb
ujZkfJWFAWbHpPJ3QP0eHIljQphA5I59lsf0ft1DsqW9imPUkUXeWbQR25OFcRwA
i1pk9S580UqqrFj3An2jQ6kdY0oLzHLRlFShGi7CWyqhlDigCe/pSpwU52AkYWr5
CVpApXMH9J2AMxOrDBh8l8NE1Lq7esi/KlrF9tWNKuBxni+AaBjVRtRAFDa0fS0P
ySP67ah6UrHCHW/4XBq8eQKTsM3gre01qYSiSsLXgZDvN/uT5kzz4wlUbMC06BvI
9XVP68u9GLzE6DI8vrU8CmhcXkX5LRHM0J6GGt9gyulJC/HbCYIJ2jIduw1Ttm0i
98v7rduwycLhPGHKXS5/jYa3CLSjXIfEhMHYNXzm+rQQooWdZa6tYzh1F0sV2RDf
xsJvjCbOiWIEd/3MgcmrJ1hDkmOoaNNH38wyV2dBJ8QeWnwBwnkLhh82Rb+xBa4f
GKd00x+oTI5xaaIzdA9XZKhW3HabM1jDghafHdZDsV9ZaZ9nJnDDuJWCssPqpouj
7+w8x0gtdfaHlnhQUbyBJyS86a798jFL1UBPgGN1mD9SEiDa0FmAyiDz3kfHEvMb
sc5gI87AixnxKuZ40CfY2TB7Qb+H9L04fGIN7OM+b8SaqiAmPk/6t+6YV0f1d18e
BQkq0A6YX5bxCjo1wQ4b7GsKkWbarURBREYZdt9FCrPSfI7dZUGwiKiZt1t+j2MW
NolbPaap+H7MRa91SHiLhacYj51mwYbc0qDpk2a5FVjfQ3uvUsQL8FmHEUUTyCx5
+vhJHRMMFkekQRRKfg0Ad0gICS35fONN7UJCRP2lA8vx5f2ipCJuv0kx+BAVAoLR
Knxx9Q76W/7rMB5X4x6dagb8KmqODzXidMh/7LXnVweRIIVav7/0APSA4OnpRxqc
U4bHttSUG//feSQHtEeR54huVuCqYbmia1aEQpSW+QXCm8TNrDKlFmtY464rpFmj
Jz9MwflnqxbSKLTjzPdJM8/FeyiInNsdg82SP8tYYP+HfBdIC2ZplbWbul7Xurw6
leV+5O8txIStwYN6jcClvuZ1R+QIqJ6ZQklIfjUvJcB7gF6dReh3SAM/pCFFgXis
xcxVVPqdbBHfCt9Vw5d81doEDmMeKzidZl5r05gbbNkYc9BWji1kT6Esr0mwf7lE
6JmNArcsuNj7wDeNK70gh0mKJq3rcU2GIDd8Tw4k9VkyuTozaOvic9dH+Rc0OPVu
RgLkaZ903+AUaT5WCQwrkBuRLHwkPbRE0a525gE/R2SJw6PxTM2dn51Mxafz31kM
jUx/wzuF94FWSLabgIRYwIfiayTPhlJMjlFZrM40gI17plrQTE+PoJA4JmYFfBt2
nRiauqBvPVIu/cvBxmFTVdF5cWtH+eK8hnJdWzPUOL3ejdrBOOG01crJUdBgaN6n
z4nzgXtSBwNRf12BgZQ6l+jesOIF1wJnEVJSUI85MQfBcKmRDjwvhBLJA74mahvR
c6hAoYkgg94lffMAFfKqc152T+dLzLvLpFwovNnEgSsoVS4QSS9voUNCDAnLnuls
c/Nl/YavsEU9kgEi4irOVr8/oQZCGVJRDPJJWcx4fn7ZJ++HxZbnDEHUdPB6actS
z5bLpphETifuuUBX/JyxCmIp00Ofv5EPjGOvsSrn9VF1/svgWD0RT5oYrfeTzCRa
pMoicZy++qt4RCjkrNDvbN6+UZv+jbQGdSlxm58TdH6nih5ibIs2jVV8RzYFzKzT
1rASfg7sfj5Tvvl6MKO0FSK2XcqXhdUL4FiqwJ5EUO9O4Agu/Dv2Lhu0YFzdwdKX
WNXU1TbbRPotXfGRsXstS4JP13s6lk+sCtKiih0jAchiYVV6DFol/YM2JItVTnaC
b4V5HEvjduEIwNuNN21/7YE/bRuOhlnbSsuAS83LkeNGmoK0ZVei3GalWgbdMGVg
2i8O62jyvj1pmhZ1aIuYRH0ztpI3mNBLchsufX0wkY4M0VHPPdd8J8KFldjTQLMi
KrNSaSE9Yk7kWnrqwA54YomOP408V8Z5HkE7+VAZB/FwROfat1KhII1g0XP0hfid
zQauycTWyJjaDOQRFzZ+4cN70YepaP8K5anzSpBY4Wxvdxim9eBl1qtc/bBBsA/Z
CktY9CKSVD5wcE2v/WD+/Q5ifWXXu5SNsq8R5b2ADYu+UYZUIsXBQhllcFFnAXtn
1tMUVS5E2fgnmXkl8dyGrVJ+RQcPXtGincqp21cZQjm31t16TBL8R6omYk/zRkC9
z9c8OW+aCHIG7QSaloLYZbNYcKwQrOvc+WXsIH579928wEiBcdBZRlD1K18WnRRY
GVseaZhm7IYbMcZScfk7sSv7hrqCjXAsdP9iUG0ZX+m2p/B8/c/yC7G2Xmzg6n2O
zal/DsfldoDcinwm6FxOj74odpjaWoVPRsAu3tTVkGH+p+s14P+Dj8uYFVq6QaMy
a3cUkt0K3toNwCaTnyLbfer3dEBSm7Q8iTXhFPJBxeDBnwExQ6YqMUXvr7XBKyqD
qk4ooUBafuYpkHJysJ+7id2thuinVjF2BN0VsprNb2OsrZgTEBHDDPzgEj6kCAEd
1fv3iAlZ9Fo2MVebmLUhawEaQKW2Dsv2gLO/uRTzsEpkHiBptEMMAoVPr199W65e
8W1LqExq6mlAoFQfq2cdFa75S6zt7HypqNvlGSXrIc9ay6I+0CBkWqNm6uSpKFI0
GdQDdE8EhZw2rHhzMjLMLRZtECVw9u/O7Oiz3J1NFi2dplC0afCidNMHk7UV6upr
R7WLRh2Dp/ZweKMbf8bMWg/ZrBgKEc09VZPCB/07xbldItKUsi+LPIxzLNwP+Tqv
9Lz2KHCrVY3Kfc0nXUXsU84M4QcVZyvLUl/4cpvPLvXsoYOsKnlHn/8KZZn+ir34
S+VOMCi0ZS2WW8sVYq79YX/yoknKQ98/BHOcXxCAgUMlor8lJo7ZdGKq8CstGbqG
xBbrnB2xojW7rlAJE0idlay6l5OwW+1lTJtSxat1FBNmPEZRRt5f1H034tod5c0q
IYXy518I4GeFNLnrSlayI0GuvEJKyxq1qmuq5jtzInEiNrLBz2NNnMQlfMYtfET8
3GrCJulXf/8OiSyDzXF5VGc34YCLKWltz40OnnsqM52NAvotlKVcwzJE+ca77Mro
/ylCLXSCzuv+guCdfaN42uuRWIiukJ74HmrblfD++4KtEQrNYRdDtNzMT2cMoC2L
Kdl2N6VfpHE18RHwrp3WAuGMa28P27hYouA1afLyxQRUfUHrnfJ4OfGvXREyHnoA
J6OjjsoOCWGgN+X29nKh7WdtjMkGLRy4RphEiT393UeAVF1W5NoSUtipupzWs3gh
kxpXUz4Psysz/8dE7UJV9r3umhvq97Dgu1ffE/WrtI+egdoaifkGY0qBcU4Jj5On
pwPg+RZXVGFii1+3D3HOVPT7vjg2ko4sUst5mWepbMwUa5Wsjr1FvGj+isRPiulj
lkvpl775ROTYuV6ZvEImSd7ArOCNWGrquFb3rTPy9uVWXaq9cJEALo4gHVF5X3wG
uAOg2F59Pt7usdKJvcIbv+RvY/LbfDuxgbYVERLpn0VV5sOWIips3xuzq4qD0Xo8
aipJF8U0jsjXmxpSgIu5FN6y+lGA9+GK+ZIHX1x+mb9A6tROymEksEgz3s7jGD1y
bcpVPueQ1thJHV7+z2A2nWh38ytPTgjkZ6vQCldabU1X1+v2FhEQk3io7SBGNQOP
w1x1tniXjnPh6MCMCyvyHRnj5cWTjeS7FzjNbzVsOSSX6kjsB4OcEbIuWvsvRr23
I3sQCttyTRcLi5bMiZykSxxbQuCh+HD0AgiT1IyYjZTxKhlvmrOoy5eUJF1jhMun
pux3rkFfJyg8XfuRQTJAfO2yW7MCpC141qQVq2A4p3SiSS4W9DVA1cbmUGtYDJO7
24eJ1NmiNqqgkeQF6o7L6xX6H+7nApdP8O+w4cDJPaOegSpqP1DLj+m3OxVsmAeV
43ogfSaIkbDGdgaVfxFUGjE+omfm/7iPvGV39op533kERAYRikMi1KVx49ODbx02
+/lCqTozoOErVK6pw77fLlldnry/mf3CGTMUwa4wMAPuHAp2uE8PDZ9wQFF3ZHxO
Y5s5nicp9laDFmIviL5hkgLmlKnHnybHKwhu6q4SHeilF3AA2uLd2jXjDHfsVPY0
YV0zwaqdIeQx7kZst9yi4QRLnMjpphNb3yWHWhwtLJXT/hCW3P5Vb2PtkA+Mjh5L
3BYZMDQN6rtVoNVOgbDKcg8D97Zg8Scmvl0299EDxyMxmo2QvjPONyD43zF4YDJa
x6rNrPxT7025vwneAhw0vvvANS1bN3gy01sU6p6oK3iJlIinQ7l1IEczRrBUQeA/
IjT/56ehhlXRW4QTRdcnKf22+8UnPk6WHuIGWUVc8o2BYU9vTCAav3J61G3G7fyT
a1DM6lUl3Qm4tLHGgZNzoMB5qoVpwGIuB26pOrw99bVJzKkr1cor+kJEG5fNaB4A
oHGF7IazpjY9iHo5bCuDTuIlmwxj+maMTJRy8x1nr2QJtKRBb5PSFQdTVBFK03DM
aig3/+7q4kkvcDC45tC3lzwF8XlUQD3+w1f4mx7WAkWKZhd2VN7uFZO2+JFkQR7C
hsQdUAATd2z/d1xwTCygGiF51DTN2Ukm2QCixTC/xLla0g5R33ZYG1Q8ln8lImXL
rzwkdfvYNR611QfaNNzhwt/7BRnAFtRxeVw8nSwwryrE6r6rzS/cv1qqqqgYEmO8
0kZQ7OdHV4lh5W/1TjT9zBxAlYDKXeCrfORyOg5Bz7gJ/khlTkZpq8YDrgr3iGCp
KjS3ISpmZikfKU5eT4dRtq2WpuCV5TqBlu3iuR4FNJ88JBk9hp74UubZUU7X0o7i
5iW/GyLIkWXGvV61QAjDMVq8iCBoqoKxpAujun5ILQ3pmltbCrUL9sAMNyqaFOx5
fKzlgj3HOAmDu5Nt6cRpwso/8SYmHaUIUxf7dz5+g7PEQK0RPd/zfAUEt6MGNym/
biGP3AbuT5PaflD32G5Vlv6Nz6fLVpVVmdFjW4jl5OymO7F7V3muDaYyLEOcNXmo
X9C7rlS0GhBVxQoXNOg8i/ec0nvsqKzMF0MyL7kTmLLCKSesBloflG04hh8OlYw/
zx1H1YPsPuWkzx2mTO3jVXxRklWMuGqEXDrzLkt8gPq4NF4g5sBrTts1+fOLDGJp
Ejn8hSniGau8NYV0kffVcYfkrkyNHMBs3Vqzx/WvdX0khpbUxCj0qcPe2PYrW9hK
Oq5AtjfPWfOjaKKtuc4/QXRu3Br3N+XbBXgBwPzp/HtDFDAMoPDuNrvJbIWL+50+
k9KgmtdIJK2/jccVpCt8x1OOqiRIeaoKHjGVXQWohlvNPBIyQYZREJh4FLiujFyN
P3IFdkpXdJqnRjttnUAdfwh4A5SkNJBS5Q1O3jQEPkOlE6MioRXEWvDXSrYquJyd
w4gIbqyVTSkaXaiTHpFK2DOwrfuZjr8dg99Fsd7oVUOKXNtYnp+C24eFS4hsMpOg
H98mImk3T3AG+2z6AYw9iBiah7bohngMZ/BeT15rCdOVfFo3pfWMgJQ7pv2efNYv
CpXr5t4ohEbj4nuhCyYa7RHrUf8McbHkQjsNVTu6q3SgrJe8jydZLn/B2dVbMSnN
bCM5tzbu9BGc/XxtKQcp7O7ZYFlwtcPDyBHaK6z6/6hIcl5YWhC0qf3dd8F+RY6q
eXDCt4Txoe8Dvz5rywfmce3Z4f2CaKTKy6SWIdZA6POo/HerPLBlXO8LEiO7le3W
5c2LHB9TfHCFsSP2Ws2Wv4TB9y2sioFgTBocRzYG9JAG0IgOoCK2wJj4BkLkhU14
Ts/k00UyOuEnjKUtmvUl76/XxAMOramsiGQx12P37Cy+qy/BOsyBbm/RB6S/70K4
c7OiVsiA6Ux3V91AjgLRNh9liQyHpVgvMPU9Nf6jwCJSj4HLYN0cKOG8FgkpRBmE
c5F1IVRdpgUPGZG/KhwD5kKMh8pwrcZOivFuuDeIgmHbCAcRFCPcR1U+/7U6Kf9J
fxDmHK/tct2tHp1lc3RlCFTvXWieVZDtAia2CAVv8/Ce/CHZp82yK7n3Dw2WYfL2
QNXevQAh+EvfBryCYrTetuexDlVdO4RzU9BzEWbvdcqahgrWeh+Y+G64p77S7Ixm
RMvxKYkMmXvSxeInwsQsXe3OOJEDF75rdDAbIdPBcIUkYy0Om6WH/ARZcNjjYVAq
QZ9fXTt7LP2OhOHprzi+oO45MlYIlRsrpbJSvVLzVGj6JpDPyL4Ed3ZUj13hcBjZ
eu48LVgsk9nJH8qaIIjBetgFfOlYx+XV1370uaN3648IFsKGjyffoamNZgxnYFmi
HDyuF3zhj9Ze8BXq0sp78Cjb7cd5BkqXU8u6OT/NVyxRYFJsIxXyDiV2dxXO+5wQ
VTY8fXxMjpOG5HjTjob/LWG4BKZ/hiNqYjohhM6iZ5Q1vHL/ThaIf8vUbVfy+M/Q
EnXEKg91ZPucEBeYB18aU7evPiw6zXVM/ajGsFKUzEoOtS7JcRjIStyR/D1E/VjP
oJFnVys4hHxI7MQLDKS49Y3gn9P9xEiJnhgFtWS+WHU+BiYWfZZWTPCTVmzoUxLa
7RHnXr5vgVm14ZnI9SeeZKNU7fPDSuFiOB1v0cegfmNqZHGJVImu6Ievj8dpxWEv
gLIFWORc7rEVmGFxUhUM5Q2jJmoEgBUlu4d87hJR/h3iA4soYJRrpZJ5smS1HXBp
sevTTLjIrrIVKCsMuMSUitb9J+ytM4dhLNwgNiDrDLlbGSr9cVciIeJHxx/bjChH
+yI3y4imj1Le/zzSiZeZdVrkctWJLfDrBr+hBUL5dFzvqi5/G9FpR5wvCpMmiAr4
WFdR734nH2YtB0+gLQWjkEWRn592iCrvX7+D1qUiAzV+4Ow+GsMem7Jz9YASY8Xk
prby3M7OrdXItRsucWXlxsU23y/klNN4rVUbO/N1NbTr9CxiCgOByrpByiz/Wn1A
GswOel8iK5LDocsO6pTV7YAQwpSpBKW1izEo2eZGLQLYHTkBhx/WgpFGOdKZQB/N
mtcJatM/6CFDCBTysXs1mB9NwHvgzcLxbkroCQjgo0aJR0/VKj43NBFrSwi2PYhm
KNe2LT2khRHkqoaypSYeSjaLabxYgzXtKli30lrWvUaHf6ZuAXwV77tEukcBzSKn
a7zLQFl2Kkg5gEVdUNtBzMXekNKnc54oGYz2yjy32bhuFSXNidWTOyTnWWnwn9n3
rcrx7N1NMjB72V56asSUnDjD7acb2ASlWDYABACDlgP/5LZnpoqOm/+KePsTXP5a
/HYpb08e+7da27jSDQahse/sCGb0gwJ0NJfQYdvjVIYC6wYJqxBzd4YVQiaM3Z9B
hYhxMTwOCR8qGoSjyw5uTisPN/XSQZpwZkqdGddHvew7r5HL9nM2RKrbrWTOT84a
zKTQ2fpj3SlS6TM976aspt33PbfpI/Ij3wNsNHNWrGArhQ0U264g+DJiMmsWIr0Z
WaBdfizyz9U2mgVcE9EhxuCS6olTVw5cC7Z8SWEHeRz0A2UPuhs0eeoAP1PbjJyG
crzNIoW1qVtzQx/+8/hzTNghNGsAGOdG0KXjX5PDvhXwSCc8PycSt+Y5JkXehmFb
5eQBlX4lFpgNrnR6N8iAYAYuFLBPq4DFwLjfS5jwo5U3qopM9zLJkZ4yqvN+UYJV
12zCSSEwd13lfE4zKoXNPOQ0YR8KmD6Yl7la2i6XpSqF45fGjQMfm2+0a6TWTVrb
VdttvbPIJLAFOCoPpe3ZTvnHP9Ivg82dS9R4d4bZ/CHLwjwK+vYzMlOonuS9JyiU
ADkhMzAJnWLDuYsGaVmQzFtwJ7AIcnNX50TcjJxKS9qXwj06816VSFDXj5WMKq2q
jW7z20as3WTVsbNCz6uuHTGuZZNh+5wx0sgcmWEHPEBxSsxUrQy3uXGquJpfKtg1
GbQkFAp6q0jaoU+JbzHsmup70dpGaQig5KKkQtfnKPBxWFkOeedngdAo+p7fxhYi
n7YqVgn3AgjQ3/gagm0nWHI10NaQCsoSTObF35dgThNk4Pm9Pz+pcsz0SjDgx2QM
spRfnTOZiY7D71DuUz7rS04ck4aLOkDKxcel58o75i3ZB2ivCvi1wYRxP8SVxw3i
LSl2zz8W6KCjW7hxDvvceVGuLx7330zWYz1JDU7MKnCHFPSqIxNVUBQ3ZJBKPFLp
OX0lVeFd9J+kmqqaNK5ynB7ojeKwxKTX47AdNK48P/RbzJKIsM4UJuBylox1XlFJ
uGCyUzIlmzaEVTvtwwLc21ErqW6tBlk4FIVadELR8gBXGWBb9sLaWjxfV3RnMKzF
hL023pgODW+0+wsvDDBBEncbKVDhcU+xuFevUQZlpPErl82mMI/aILlYJhS+4st9
Z+HVZ6CNy8xWLIbRyr1B6jri0cYXiGWmEFkWCWpx9yRwgAEjAAQaw+nnNXpsrFYg
w7LeoCTSXcd2QD96WuNtAC3PVUgpON3lYvFeXYaxDjwfC1W4UNviTx5zLeSpfigq
BWulCTvfSRfRfRw6zslDbFjuOjG9kRffMaPUP2a37gpnFsRXV3qMDeXOUPz/mHLK
Dqlr3Hap9hmcSNh8nFbufNS6hfVmk8iiMuITOg/eLr2wZgJ7FtHe4/LZ6K2JGqzN
Z/XmXgo0sV9Veuimfr1sczHfbKu2L2rI5gb2L8M3TxJ/nit761w8q/XcUgl1d9Qo
ImdAVCms9yeG8SrM2tmgjeltB8Vw2Rz2+zeIQoIbXZXWBkzVTHkeuJwarOBpOz57
c7xQ3BzgwiaBXVsraY+rFvm+uYycgVGdgANLOtiadpVfnzmMXYVl0bCincyH5zZ/
teKYNnApQX4PmTUdMHFxkBDHOxvvkWFYqFrPBMI16TiDVvERLOc8BfNTtneZbUeM
bO8ZYIo4rslnNZkkgr60V1irHLeJ2B1in1olvMlqHM59j1KRHjb8BrnGqeTZPwnt
lrkdjNzBK5OLv3SbCqqprNofXjYVh+UQj6Rxz5eXsOuv1uhwIy5iIPSqKKb5mbr9
CHoC+W6O/vAo9szDRs875FdT9Y+36EEMTv7/y+yYOdmRDS0QppZ/jg/iGAieDZup
u6fKtNdsWVQITaHstbZN7e+FJsMq1TKhq3xIUQ9ziV6jACS86M+e4K5oHmajWBBI
d4RfIpu9A6+BGr/auAsBXQSEztrrQJrbjKC1qSlih5vY8s0FPWiKNqDVuqpoYq5W
qQTMCKeRI8xAdQEfATen735c5fQurF8hsyHGQ1jq2HBb3r6f25A2ah6NhrZRIJeV
T/NYuCwSkVmLySWOJeumq2XqctGJowMtUHgI4A3FnRNFMS4QWWHFKx+jVCYHGvPg
d8CINGpBmtsQGiu6Cd9R0Z5PEkMogg8eK/fBAeUGWqsSISjJ4G7ZZS0NBRHm/LVl
x8w/mZyHZcpjhc0OW5liRCeJnLPfpM8N5iR3RoUvp4STwLicF+1A14aTSR6VZHB8
TRSdPCdbElEZmkLWEdzwTZTUWRL0gfKLPzXu6OzVn1IXpt1/kW0Ua83yQGmD5Abu
SOrAdLshy6GVKBWkoRVPgW4nOfUEv8jwibIafUQNznDo0hzRAj1z5K8HcLBtGIaG
cAlaICwv1Ctq0DsWq7LHon2P7w30k/WAIsQxUaoHugMtldNPZ/SK8AKmg0x6yQd3
zmLbQxdUyMt+aTvL2Ld4FYTFR8nSaGnaK02hSYqK0bG/Pd3/0gbTuVrx5/wb14Ux
lbSeW4HEgRVl/T9og8xE0qGxnPBlvTV5HrOcg0F/tEtfKzkCes0gj7wLbvAIn2ur
4wYFZPGJRYwqcRaHswf9Ji6V82MbnA7EbXGZstCTBBZTnOkfqNmns5kezFaojfYK
dN7HN67uNX2ibOC6luD3p8AujOdi/AyBV4lzzMEIr7iNjeggPq5rci63rinl4onK
TUoREKuo50BJMS1x7b5yO+GCuPDPMdxu2pe5pApTB8b7epnHpeRLYBGIrKtUMLA2
u+vs/yI1X+l/ZxOYMKTYStHbTPhYaomviXH4IunL7YAuzrHEzufYCtErQY9s+0UQ
UK3kUvNY/NMY/L/IHZZomMEYdRtSecyftXRRmvEvn830LQ3YeS6SlmEwoOIi1jjy
In1jtElWpPfhwoNpc2vrlu5DPY6sd8b2OwWK6cULha5b6A5T9nFKJkfMKaksWUV+
pQEg83a2+gZKqfukwu+z+pjZQc57L1mfac0XgmXWXWyTw1pvKQ3cRP4hvELcG5O2
UobOtBQe89CapUmpbSm4UgEeA5MV7XIfABJRfNLolkm6TW9UVZON0H+MoTy6VS9o
yjqz1utGS2JyuMUXwdjInOU/IGTownmncP3GnvMtvg8mAKos4KQO1BRAA4Kz5NaN
6fWXF32yP3kASOp4WpiBg4Qj9uRZTYErwPS9lKmXUadI97Q44JqDCI2XlTp/zmqW
mj93ghTYRhyZKil6PuhlkwVtYDnCWit8JXm2CQT3wbZpqKcZLNr8ikCeD2QKyp0p
pP0J5QokUX+GvS6Q5J6VaZ1PbxGiBhnE4J4aTySkVVEdHrcwS3h88NP890KmlUI2
Zbz/LwKw/Jnrzk6/vn50MNITatTqJ8fAmGPhaXgMjkrce4lqV3XVSOf56bvVuWKN
CGowmBvQAOR23wi4DqPwMWUs+Eb/cGFIIoQzGfd28+rbiqFYwLM84CGK1KI7V/ti
1YWaAThhaEX7UCK+qvcFB7xSgZZ8+riIMqo6hMnot5nnVRsqa+VlpMj/Dsyw/5ei
XOP/rujwdmx25mfYznrpgzqjdCL9MdmoN8UoC63Bix1eS3I0lq30FBuSGbFzDbiS
ygeHcE5iKEiXDWhqzUvX6Oy0B2COws3GVz278J4f76+QKpgiKmOJRXeUrX6xhkuD
aKOrNaFsZYVcqZXi7xbxFYygZPMZsWRhjTSjBR1k0H8S8LiIxNZcXi4crr6/GRzM
HTVRsC10SRgxwKYl+thRvVl9FIgVo6pz+U1/gr9vhvu+NqxOW0QVH0mx/2nGwBKL
KmfpjrLuFmxwW4Vgza9bIuMWzCusq5yMPzgjD63hXL4zLa63geM+Pi1gN/wHe9En
vA0PcJzy7hH85V2L3HfMbDkGFaCxENcCbyWZjJnVuS+TNJ1H1i4kc6fpoOWpZ6Wc
P7fm6TRvId4Mey58WYbAlJ8yQHac/+fAjsPNF8oRR+uRjHWAEXQ3rQ6WR1eG+n8u
ZsQP/a1t0SOZffFgd/ArTC+48Bj9IM2H6CC7WmI0A64Uy49mHXI7ayrBQipL61IC
QFKFkNCv/mQWpA+4q26i6hDrsWxPS+700k5xZJglmn1do9jaLk9/rwFxzCHHDvVj
Sh/oZyjq9jbdYHvsDGtIcUUsZNINKPq2ZWgNA21dOFIrW0Kthm3BWolsegqZ2f1+
cGN+ln+F6i9YQkSCZQ8wE+04zVgCEt0d8pARaKanZJwTycVi3tZV3pfQyCDQpSJy
XE5Gfc2KuNU+MWufDjlS826mUW/9kSYjnEjLp3Rf/4StNoT7g3a/2ZQLA3DrpYZc
/ntrhomyMyR9O2NWO8SbFp/fDtM6P3G7Tuu+wKyKLv7HZNKt2WOumTo7OPJux1EO
gqRg/cInAuAz0WINf9hbvIHO5LNpqniVA6M8b4pH9XcMS7HziZbyDPbwqcU0Ly66
IRZVoeTPg2029rOd2UNyFHlR3KUcWy71qrQ9HTONVsnCH3JtsmxMJdHJlBOlBEC3
QJ6nedFqAVcCx3XLgjzlNcUmg1rkCb2kv1oRGp511M7iIvvOe2JOB/qNcW0X6bw5
dtvb63WESi3OUjzSmBF2eD5aIVrDXrlDjrHZSL64XNeCJb84Cbyp9w0tXiUDpRLW
+Dmu6lRJUm2+12Qh68mXWYTpgmfuQuaTQHd9QjHI5J+oYB6A2JNSHOiaCPMQo6cU
GbGvlNyo0PKkjkJhw64cDfWYq5X5Gys+LOA9ASvHJP3FXphf+lkZu0cnqZtnDkD2
Jjkromq4TfVMhWNPYvTzoGQZ2pM7UOQCcTPR2Vk4FS57WVSR6DZ8NIbEh7E5XU5X
pME9wQNAmBDivGl5sfE5+TWI6A2dM6EB8vJZZ6n15MxBBTGta2z02VDJm1zv61QI
Jhl51Lrkcb1QeXAxfGlDkTGxXM98SEdtu7XGM/EXm+GFSh82iGCZ/BkJIT7WiNfk
qVLJRkzc0atXsmVLilgKWpZvLYrsgcuxi9y+NkB1hvxWFb5/K0Enf0GtYMVR8kXm
Uptv8MWrC+2IaEV6gdT+TAlaRmi6+/FDVxhT4o69c046AVJmQrCn+oxCv79rbZcb
uoJlHwY9YiFENu4qV1+mht8R/R3d/w7UylWeq1Zt34CS1IpZDFmiPoSN3jR4CrLs
rE4K4JTmgtHud2Qf+3vM0FEjHvbwJNST2J3/4tU2qETp+X2XF5Dpq6RRSECWf0YE
fZbG/jIRIIzwLpiTjbS/qlKJ/QjxjZFJENTSUQCVvXrjrjNR7ebtwfRt/D9Wb3RM
XMe/FHXfefEP1GF31VBp+JxYNLvFHtDkbopaTc9xGBqTh+EzRS/vBF7SZxGyfYTU
sLzlDGFbq3uT46PG6DfsPd7C2CMs4M65Tp3w6oKzRGZwWIKGW2RrRw33FFUD//uX
9ygofjTpLPZUQtC1iMDm94EeT8N8TdUeNL4PqeWAkCztY6+TVacR5VWh8+OjMjR2
sO4CygEHYl/1h7Pq8x3+RVrq2dARI5bn0RiuwEWIbty4TCkh6ue+cXSdp9SUaOYO
XcGmR2k+vy1TzmCoCXLlS3Oth339iIkpfhcwZi2sgn0JKbj3+JLcgJbey2KDt1ui
j/BcWI4+sKItJ3Ak88XTOdGDKZr/bW5n+l7LT/2bWnX+nYA3w8jFsbQH2PgNykGQ
ssU8axS1EkmTY7D6+4A8OT+XMJRY7pAnZUJ2bNz91Vd0vPbl0Tj/VmVwwElHZguB
KReoZIHBfkHN8dwonZzNOGn4lpA4f4XPpjeVg4CCshxQS6AhM1+7tABW025VEaJd
jVRPUnVlmkyR+3/5okdQy3PUvBofjHB3Mm76cIzpkanjQVvEH515SGsY/otW/uFD
XyguJP/BmuilEdakAlP5WBPyIz6XwkzxGG8rvghjG125gv6PePvtOL1ANQLvdLNc
4IWz08EpNQZRbIhv9sUs/atkhJY4vNacCDUyyJQisv6+4Li5u18z/E5zqfLAiLU+
rlteDrDZNGir5cdl7yT8OiZX7pebnto6q/K/AKXHjOytknc6SMvfEFYjI+2yqxS/
dE90EljTMA4hIc/opJWiMzRVFp00WBrWjPrFmCSAZb2G8cToQtzwsTOr3UXpFIFg
6GBc5v+SLX4FcsLb32dzH3y/tKKFS21U4y97OQN0jw/Zg52wKm9pQBDDfMOEz/WA
sH2UlC85RodV7/YxGZpqzZHaEURWUe7sWLJ5LKSCIEnwgL6zZbhsYTidWkjnK6Mn
DQV00GSQ0CBQ8g58jMdr23XPd6gYZLb/AIE5TL3bn22S2MhULtDwQfZedDPbWass
JcCYYPdVasUJytMhm2AtFHwGKmMVPS83fi8lcTQdz+C9F1ozojGiMR8ZfZVmWY3K
wbqEwwskr004LsZQlSCUUaH5zO8Ih7YxyZJfV06r7Flpwuji7kOUldg4ovKYJve+
FQcVdcqOmw33zc3D/Y5jsr3R7kapr/B9Bo0/cIIY962EM/YeT2VE9SvenTF+BVnJ
SeB6rLgj5w+aTWyCV64uhFu7JB6gQ1CDG3r4aHvwy4w1x/0fDnky8z/rLkIi43Gc
Vi1vf0PANh55YhXXJWyxde4D5mvrv7VMpr0mEm6m7pP8ykCHpiiBv+4sLYIjGFYm
mKFMv3SDrUc+geqh08E/h18DEXUbwy7BX3FFYwzcSlhz3XsFkAuYAhcZgTdPb21Q
SXpxn1z6BcI7Z0Nlj/zfIVcY8+DZrNOo+Y7jvSlxIt3ZKKDrkdCNGnRGRTgHr8+i
gNWmdOdCzYjc73fU06YtuQKkua+xFwbjYXquWIn0pWzMfetdidnE5nvEBg1va7dz
07Ga+wf94Hoh35a8PLr5Qmh2JHm+oX+6fIH3EZXPxL6pCY6X70FPHFi7Exjp9ILP
VsURjwzRLi/K55LTApRsUqUL3K9Ia47oIcUHGX1eNW2GzuTphXzxLZYCRd6NSg8A
BY3IgvzwY46qWG6X4ofdC122pDByP0GsxiYe10LWzfPB29U7VngYV4e4cG52Oe6b
TyfG+RAM55hoQJS38y8kHWaPX9QL2Gy6g4+X4j0wh4PHMx5XQFt4li0X9ZSC5LSR
eXAmIO+ILlVNKK8OaQKUCzLDGZLhAy/XK4FMBg0ENUo+fr0mT/ZLIOitJO2LA2Mh
TVd+l76CfInPiXaxMia5IdaXn/CFgnZCNOavASW68aTOV5MQPL6oEv+zCE0jHiNS
TF7MJZ/mqfqiKHGYx45tTrtYq5KXbcuz+RKAlJiCLgHDbCMjM3HzIH8SvHjFXxvo
jMcn4zjLexz9VPTcF7hpgvlKSKqPeA1ixgH6pcHJ/mjC5Y+uxx4HJLI2RCaxnGlQ
gaJ/X552J5ejLB9K4ETsBGAqINEwEmffJLjaAw3MggWlVRnUqkeOfb7x3p3op7N8
1oIOXAP76q3zut82b077VsqqkGX8Ecwb13HFH0Ede1NoiSNGbzuQKYTDz0aDwK84
s7JCgQJHtyMLMO/IIjJjtctMi5cS6qDQYGpzZgEOcSEZGWf/SfScQVzuWjGTIpRe
1sKKlaz0mPTKttn3esS0nwDpmTRMttR6DCXlrQRYHnzSn1jIDhboxhsNC1zWZwVK
3sYHsI9E6snwKhKKEJfYBBCYEsjm8wav450DvId6nlA+Vso0HbNC6MQy3FgLxkgV
UAGeGvOyV8ZSPVacfz2HAyctxh/2xJqXHZDj3h70fUMIs3A/vQsbYBtDrxAHCzUm
7NoYebt7fmMNBr3xZJkZZt5AzlZZfqHClFv+Kamqm3jue/JvRuZyyg6PaKeyfKSz
8MCVqOWALOLhTE9EyZMfAjZUxfeokSoeaGcrPYeP8M3057LLHadnnlbwSnOsleGT
RUmrhLKZfpgqFoLMc7PXLnOr9m8hajK3c4ywilSix2qXkpHQu4ocD5LGv3Ao7AV6
j4QGvp9B8he6mHlW0zNCI5gbEZ5QYWlAYQ6jSBY1YEF6FP9RsrsJd1cqFCg2Ix4E
3J6MDiIIYESVsKfv40kS4T0wMsVQpmDhPHKIWt1v4TL3tS/zM9F/WT2GNODnVWwn
EKCgBsvOB9w11yAaqHGJzFZg9I9C17ZxcV/hkyhl9rcD1ypMWPix0G3DFbbWAfFt
VE/K8bFVoDrUR89trmiemcD1oHXBaPDGv1kMabBY2Ovswl9vAlbb1RMN1zo0oSWG
wLHY1pJ5tPIMoGIRMrmxBxB5e+6YtAvVXgjA2w5cknYW7ecBH8ZAlHE+9IP3cpf/
cAtybapsX9yPVN7+wHx8+fASw229hqPK7ilMPCMCKqF0KGuD+sEs/juACF6De+xW
bDw1Ynn3sHaHZwZkouj30Xpid71Bdf2/a0Xk9tsWSobp9f4zDfEUx7ZglN7lkiS4
v4GV6tWv4Tj3Zdgt2vxYoAHE4oZJGbbRScqdFW0dFqn0hQBIHOfry1/XPPCHHyR9
1UXBvTY7uRP939p9TQqJxEi1/rFrA6ZqkEhLtRAPbJYleIJMpyp1dhUEXnUMiKQX
hVFx/44IeDfmqwUc3n4PVhtzFZatG0G5Ux5FU9IFS/G62g/8DHqqI7MPUBbrNBIc
TiABCSvSw6+OlOlmKiHEcWVkqtOpSwlwceMTAJqxeM/R10p7tfZZpr7yp6/BGArs
x6gbKa8RCBQTwd1FYGSWYvJ87slJrZLUiYi05DrsqvkipPvG441IuwlAf4IDqkon
C9vsI/p6g22BN5CvaK/JfAqHzi2SPfTaF5HwALf6go386zwv432RBt4v7QVUHpo6
At5p23iuUs6YuwhMdqoXYp+qxbbGUwHwscy2Tet0jb3ThpDOtjW0eDWi4eOe8u3X
gAlYg9rTkXRpyIo6PeEYT8lgWq7LyrmTncm3qHVUIXOdgBh74koXHYyPthejA+Sr
wjXPOqwUcY09eMopXefM9PKiKElctNXL3dUy04Ww/gcrZtRruFPETYxYX5moVfSe
w90TaEkWr243PpnJL46UnrNhUvIipntYR+Cj+C+Wjx1q0MgWnroeAfob/qM0QsVQ
MNP68JqnKvzbjJl9GQl3mFzbQB/+dGYQ1DSaH4O++yBZETQm+r03CsWhj+cm2HoW
U0WUemuicLU+pj+X1zFmSUZjmWX/znTS9nHOleaN/ZM/o/vJ6mSvOiTBQjbPNRHw
oJNLgdB/jr+TMxKekf3fvT2xwtqx9WRo+jcgIe9YlL1k7EXzKc+wTRoPKQdv+ORW
hqXqxHVwbGBloCH01BuAcve4NPNPJv+Jw4pA+/MgphjNyh1a/dc0p/TLCpqhJQQJ
BQS5L1p3iS93sw4ncBf84ff5FEd2HEDUJwdgEYqocvpTK91GmUTIZWkrk8OfFQdt
A+FE1AZ7nz58xQEbwoNEoBCxOjIxlr6mvYffCyxFpKfFh5CgUageEHP//eQXG5ke
NSgmZCxbRVn9cr6WKOnVfiSpqhQ/KM1cO2EGlljUoZhyr/FDkMOdo8uroTycI8Y4
GRBL763DN9W9ERji78bSk38i+HiA/6YSMevAzAAdomeBgEplYcWw+V4l9ARmRMcN
ckEpCGvC4P8/+zYxbu79COyoxex9MW6VLu17tNMVA7WD7nF/o2zRDsf/esGOHftP
5Bho89FV1bRHPAQn87/HalxKl1ZmLnyfs10svJpo/sbPDo72wlqEvHp6epGe33nT
dTaNrmErcrY8/4uqRWYfg3zjLxFwaOVpYY2xtmUXSToEUPXCPwc/LrSLnBAYteJo
tlPaiAaBaa7rxwImtGzABG6s8XSwziwyezf3Iafvs7rVUVq5cIKJRx9vbJvT6kPC
jb5S/8aT3uuA/DgOLbHaSRQrlOfoGhX9kMF76wfqNtHqVmFK2R8IrKwkw+nw5CyH
z0hExGp4+QleuJj27Y7MN9x55dfTc6c+PnNz61EocppqdRt51HxXuHY4TZsE0cd7
DDki9DChQ0G2UxhxNxsJxgCASNuJP+TA2p8sLlELuEB6nbfjJaX3Fswg2h2ugqEB
Z+BIYEP1E9VttFkvYbTMzrWb28XUjVjDfzB4S+Twc7xFQ+2GCBcAhXrhrQ2Zy1l1
/grDg3DpEE9YIv55YeFsACWR+VWfyZ4cIdiafxZVpmwXwcHhNH/yzQs4WTJyi2uN
ROdhlHkifJKkZ1laRDGz+dySnvdm1iDygGm2ECSBcahFunUmjfuVfho9lRau8feL
Mz0wAPotgYmlB26tERcaGLo4UGccjobbgLnJTd8bZV2cMU8ASVMEjTxFHcAyg0hp
gJV/sNifzZBnBRFe31d1nqLWhD9F5G7D3VxPlbDgWq5YKCRQ+koZpceDQamEFbID
TXDoQPn2fbQlizWRYbLneCL9rJwkVFOKqQqfg7dcxj/9hK8A82QL6mGBv5uwJmMD
Y9MoZM8b7LthiZZDCafYkJSIWvzO7K2cR4SFbLU88Vp0aCuGpAUX2af3ByqIdkLP
y2+DeI1xTWIFsVWKMnV2jkRRACTPoPka/RAayW+MPfJsv6e/2t2psl918g8ko+NH
QlCZnbmdPRIXFjHhv8vUUpcIcaCYrgq7xNnjELo9KTiJa0Qy/Cjj1q793b1FkA6T
3eWjxhQpjxUTi5xhIXg3ZSn8tv+rocyagQNkUN+kh83kzOOrdYTLS6FY7JTJf+3C
Q3qgD/hByFhTZOVJzZQV10Lno10hLY40ed+gveWy/g4uDB24SI3F2AgtX+GTpgxm
dJfvSNrmdQeTgwIQL1j+8oU39GT55wJVux7i9ht1h2yNx2KJAcWE+0b8UtQq0q+x
ci8ruNcjasN1DpLxNVPgYStC6dux7mWRZYr4GtTkSiCs9WFzlsuYhe+4OQRnF3Kf
XfiIQ5BgSrNdVz06ldSBjpSIXKFKWZOuSee8Yi/tG6t3lask7+v1pMtr/TWmAJdk
/0+Uo45PkGKPUcS+vzZFlDxlU6M9+a0yypaoYE+/E0PoDQRcTyDKpppTez7S/yDi
A21bpQWF0DFmCfblvSdwf0tdMX1QJtZY03TI2LZK/TKvETCmP0da4yJtsvCF55A+
zCesiJW+to3sNXF/+0Ebal0HYNDirpWZNShLohHBYIvmgSRoHW39Qr5baSPLo1As
D2Kz2k72k4fOPAJMMdsSvjcryQTDaqYwQhmRGQTI0/fqOZCOOoWyE+uHStnapTkw
FXYA25lHmgyeVM2O8gCDUlcTTa5rsnp3A4VgujZchBxCJWMaTV2A2u90UuqHh7Yb
UUBiq/8NTv43LnBCNDZ+o76AeEOGTEg4QScPByGRjGbqQW5IqTCL5j639uF0a+e2
rJfiwrW+m+spf6gNApQHhB58Diz01ieBiKOEVaTsomGN5DeZs1m+R4CEtVxZiQ6h
uGurcamkXcnGKaiKIC9eSHuMyl5UzbJYcY8rg+JA+KMQheMEpLXlT/R5YrEV+xnK
DJ3oGI5nQRDmqnWd55c3OXx12ma61A+rH6vV0Os1ROHpo9xyyXpP3YBcZ1K/jGzO
8KJlZnd/Rxz7/O6Ri+DMhgNgyfTjL6uPCc8Fdmx/ISkuTANgyLMkLlDJFf7QwmyZ
nc/i/raefewJeGQu9XdOG4VRCh9AeFg3I+xyxEKiYjpu4v4zCrghGiv9YRWhP1qL
RARO0vqMOmDYEPGyLpuUSISuCj+dzW8N37DfI+RU4Ylqp71RYR0R2GbSwOpf6u2G
g5/aecvlfhrUXhC3RzI0wOuewuwIThOFH1lBjr6EXm4eaQJouQXO1yKbrFTpPvdV
RczuqEMCVq8YStaLh4Yatqsy5p9AwYiD3MF0+ussk29d4mwQ8UfNxYkFJs3AwkkY
3EEC5l6SJZWQKl8y5ZYsbjvjBVfOkw3fQ1pa5l/saEBUYFiUzREY4U12wI3HGqI+
Qf0STx6ZEQjAZhr6T+u0dYPfZiDeINMdJA6YvPj0DnKvpmpd1tve1rbkl5VYu8nk
qIBtznMgDC+UbHWDul8aoZlPo88hN8F49FpTrE/JnOIB11F5Sxy5J2zDAyMGt1gf
mGv+xi12abADNwshjA/UFEW80YJuOnlZLkFwHmreckLWqZ4g1kv/tVKHtcyHu3IZ
bxIFx/BAC4kTzhjq5EYeu5dimkeDNNUeSv1+bKVpp4euUK48RTmZZj0Irn5qCKfE
l5QDR7eRXIZjaFLhv9C6HlC5fPhnCwA/iERlcaPDoyvBrzy+ia82hqUNoHk7Pab+
KmI35nb3Wh3pwaKosApQqVrnqt/UoH7ES+dseqXtzelDuP9OqXQ4Yfxqn+GyeBdZ
sS0JdJam/VZqj/HuK44KCvSuAk+zVQ58dafu1Za2S2rE5YOxaDvgfYb+ofdRz+iP
/0WLEmaAD3dnPWi1Fs2Idd13rTXQllBuSFv1XVy5QXNLv4RBsfPW1SOFRpdvEgJb
/zV2qvLz32tZea16CXH5CyInhqVjo1GoUb7RfFpq38D+fsolFU0oWWT4gGtgK5lc
TdPXLrsU+WIrEnM545LoaEoOQrWzgDsI3tEP8Hc1Kmqahf+TN7RsNKqLY4IvQfEY
TDugWzkzEdu8tadnS56kSvo+mZy9wxKufKx+wlPC3KFw2N5MHp86YmbMKVBTZkEu
SsQ9ezUp5xVJu7uqrMKDCk6vnZYSP3f6f3DjAicP3Oyt5pusF8kPjkRhu4t2Yllv
YbV/clChIyW/zpe9batM3AY0v/Jrcu6/TkdhQc7U2zMXD9YJbZRX9NpD01+ARHOl
d04auPkqgH16P9TlPH52DNCuMn/wTO2YtSPIs0oDE3CZNUQrtvAtwrHcYu0KZ+yC
egM5GQ1lmOujkvxB2dQbW5hT34YZ0O/4FkhUEwRYmOywLC6aVZrVwZlAkEYkdPO8
FJMkunmH4M2YlRiBxohtlFF6p6SGSVWHtdaRAKQOFmRbCn1mWAdGaOUpHlKubPIL
Ms+degQ5cwS/bvB3L+mr1hh7mBN4yO9GkYTpd9CKjaKp/2ly/VFyakwfoJAFllu/
W+ykzV/W2VmwVlbMsjKy4yg05XcoTZob8xLs90dhf9gt1rGfeEjH/YJ2GdPQ4nrO
4lFQA+p1ELYrA0vAQEpdblpht8EAZj7KqRkoNTsoRsqVzJ2xrGvQbvXTUVtb7RwK
SMaAzW8IaH0gzIpKma/Dm9n/F2R0rUxYmqGh0j9gKmCMMTLrsIR1EXUpQGb7FCg0
F9WbWDplT1yqych+xUAO5Hpa7Lb32R02yWTucMTwHEqSBDkWA4QkttHne/yhpHSj
+cl7fLPxl64JPYjBkeSPbE8ps+TpyJQt7RbJCSCdAt8f6AExCvswMKoLGvYzEm/u
IeVkey2l+iVBZgEx6vjmwCCED9HAv9Abwnag0VDXCBUTFuy0rFjem4VCUATvlVom
9ulT8eHyn7HAN/CY01k8L4eFw0aELfEQ4PWwyACMyiKQv7IyICwZu3wbEKssccI9
OVZCdIyHnrfDSM+qsx5mpFwgZFFy+VpbwFIyBUSOkfcH1WiEQpuVZob79QwjCUJP
ZecQY+s7JgJBuir3RpI9OW94zrdKUgQwh4R3WRMSdDgP9FwuwrflOBFGN4PL66dI
oSKiunsFIUhDvUKCDbBOMaGCfN/Bk6j+oruLzYa6CL2B/PAPw3LirppGcsRL+DPx
qV+QzxmW2S9j04cG1Tvrz1oCUCrL6M/Nb7AC3M+mN4V/mYam9wO+H3eDbhr4UMq/
M5QxYiUHkh2KZjfK9je4PpZwyvThEoulxB7P+mmOcSOleEx+pWh7wJa2l6RBhq5H
zk2Def+9d3F73QTHwkKP/0kPWDbcXOipb50ADlY1/0B+Yc5m5HrsASjcWdgqKPdV
6Laylt/mLycu9ADbqs4Vlf7BWQz47DdGY0gw8NmSW0IM0RgwaWCcyh00HG27mcVU
vNI3OjLGhE3djXZLgld0UWcAjGw5bXI2IyKhrcsWbMQu4m5KBhaXef1Bl5BrWSAO
AMeiz37XQmLc5Se25hCDf4dPyBhDBrU76kh20tLxpa7L0LwfaEIwo5H6WHSZkf00
9ZJEZhBp4pfuaubIvLUGMkPF+ATbgLE2DrEbysbZ5m5HHnRZjvNZO3/wu+63CjIv
k8rK2RflvrswRZDptg5uORCKmCm88p5epvEmop/BHmmMbrkdre97OsdPsMZfZHcF
jGYpqgYfbkX5myhElqxBAgG3FQbGoIIKpbMVBDpyjxTOpOdX0gMZ6nc6KjnQkyPa
ioDk+xBIQTnqrS+0l9ZxQ3gC3GFjIqKXRFD23I+UhurUKRdS1a/XqL/fGQkpdK6P
uI5CBo7r1Q2p98wYtkFVcl5NobstDqx9yQjDUa7rgRYbPMYEwbsQbpig3ClEQByE
i/UrN+pP+5EiH1gsk/AQvT1a0HYmmUgzTXQBR+86YzAczKP7ZT1GBz1moGVrlXbI
79DUfqDzMjuSK4MNLhp+naooTfMAQqPxnHJP5ouJGclqNMfAvnxJozw2gDWxG/FN
sjESERwvLE748bXaMHU/fHVtM4nyzLerKdXglz8hvTKUz8q8g8PrqiObQDbvk9aY
kHulryqqUZ95uTMTQZrxOkzKENUbPkSc807F+/nBBjsUStWrwQBeg5AgJzKDxGFG
G2VnDM6AmNIt+x+ikweI8Z3gYMtsHK4HBe8P+wAzcrs0rB0/o5IRmUYqn2TJQ/jB
HEBYagENIPqMppFU6hJ52sN9V2RBI0hubf7aU4SeZbB9HM2lufBnckU/9+CbNIQC
DjEeBNgwPwLuPVhSnkpgK8RdFe/PMRyiLUYnNP5pJT/3NaxO5HjufAfrJOWx0DNm
HkrV0kaAfQIWjuqh72VMnbTnTKEHC8ZGk+sjCGPcPC4AtPfQNEVxqbhUlRXog3/3
SZYqffm1AzzKr3z1y7yvmccNbO1J88gnO/CjqBSlYI/PJ26pgGIrVms5yFOMwzHm
VXjOhxDvbp1V9W1B/z6iDAttozPrPZJt75UOCk+7fdKkLsHrkUc5O7lxBH/+d7HF
k3aM/L3Gg084AKsWhyV74oRQ7My7CHIlSQ3H89luS+SYRU5XGtXpecOatDha4TyG
IB9W9EKSNfGHpyyvtOc0F1cBFrolJkzSMbHHBzBoXKn++IX5xFNhDnuer7YbMbF8
xhbMJh4QfZCnrj4LO8LiYtdcz6TrdZ1B84HOl4PQNEGWC6Mv9YZFw4bx4b4kn0YS
ixHfL2KSVOG6vu2z8I4Sp4VZyVV9hDqgl3h8ik01h+4KSL5wM8gSaZImOdy2IqC6
yH2tbYPig8IUzhUo+iAjtALehYYf9faZh8A1X1zJ0pv5Or06aob8VWOFgIMCoRHb
/8+s38XVDlXGMSuy9P/Xis2Gp0oMKCIlQCqRdJ/9MwzbZGkA/TyDMmyxRj4iMsXT
pXJ9Yakw1yW16hs1qZwkcyG2tMehRcJSJAjjf0eDZXU3168lhyiVGTYMUrcJCY88
rGDhBGHTCOgOmOCsQEsYLKoA2nH9s5q4WLbdNu6Qi2NKg17ZwbBfxRo5bxSRjH5M
bq6h8DZFgTbh2r4PrWt2oXFS6kybfpXqc4df+MNFc/TgjU7l0Gmivc4oaIn40kVK
izeWQaLrZUkrJ6Tru/2MaUQE7Q6zTWY0g6EOQY1jnGpBNwHySb7IaifYz9jNT5pf
kBt+2UtP+Sr1bpUgoJKSqio/OZYstRypwQ2KQ0GDqRI9v6DwBvB1P5M4Bw9YurrT
Iyyqnc4A14ugJDhInMn22pk6LKOkDD3jg6tcew5Si0IqRuZruLQ3i3M6mK7HdI8A
53KVVUv747RCnqnRoIUui/IID0iOG0h81fZsvN75UahsM/9lgBHnYJ9g5sp02BIU
QBgSH/HddMavhK236NQTSHEbd4EmZ6zjUi2/40WSYXCwyaWP4XkXsc0xrsoVmHsv
PZuzp7JB1B4ik6qgrUidIiQLeZAeh/swjfas8/zDcYQkhM3T1ANlhJVizSwqt3kz
KZkPhamGPgI0gddycYlrTg5zoDE0/OaeaHp8dY7OT6Dv/9fWuCDv7VN3LtxP8L7b
zM+ZpiONFhlBKIDPJwowAjzySnUUrb2rPbmCkD/pIcG9aupVAl+SC+5EVthHsVOl
7RoGPehfzdziCjEuxRQ4mYCfXwyYWmI4qf5Y+2ezky9krxKNkgnFXHzvswmdMhrd
uWcLTzPCAQGpbuj7MZoG63vsMPK+FCSeBm0Lfasnx5PhO2eiCbsUlTp2WfC6YzH8
p035pKhryvTxRJpXp5kmHIsqHtPl9D4LtX5KAzaNR2wNiUgUXKFP3JbIJJj1lJNv
fYrFEuh/znTTM4Mqq882bl4AGGjcdY1vzkGTIF8yLnwkznXkDkTlr5g8N6nBu1Re
lfl9AzdhfCBMy+HMZ1+UNmKoeif8rhW71p3uyIzPPDfMoKdLszlTcklU/L45L+Iy
WhY4uohyU3Mazt20e0htPQzxBz3M+0YsZMs3TiSpWPIpePUiTwtxneQXF0QBg3k6
vnEHfyfFliBGHoCwjmMIiU1VJMqxxP52EiKeYRzsefUPw3hbJSEVOcLYqW80eRuQ
4amE1kCCcc4JqqPN5vfqWfCghsQNsucVZl7vEcXnt77U+SPvT8T3AHzGkEMXoWyt
vcpFzOeA6mhFqkZBM4XpfXy5736be9/rOMYA7bVeH1cUwmJ0DcoGaO9SbNj1Za3u
AQUVDO7a5GeVYG78iNWMRkYjUAV+oCgorhI2vF+vb6w3Xhsf74j5TmhdzsKaa1QU
HAFcNzUbmQebOV1wb1dmgO4fbS/LzgrGJ/OOKfTzQIgE4YLj8usgshqnGBd1nhzQ
/fxRa+FhQbTa91lhGZpSdVF98pIN0gZ2Hfbl4r4i5Kd/h/6CCqMIeHynhi8EvwB6
mw6l+Oil3ViENlwUuVj7pBC0+nXf0BKKhfgxnxK2oCwpulqBeHjWaLjaPuRg/FY7
xDXpOwJyIZQTG0NtzhtLikL+9JF8yinxM1dLVCsLA/VAzvFQy/z6V8uFqg1tvFvM
ZBQ2qP1/OtN3p15GyEcg/sz0vtfjVHMEHLJugpC1Z4IX0VDbNfeHYs6dlQQ9PUz1
2YZSL1o8b/dDkOs8il0VsWt/QAyPhbmREZsa+zSvgqW5R5v30ubIAO3JgxSa/13Y
MGoc/swpIcsWA4PXh6A8Ji8WXOmQpXJyvTdG+GitntXbGYhMI/cq9+NrK/f2MpNZ
M8MXI8Mq8mt0d70jw360Aiz0yyUeI7IL2CV/35pfPgYhlzmtCYtNQmUxPh6b0Jeg
8X47znFegUvYAJ/6dFvXnvMXlvKyukhd/Cb4Bc6QV6Mz37IgVWQReSrxbEalAhnK
MWMarszmAyfKrId90aKbFnZRoa3Xl+4E0qKQ+1f2q5gActvUO23afEOXBTRaEVuH
pwNwc2VhKDUJhqgpLtaru2RztrDHv/B881MlQUfiQ7xzjqxZRsRgW4L1HRceOUGp
TemjiM51ifFzUb1pd2VLuGA5SoVRGh2NdeVTD81Kq148YK9vMBSy/eLXT4s+xb2R
6h6MPpFnL4Z2wHQHishdMF9F10bjbKtBj8ii9xa2XfHVvFM80tgfMwtI/faZazN2
/L8Pknzbp+lE0U6SWnDXKhwhntPl15zAKDS+OSP/oU1mR30Zi7SWgo5n7XoD99cP
lqXUvEHw8zKm+ofOb2ICRbcaSYgWox9EE766aHvghMVxLEboQ4/6LL1GJTGBCNFY
oDDqfsqaUYtiAAAGSfcFA9mdcoNG6JkrGcYvbPjaL0vm9BVT6q2EyYXcXWM9cMaw
tT07OIvcJq6r3WwV2J+2TIXqjqmrGqO3DbWqVPvwb4xmOeK2z/Xi68MKMhMriHZ7
niV3PxF+rqo8BeppjEoty1heBCa3kD5L3Fay60HcFfpK6DNkdSDNuwd/S6NiwN9S
JZiQje6/3gVCnb0yl2UneEVimj0xf89J7FhcFKtiH14v7ljKkkfGK5PoGNYHOH/7
CFKRJtSTjlvrYNlPeQeXj8Exh9gS0rtN6KnU1UmX1ZFzdH4soxQAZ7uppj7wPvMz
wDnukLYp/sbYzlMMxmO1MsFpWwMkYAmbl/FvdM7tkBbJWCwlRefr0jcZJTFP96XF
Z7QLvpIR4FyBOUKyItJ76a4CWHlO/270uKK+YyouM8IHozxrh1CAKjO4q+dO+ZWJ
QPH/axB0IsekyiprRR+aUinL8GvNfTvAXoORvQn9vttE5vNBWCzh/x2OiK/fitIZ
p81qvI5JtQY3jc1rLRiEAaD3VsVTiNlhGNp54nflqFQRIzhQpE2UZ2shAQgw4xkN
XAL46ySlIYxqI6zwfdd5gxhdiDMjF5eX7Qw+j+3EPXHshGUcSXbQP4Cnjd6AoTac
+8QH8LIbQL6pYU0yB+njjO29DhKiJ/Q+VXxNfh/uJr84OxzzHc5I+Xh5Q92SBOGe
tc9pIql5RglmnpnxL2HD3o5KXLTvg0Nmy1QMVMTsjecOGxtGTyFzoQfO0dXDJYWj
PRQl955N1NUwfLbou8Bfv4yQfsHDm+u3LAHAGSigHelTClq2wqJBENIw3P12dyh7
dyVq9+wHir0BpWx2W1Yl07GP5lVekclk7/0HlIBdc7eftvQuPomUqZpZM4n48Rnm
PiESuhpM57DjwaxxK55hbSKPU4BX+cjqPmnExvq1yma1EhNRuXWguRSoVKYcPNsN
ij1npdfeyf1imFLRG46vybRLBElOpBo8YrGZpH5xgx7M2eKar9WFltkzLNbB8fY7
/RwAyrCIJO4dcG7OoiB3KShMkhy79R5JBWnFr3KEX8T6TAsJUXdbSKPjKBrK37FY
tPRxQtQoMIE01eaSWQE5onqUuJzr8+/zvljMireNu6UIOgfjpOowoGjF29kqGr4s
UcrJeo36dPJyEP6iQarwA7O81mJryuObIjpplmQGD17FFiX5pk+v/eamLh6UE4Uw
RSqZO/4R8aty6dr8DS3MXQwwqk/UVrxmKA7rNv9gPsFZBxieIJmv/wX0tRBJVet+
x/6SDDW/71E6Is9p9wBm+jLJ9abbwltWt5+cfl1IarM6BwdVw+1dUbZKFGi4hIFZ
l61N/bA6/HtwS64HevGopzV8bU7hM/+lgpNk7Au+kSozy3sMYMGAs8l5l7PzbBHL
gNXwTEW4EXWZnmYk13ZHnKxanR6cWIy57mDzAKIEXN8sHWfqtdMNInB4um1f7gAJ
sEvkvf5v+NkNfC6CvkpZ9xYXDzMP0Kl/p6C1eY0QjtWgQUp/mBlOrpol+x9FfmDw
9CtiuPdyrXbXqDRzqETiITInodwls56FIgbGcgpcvBziyts5+dFVU8RmQT55d62c
Miq8gMLKU+Iqnm3PZUVnC8YGGTVStwgzQHKylqBth/HmenX3dJwLuP3Zrm3+2g0A
/BT4KVQOV6f1D7I53meTWgc736Y0XhXwVKhWzbEIjVf3XROU7e2EEkmmZgbPWsCa
IAbsVR3oCHep8Xm/IbsuO9JCWvQdXpJUSeIlnngWRw2T7o9a2e9+O2r8kePEoQ9R
quUHqLvD8cjs3OOAEyzIA9ckWZ/m1IvDTRNw9Gc6MFQXRZzQxa3zjWZyYMmWG5XY
VJ5eNchmB4wFQLwp4SmkxIgfMR+YRXZWgX1Y4IgqOCAt8lbCe34vLeNogW3YYppb
64JqiR3DoIRdzvo6JHH15swJZ6CS3AfU0GK7GQx0ykZMjAeFmbrfqHNBaykKtX31
UZ4cegpdOIsCaag+KYJuLDhSmxurXOVRNB0z4Wd83HcKKMiyafY7IE0KwlhkRJcC
BcgofyLlgu/zyukqTmD5vRjle4tGRolBeUfv1hBMYnpul4p19tcLNTU5fbZSIL7r
FALuVh+L00BGNWrdvBJv/c1uKqGaLYZi5YzQEkPTJ9dCa1qowlfmhwzBwSHWCbad
Sotlyr4+YIc7BIXcxNqAd1lZY/nMT8AkBVBPXmBtOWywbXLzsxOasfsDHdU4h9XV
7dfBVPgrmgnuFYpUOVmJqJfN3k/G/arjgD8+fMvGjWoWFVHgZUE9PxeZukFMaMQg
UwxqQJPd5gJ4325rysdVlwzirL/6BdqPgThWNhaFnEVrm4V0ilDXa70YdOz4f3HJ
a8iW24PaYfXReEebKs1DNETGiGkQ9Ne3bt6DYtptpzURjz6s2ADCA/bPG+XrB9SU
lNuHi47NnZjt0zsi/MPvvOz2pl1+3yZeus6BeTJ7oCm5f24BoTmyFSCKyEQkfHsi
gHr4fK80HXx+C5Uu1KWR0+Z4h32wPA9F2mVrsV11dtkglHYoE+TlWXyyET7wOVQ0
gXusV32wUdTVClIhiL3CvOyquVrLD415HQGKkDG1RDM7G/z233saPvzPNAOMG8sN
dBcWQSKbEfIj7QSIkUBDuNig1/hJyVCtzbts6DHYF+5iG+WiFFQWmoM+eubfaQwj
0BXCLuQV6VAeWYJtGcNmbHZ2koyw9aMQoM2JCX9rP3iaUvWQKeIynPijnyp2+x4r
Kcj1aKVVjQJlF1d+nvbRwQtLfO6O66OUqyUof0QE2smoyE50NlC3EFC9Lgb/Ffgn
VYwGq2Iy35qjWwNADbWtuC3dnA7a1xtjUomKDz2DaTIITr/CfRmQqf08drO0nwpz
0Uk4hApK0P/U4nbd+8lQmcj6IZuH/Z/E0xY1x+tHpDuqaaZrWeDKGCjo0TAUnw0y
JlJsaIms/Ktp7w9txrRyPxqfYR9vpluMaIIBuWW4cHOZv9/X966ekkzuHB3XI6sS
tYX8TAWg6ljT9VQrvSl+v8q2YSvg7R+IcFUbVId1OZwO+RLh59zSkBAy+AAA4kB0
0TmY5sSGgNLcediBmbtcTUENK5FwM+UQysaaAlNlHTeUPszsox+n9yPqJNSUsg2j
k9OSNtCyNY8CfTXcVFgBQUDAI1ccDVnZfRw61aV3t8bHhYlEPG6NxpJlMU2rPWti
OWq2nExnu9EJg+YPmphnyuqVh0NAwxKmkKRUqAy8TcvDUgqa3GISXGZGvnaW+JEw
fZYamCubsTT6LJlMNhAZ6EWWdy4WlYThzS2JcVGGYFjMbbQMAc7NUE/OlSxYx1RS
4IIna8tbUufP0XnVnqrHfERaYCwG4ksFNmUZj5AHfjt7M5SRK4mJ6/T5hCLENJOU
HljkGnPpj/W6lBGFSQ2dhJkPTCR8AaO7gvgwDC1rWYFXJT7VbCwUJVzlWEGffNF/
560j85lR8Y2yCkwIIR109tfF9j02V8tq0Wa1MsSGA7rNiD2XUuFu+BO04peJ611o
naS5CihhT0etZVx8//obv6ibywVtbXWkrjgu+PvRWOCta3KrGYpSqwHTyS57bRQF
1q05wZ4+ps84N1Pt05wBVygnhK2jIKVuk6/0qtsjVS3OmNaF9DzxKmJS909UUtzb
VHy9iMLWrYBdlua2Q01yaSBDuOOxyYCP3z5tM+nW4D+U3uKw/uz2YbQC8DfJA5TA
bjSnFheQfXZtnyxQkT598TycZ/LF4ST/892WW4cUCNZdPdaVO3xu/LUs5hkXvPb7
VSawEtEq1+0R+lGWWhfAqa417n3JXLpRvH4jENYUReh61uDpvMz6CpiqalbOKd3O
WSAkAlQNP+aQZY90H3bquuMT49q50RYG6rzOWtuUSIk094s9Cegg2G+KpKsRTkGO
yhIXF3j3Kcs1iS1uuePQq6qBuDLPeeTwm4lCsESzEIsFpjGkXDF6HX2Pgn6vcRDM
O5BhwKaaPifJpLrwtkueTTXdBnJblKP1vdOTCHVboyyzUXl8cb41llZEU4DwnXmF
jzFrw6ze999ExOwd3A+95deuWOZ5YSEs0iwj/6+MatOVC1iaO6K4pe7NT/4nine4
mljRkwwZzYoBECMdT4XCNt774qJii1N2WdrZHuVCjvQOwQI26x/x4Osj01XlgaXJ
ZBH2BO+JMEUeDER/11Tos73ukW/dUNGPzTqxJILKL574vbLsk444ahS1k/2iS7Cd
fs4ASmxEi+hA/WixHpd3iLJBZ/D96RlZYCyl93B7zrLoukc7HElEIDMkA5TxXEDm
+J9mjVcd/mSrtwmRmSUaEMTAgnDIvV50nF6tyQBBovhHv7uN6gSHmiCGIj17OcxU
EK47T78R/jAyA2NQsNHw461KDPqiXqRZke9Vj9UNylrkhKwTk2R2HVEHjVaE0F0k
npL0+4I/W3om1n98Vbu7QA7tO/ObaWPf8lz6BRiC15UtQ65wy4fObdOwe4D47mAd
h1HWsTwwpUVAKnJaIZgc4jURK3oqLNDYel4ZMnRP+igoKnn46PKNwgba7STiMsPK
8ed8ylzWsUIOR5Cm5TepkzooNgo3lPxw6eMf9RfqrLb+EyFZ7uFvplYPebJQaDPa
3opD3X12oL9NLGU3sNVLEj+l/yge03QnmGJaYpWkly/H/kHMIhd2JxLpZWXf2i4D
JTGBb1OWcZ5lGgrjpmlpSA+D5yajBidAluRVx4yTtH6ytuptAEz/ZF1WksRAGWLC
uY+Tf4ldRt6Mq33nKgeoDwBeffhuAQ2mhUQiWh61Cbe1gvnPbQnodjNy+yn9M8HC
PTitClJklZkVqa45GPInWYR3GoMasE/5TPuXU6bJqH+X7iXMOVaVRwZ9MypKklPM
TrL0HxunX/GTHldrILPuT/gH7/6f702yQTO9w85yIq8PrbdVavA/vs0NXWTgJJTg
wyE+mqUSxi5a4b+KEm453Y0vwr20ZX8W7sedTzlk53YFgXdAR1Di+GaD7hBY3gUu
huRca6bpWEHOpptNnh1JEvZOk1d3NpIUiC3rn8fu96PjtThDyXRdnmfNyNn1o70U
hdzAhn4SZ0DfRZuzrtSLJg1fF0zny60pAND+is2ZNs5x5dQs+625+dNLMmYBzQ4F
tb8ZAxOsuumiIGbHMWX4OZ8FQzwtZd6PdfPllcVYIYFDXH7rre2+AmFOMfksILAP
E8ezuJhGyOa7qk5IPkXQ/YIoptHhEJJMxtrKBu0aPyL1NFmgFbov1v4WtDS2c+OM
k6jlsNskmNYGNBlP/uCrXyqqRTjj/M4DGStDfj5G3ZlUu9dBimovOHwf5gy6AL9/
zDtWbQiWC2TrVOFID+S5/7oKKwCl8/wZhVV2ErwkpwYxxYvt5FVELZ5B3lw1Faoa
f9tyZzU2M4yBAGlOZeF3257O3t/e3678QJUvEpOTeR37aFEIRbA0xvpavn9b78Mt
NByJyGk5j2fXlYzJGa/YxkW7IWV9Y+7x0B7x33SMxLmYsIWDob30s3vQawTDMmBr
H1fBXIp/RMaY5B6K/d+QErot83IfPAMReb6ni2FqzQA/Qu3hSVgajYz9ZhLVtaPS
bxJzXF0HwWZguQ3OqKf0fnXT/uXKYjOow165J8kzoHGwwnL3JubL8eufsW6Fz8p5
qhe3WpQ69kYZWKJ5dQKejbHJMZmAfaffOqP3jNtSsJrmOO+HAlWVT1XhgItq1g2f
g2LauYVPO2crgGAcYV8DB4RP3fTb9HPLHsr2EQN8+Xl3bElq5FKD37/51umYKn29
sFgFV0Lq2ks6dPXkpPFTSWvvRoiWy08dBR5o910zOH2+ALs1bk5pLpijTbtiSboz
X1wSgyFOAOEvFiURlJoydE1KoQ+vCTJiDzGm7a+TNhab7tOiuDFI8Q7kZZKhcI3n
pClM/J6hvKTVAxu1pweCCNQfSwZtkKSuiOG4ds1RgHwsIpsBtqKYmsatUQjvF3BB
2xvEc1K6wF9CeGRW2B/9LAe1JJzuO5SVhUmIVUU2G0o4ruuhaXtVf9yJnFwa7K+T
vstNpBAG8KkJeE7xpL9wQRlwbe3Fy5jIJQUecNfPBMyhImmAeM2PbUiolIxrzqoA
91TWdTQFeZ1ZGdlGKDyBHQMzSd7UyioKhM/+ARsZhV/BMJa9wwM7HEBdCrmbBvFV
YcMIyFvA40xmcKkSU6c2ZTGBHhnXscs30Ff3pTmFHZZT8UTiuhglsA47PyA8wRRF
xlhV36hy6Z3G5A9fD5UrE5TDhi9onkOAWbx1snkKtQ+7ezfa0jnxyvY0Bzgh+kN5
+64FQqyEy5qEMqiM1h+LJwCLgPqCaotf0z+7lfjTiNcifZVjfkZiMJP5WC3lMtjK
35vqgs0xJg2/7jNkYG0CpxPcpK3aoi5vDAvhe0Qyi73Z74s8juDcLEJCROx6VO9Z
WdCl0v/yi2NYVhmVUASjT/TsDALyvicWs9YzdQk60Kkt9+zFg2kE0lACUTsqgAwj
UOdyX4ZVxPlUR7t+L22DUTb6IsVs5mqwujEo2c8WDQ6mzRgGrsPqFxswEu6+UhJ/
b2d/jSowSM5NJOOkiMm/q0bpdD7M8uGrltuCg3WvY5/he6+UYtlNWphx/2mWujxU
sAusvvKIL6tQuVypZFb3y4yJBAHLCpSVGhZVLqxqtDsJYPiyVEtRmsQ+/yjf0vqm
9GhoZ9D6oaBmX3mabxNECPPoTk6yLFQFY3/uxvpdju51+1fF3+jyLbgBluGcapvm
g/QZBDk3sColj+OmnN6qoNqV7S4NDLSYyvUMIxWnZ0iAYYbJs0LXJfjXYQXAsDx3
FT7hjYdtVxQZogi/VpsOJXzh0jvHoLrByvrabSQeQuHPORP9bfIOiivim2CNfxP7
zMfz4aLIBYqzyBNx+XdK/AZSQdv+a3V7F2QimvpRPe2AKPmY3BdR0tGXhyXzh0A6
0F696W/1TuqfjaTNs5f4BwSby6USIJOkckdl/cqVRcsAN/X0mlPyj08UqtvMgi9p
h7G0oRllpouKqJijbtZ/0C7tt/eIeFDPHzYi04MXEibFSbjiiV7MXOmmMgOPgSP+
RgPopmibo3MrKGfpR53aUDCJX+6DgncyXEjlosUR5wYa6c7v1zdIERPGfxEViPZZ
BN5AccqcXvvb8JocOANk1/249n6Eb5HDvJfFgoXMub1DfUgi/LK77LIihqyGdJUN
rD0EIEKXC9Fv0scgGWFDM6yG30l29tjc2yB4SMCONVqqxdOk1qPm2qS0vzpTcDaZ
LmOBSCja5T4hWdsLROc2r6KWb/H+8zzKVYMkjd1PwgtH94KGaz+kzIREp8V86xPk
JEtuIuYcWMtWtzY1zH4jsqdgi9nGfm2XBsiVJ4IFPdHPJlqJtpDvUIIAvbgPsdAf
XfTac5Ofjp5a/l5V6HXIVRAOckqa2+B43mEccmdWKWJ15G4WRn35PN7Da10PboE/
lMUaS5zzJEaR+R7Zxv1UmZTNJd9UgspZqEtf+YOpyoekChBh6ttoIigP75uBzdTm
tLK1VVtT0WIvpmmk2nyQ3VBNHhqwf97mRtkiaH36IHGmIguBCiV9xd2DLPF9oG3a
qPvofx7ei8W6/JqKAqkEcrCEIXDLPz+Bol7QX1h0sDIxH/HxJ2JxGrtHrXdLcvMd
kA4MucY5Ykj147n5O7+iPaxXkZgAnoK9KnPvxtWUpnmt4wMskb/xgeqycFvp14z6
A8Ly8h4mjqoLEBo04n0ipXroqnlZXOXbNcmCVLPvFdLpzkO0yBBJ3HwHzHuaHIKI
rPj4xjoRA067jWL/m4wP7gPWULV5K2ZOGM42MzzOuxopZfe9xWAOeQGek5hMGq/a
gYuGPPZHHHuXafR469+yTga9Cjq9SI1OAfwsikl6I8gQzUVzThaFWMmDxUsxSZNC
lkJHiYrqraszyuhMURbjij7c9ZzlV8rChlou1/RLELB8Qe9pNSjeCxiEg8oCGmKU
hUpr44AyOxoIBrQhVJVS9zvtOq8qabDm+tUieDKJw2ygeBrzY7LFUJnFK/RKj3FT
WAGOXl1dfjQrIsvigG8rpNknW3k4ksRUe2M8YLy2+290SI66nf6ov6rrEHaFnhig
jjkBwkUhsPaH1RCFA6zcLm+7oZUTovH3HeVhTBemZQEbj9Urf4uMPZZpEdWvP22P
ve5dyT+M+INGg4MgxIGqDI0V2F7BJrVpuljmm2iBrGzG8bsSZ+KTdaG9gifm3dhH
syaemxjc+0IUMr3Z1DecDw89Uc+/DT85NNY9MlaU3QmIG3ZMP5kBlbMYwl5tKm8a
33+Ebl5f0D7n53GmuDRaleArdz5Vsw7K3p0nZY4DJxk0GMOWQPz79DloFayYbSdN
P+cBM+fjz+V9xRPvglcVrvlPXI711NUNjRjNoDry2cy1Ip3urGTLeNzMUf6MlKtV
f7e1C+EebwRujS7qOivZwnP1Crv+w55u+P++APERo6kOefwo+LpZqBoJaO9PXS0q
LrI57wil7Q0SlwkQtaD9JvdZq0ZSzktfam5glmQAI22SJi0nstKrotqbrFbCKXui
zWW8/bYUc64/KhCVvUjjrWuhCscQHXxvSlxqOObqgU2db8xV1IRij374KDUkU+Wl
ipKMVPTA0Lqh+t9qKR5bXm9l4F/io8EEpBvuQ96FNM0LSA+aGdQmBQWVbWXj8cSW
FAqfV/h73zZcGBRkfSRI2Qcy62ALXH68rYikl+VoCVFrpOTaCOD3W+5jRjq+zwiF
8vQ5oq1pLz1g4S65WZk5AhrG9h7J5gj85CPbVPyVZ45RwAhoc/qFQAddgFiNjzU/
bL8Te/hM4BjMdNudkotC2rLsXg4qkn6ae1s+cJaWJ4N/pZU9ItQIWhPUmQKUdfMS
jUqJugQmtu0FnfvBELHjnO8p6uxElIka4hqurtV2w3kDk9iXr3m9rV4N7UqUt4Pk
p/p3gOLyHMG/IM862hcT6Zd8othcxB6Rw9cktRJju8HYbUMSqJM6YGT/JXpI6gvC
92VcpRjRDUv5bQR7BOgx3xu4blrSOSmGYZ9IizRHREaxGsO+C/pFymgOW4yE+Fah
EwplfD7uJK7KBJjDxswAxG4mStv8VpIcN00kaqNxEVw+0dhl7zlxPfvwOBFi2WH4
mDSJGUSx8WxEXUN+lo5rb4mfb9KZKVb2nGt2S/zMmgyxsEbbsomAATk7bBdOaw/U
0gbXy6ruNZRf+SGyHFSyMdkp9fyZbaSW6dLia+ibESjcOjlZyhBprTA8nsAp5p0j
/ILXdW7rzJd/0qwC0gTBAUwf3SEzgnGrQRhPcKOeOjs6AOwIe15fCadErgPwVI9s
NiT6fTkSosa++gb5Q7JHrR2t/wQu8wH7/ZTztOXglEfIj1vxZ9idgYIxjvFAGs5b
4A1HwFavi/Rl7tM9uNiZRUi4jY+gTSMxMji7U6Vs9pUcWFx9nODPSl01U+lBIcRg
rR3UV70qExqVt1AOk5CIPHvUiXOnYPi0QqYtepF1UHzFA3mcDVW7ia+BKe9fLNIA
LBimxX7zg6sUQbWAeiJA5S0JyEmMmzTCjEOHyDHZDY1zzseY72L8NJw8OIeyqwda
eallchYAee1+H2VgYpOFF8tGHyn4d/gU1nhsi5cTG5snISWOPbeIsRoaZK1WgE5I
c4rtp7BqkV3C4FEvJsqX77u9YpqcpHLg4S9L1/yoOvCIBsIuEOz0iyyI5pCUpwAz
8gvCeABt5sXoQMMveRXQahL9BvA9Ggm5TiXw61tWd4d31W3V+TxF8CjwB6z/XXxK
K5oDbjP/KZZtfVwNQqViDYD76tmA47y4ayQibRZoexzperRfW2h+G2P3lF5Av4Ch
PlPJP0lxUw8Bu9lM5u8XfValKC1cQ/ZbZNkTcyZZwfsFA+MAXoBwOwJcIIPCRlgF
mqj+T1HzFKtGjKXt8ES9fDj9+NDk+ghSR4ijU81CfF0/RQs/NE54h8if3zd8BZcz
m1KNKFB1RwWJBjhqG0Ez8cTVVmg+1A4usq6eVzy3zfR/Ram4H05gTTA9XMUoEQav
kT+D4V+cTjZoTwumWmFTZT/FDSc3K+yTtaJXNyS695KqDXSx09ceMria8DYwoLka
Gd77yy5aCLlTO7eOcv2HGqNsZn0NEOExNkIndLbXrEW3qivD+zecPv72JiAriawF
tYS+uzU7Vlx/4Pj5/TTFrKdoKelkOhgEbNLxrGG5CWsU9a1X0CFS5cAOIWDCWkXu
6Gk8cUrW+ZuKHX3tRwyIhYlmPZYHWMHIyeNfaASLnarXUF/RhJWSRP7AAbIgCZzq
lh40kptW/orlL83y/aTgzNnTzI/xsKldq6uBSECHfvoTLZikI4Dy61jpqJAk+eR5
cMtTlqcN0oHnN4xaZzbUXyvA52gUZqKD96n6wm8ySOtlWHAD1qiiWNy5NRPghzSV
9L0KGlZuR+b5GqCO8DIleoAV7/fQ6XwSc2M9GawR8a4jsJMIuhQVHheqK6KhQP3O
nR8vMVbOF8SDauyLdx/bczxbT3qbGI70iOg9Ic66CVxMSCLMlwCSw3exWRgrr+1l
GPPQrOIG/jc27ofgezkw9/Hdd7ZkfVCtj2Vpve6B25eLrY/qmc0nspPL7M6VlHOp
xoVv0SdDQFcSPviJDYJAXsCqdvLK0dlWdmHkUsbSnjj/zSQrBNpEU3dgdsOY0RK5
cLqSSQovcN7cBiqmGLivnpYYSwWzzTMyFdRxx9+NJKdySgcXfUAVytPYWSu9dFIn
ckAAVw6bnUxS2pG1HDFd5MwrMoKLpUGMT/nWtozb373+JL5ZsdtTJBhWe4dfk1QP
QMM3yMZHv2V51qKVV3Krjm4jCWyXF9/VO3ADFUubON5KAmfKQWaEe21NSS3Wb0gU
NqspkpiUx+Rq1ud7nnhWYCjytmLHzEir3vFGSzsCcuJ0CdtbKJb8AfNpDpoIaPT0
EWKTFNGBXBT0W5ALe+2dlNemMttPTUfOb0/IP844mzW+iwXYWkZ4QLRKxhqlb9IX
XIOHALULnezTmcuvHBFrILr8KcWOfN/bkAiOZQu3LQS/Ad1CJ8LbrEmpxevkPzkP
8j+FfQunDFnpiUmDfJLsaSI3ZRLff0WU08MzzGICdYMI0gGXxQg88wQzNIMo07ZJ
Ki33X40EoyNIs7ZwHN3B63dCltBDjalfekURvr7XlHIZU5XWGGUHTgEQvF0zkjo/
Nc6HB1cLVpQ3d1B2q7ZurrR+z7hgm2wwlSMt7Z1Np6+1Ko8qbSX1QCODs3z74x7I
+rmjBFvPLQPnCFlAt8Ia4GZQxToZYFwZlyqUZHtHZ0S8EyNziBIdIirHke+Tt1F+
utuuRtTpggvaW6w4EIVt9J0tydqM+J+u8dul5sZA/hyTZTfXp475GmkczPaLnGkd
CNT2OaXmj9go8lYvPumdD3OK3HjacL6+MI/JaVk7qJ6Z+q3zQoy8bQEBvoSoDkPc
XYd41k7Yt60Z1qI4jO/u+GASV4YLo2Iis8kfliK+bPYwb/D0jRfVSBIdxRojNVlJ
vaJdZrDAnWtmAX9oWpRly7Dl3y7zkUWwMgqZjajaY2TgiKC1Dwfzpb6edjg9a1kN
1wml9MRPrsqYeF2erl/oWLCwTXb9H4s+c/1i40T54pFH7h+o07zhc+zN7oTDYGkX
v268O6HC82io82wqf++cLuDCWIwF5gQ1iqM0Acbotxy52qxRDM64SU0eIFga+LIl
rc+hqTFOVZwCbi9O1zVQVk9xrD8kHyksUwcib2FVtiUB3tK82bcwzwm6CnHYtA9t
5JGKsCVocWV87z7QEMaom5oE85vqxjaOpU9zNEbdo33xcafleHJVy7Cw7dAzLe2a
ByoSr0+MD1QhhUgXKy7U0rPzyAirKoHnlH4JPBoBI3neJH33akd2zsMvXy8WRJfR
Owidh+fSQKZbJON32jRTSDkquB/yFleahIDB3FoAkR9myC5YBA9nWV/rir0Txjiy
D1WB4DYhfgMTvT7etiWXzNsLlZ5VhCdS/t281JO4YbQ7Rkwkst5Ky/XIxTWMlr6X
yt39jJleN0up9ibzXmP0RBLbbUGI9x5D+q2eoDDo7okBDr23VX1WE9i139knl8Uf
B1NxfAiHNnXEPBgP91bwzWSIp2QknXujiCN+s9xj9RYOjMYCXI5gx6wSfgKr77WX
D29zoomR9/5pT0sYOfTaOaYGSpsjvaex17dTID70V8lUSSorWVxETE4wBaw3hej7
XQPwMNYH/mYahC+9C1RWUjtEZfjsdU32VizzoHoLsK96ipVyrmwni0lBzp+QP5uv
jUAg2ywAg4yAWEg3jyTaqnTse194LQafU4+FdAc48i4ThiG1mjq3EWloJ/o9khtw
3kBwt0XZ8yl2VB4LOaBqNUcNtTQAsb3mSwlCbVThKK5TMEXVFxJdpakX/pR5BnwF
X7wJKbdq95uOBFXnEZyeYqQc9eqAs9oUPMfiqUm6lOihb5Sn+Q4P9DC3C2jaze8o
K9S6fh3k53p9KqRIzhYhdo5zNesXOEInHfeJU902GSQ04mDSOUGWMtfEVq26Z0vH
ZsZOtkZxxljBVZ7uN2DNHXqCSK1Y2fHVGJ5V9bMubKiO48KZrUVOQ0nkaLOeoHqo
AukIACnh4/md1hOa8HEJ3cBzi91ENBJlxMhwLpRdpndguOWiPVhpedRFceuiCGdT
dmhXGsuX7VGrWrWzpiMqWdtUMjZc68z4rSA2qQECbj9J5cGMykJZOoPVp9n8f8De
oyXbNCUdqfoOk3wbMyFJUqZJZtWlvKcQno1fyLL6lI2UuYjErwscPSxvjDzy6rFj
vBvJRFGw3tm0Is42IwnEL8JFq9j3Jiyw2kZQwykKRnkNwyVl7QDOPn+BtQ7Okner
4Kq2fGF38AZkcuVzK7jffWSJyJ1ojZscnsVELWzmrjLGbtnhVjN5TG9oywIOCNuT
QaioR2eIgXJOGJIofThAExgABaIX+Ip9eng0ZxWlgPWVc41308jE9prlCuZBlIzP
X9khRNSv8yvmIk0qeJm8czF5t/YzOG+H89acbiXvyV3xugZoRVg0zBQguOLVpKTS
oPjPoKXf/a8HkX7HL++NEKHviAUvGULTex0NCl9/Ksn/kOnO9hbHC874Wu/FECTH
MBYUPTX5Yp/NYxPnsVmnWKDqi2HWqP9dSu8fTJHNvhXkscMXYzw4XraUD0wDQjyM
diV9qtYt0g47FJ4pO6/QimL+L/7UkC+xCHzV3jCsJmkHJtKg9te83uMZKsE2JmN4
PcPh28yfzeekQBGlQY7ZOHvcsSJTrLNUVRaRQ29M380u+UQ6ZUjqmMHBryUdJ5fU
Z1Y/lNExJIUL28mYhIAOEG4hjIzVxdRFjMqcZUcMxkIwbMcWIvj9pVO9PucHjNZf
WGZVjoJrEpYyU8cqzF/xNWCDYeVz1lh+Epd5DO1SlFHr5b+NYr9M6euS5fioYHwa
H4EAw3t4gMXyG7NU3l3GxwCMXYYV4z06jJFPhO3BBC7MOHebgqwEA8bxN5ExzfE1
Ar8bbxKJkJ/pjatfriQbl2AmIKO7AYz2fZv+dFxf5VelPNgWAAvy2HSdfc2xOSed
w9O3AiOF3S/BpQrvUN3zqi5odjDcXaAqmtAVeMDatFf62dLt8YqRUuuizqsbxnb8
AN8gXIxLDGFDZZQ4fNd8BirVmKQd+8opQujXL1hK9UMfmZIKjbvZUbMs1ZOvGAfU
lNvjDeyIBmdwnyCqoPGpDPl/OHhM51EcycgiHdPzD9anX+dpqvvd86tCIstIMbn/
wjHPeCiuSsZcf3w1fLfX68bkm1YxODA5yeHdoTTkkmgFYDs7w0Xl5SfuGLZKSVWU
6Rk4qPFo41DAtbAI1Be1OGxx0U5yCBxxXwJUl1KkcmEaDBdWtZMHPxR6sZEI1NVA
tg1PRQaNpj4Y7dxRp1WrNsp6Eox9EfDWkw9NZ52FCje8DgiYIVy+dqfCi0YnjpVa
egDoCHOgrFdPIVaQi5/w7F8RlAhcDru1nCi3/IF4hTtc11NFfRkgasnQHlX8JOHW
yKfVom/lLPIUnPciTnKbtaGdiW++1JnivoQtXP/1s1SFbRT8rVFw6ippwUQ8qQCo
v7qhwL9L3OGXBBQDiKjvJ5D9JZKLRjm6hd/Nd8beBAXw3Q/i6oc5I1P8C1B8zX99
iWpFLqNptbxL1t05IQLe+t/2YBYa8eJdGCBI0MVBBV4J/UMzUfbbDk5b24Tv7LWg
FLbrVP3QFZjRfD6cdDgWlqdsOm1JCCf+W/6UszMjk0J9xMB9x4c2bAXycfNC3tDi
AcsfDxDF3K182RDSGk+hVSlOvjRAmwcLwHGMs2yooJojTsg6ZFHpicg1WlNxR8Fj
0jehZo0imKmzoFxqgmY3+hWzazAs8aCzMahzLYYsm6PVoUUJBqNFRFEYzGe62r4j
rKIHpzq1tGO9Bgcp+GPg6ukK3EXJwbPV8eerfYq8iCmWxW6v6pc0aU61Qlh7u82o
mqWNzRbOWmg3O3wkV1y0vc48HfyDZ6FZf6KvxdqrWnmLsJXJ7GS4aMbbZ+Yj5nXu
kkjE6oE9oD9HfBcY1tuS6Ba1pTw3wL9iNsKgToZLTjLXyTdvLXQp7Oca6HcNu7Q5
tL7ZH4kj0ooNgJbNeIuoVlSgD5lzZNfnmFo6HqbjkZjhyO5xI6adYxmuKTX5pYMB
dtCx4WBu00SyQ57o5OmR7z2atPce8DLgMPdaTTiIbiGgML9Lm9X/Ua7WnQ6xgFxU
mXPswzBSSBzK2GNwzzsz+a9m54rBWhpDuPyQLmBRAwqjAqE//hrzazs/e4zVLKCQ
1WoBb434hSLI70zN8G1C2qHvabkasQSX3csFyuKYvFaxJsKhkO/MyW2imOD0zApF
sfpAT0K1vz+Uby5tNWMuSQalou2BZheZswvm6NJ5bI35YwC3/zlKn2++KDay8tdt
0ua8JsWllazmQyyOtizoWXWj3hU0Y+Dy3gCwb+D7NK1pdzqHgrZoenD9b+la8UmS
6xPdOv3DghWpt2HM7ArOVg1N0sy9A1imeaRa0HrBdfwCfhgJo3HvQumAps1ZKGRI
WXYv73Zpc4c1Swu413gEkVDeyFold8v1YPalgkc9XmBQW9apoFJI4VeDfq6UxMgh
hMYkK5mbN692YQrGomIE1VLNQsBp/A0bmE2Ga30Bqe15JqnwumQm5oSfyBb3h6Ld
LrzWHU+VcF+nedhP5JF58DKJ08u/5dsfFQj1Rw28JZDt3wIclo7y+lS1gITIeUwY
H/OZzgFYMHmNfHa7MBAoPjav1GHm0Z84h1BbdZPpc/MDhr8hU9sO62F6ZW7icYXE
oaWcghkyxJ/iISI4wToq1Odia+a6MEcFOo4/zXO8RPzEXIbit6rirUKIrITsezH/
icCrDIW0289r4XFqEitlqu5HNcfnTQKsLWoA5XjXOkcWPF4jvsmHINHkVzb7rCid
h49cxEmcd6lLWMkNZO6p/pSPnOj5w/yls8El5wqEeu0lWG6SidOQaSZs4tFaW8mM
xU4mmTMl9pS92zVMCYp6R7jx+hdDfqoewpye6PAK72eEIIXI2fmXx6kAwfz5Nh2e
sJInD+4ie5ZnVf+B7QEOViPflZZR2e7tOvjNdiMjDpF51VYmOEDkWi2WknlXubVw
loJU5Mweyo2zk0dp+fHPzx8EhnJZVYONuO/ORlcneHT5sLb2U2dUqUaRZnq5piqW
TCXPaYuZ6QX/pMNlikmL1lTp122kNdSvvH3H30T7w4//vGA3IBY0aZvaidqLMaKA
CUpDAbC3oxTKXVYri9nz2YpVYj+z/+7l4zdZFINC3tDiFLP2KwdV6C5bJNYbZKVU
bXdULMkUVMutZbSm4Yq88xK3+GqgkbCkEZX1r9PzS1Li89yi8yQQ9flp+e27bz5b
amz3qeooF+nGdChidkwL8LRSxFKaX/DGYCble8sR7vxqWwww2caBzzF9m5e6GayY
gan76kBv9gZVUgl/QgmkOUGtt17m0tzLcoiZ8jS+ca6zT22qoKCAWneNNAqUYRY0
S9/7/7zj/EBMjXP6O6tZO7zZbwQRWka9R2HurOQRfLvVLvuddQ2PjKsYHSPBUo80
OpiG43kIQGbEKRAkm7IqTkpVGZboM3ocwd98bLvHoURoBieGwW2V+AYagPu8//sG
qiKnCu+EAfznDkMVgPMf1fJwHgGO9XNbq/zAS14IvnAOSv2tU05zblr9YWUnRxs4
N6ZXnVyE6VsD3yG2Lk4BPp5qDvUuQMyQhZ1OLCN1aMLD/ddfC5uUAkMrUD/ASIdg
DRsNg0UTuqFqLfZ9UKQyiaL7r6apzdHCNA4Z8hSiDOFMGlQjd7pXoI1shBbujNjE
XwvjnDLSgXf9SvlI6D9XGoSNJJS7aDHshPw9yOBb3ipUjYvTFM8AEPqPPkQdsEs5
GYcg0fgwgunT4HTVeLazZwn6/c+f/ZTwlBt0sk8dxd2BAB2DFuK878L42338OMgj
fxG2gjsoVGFpfQJBqk6anj//KM13MiCcELDE8NKwRwVcK2Xxa6zLQ+X4TSlmfYs4
/yMAm9vtgCe+mLuz+Ceu6pa7h9wxLU9ah5LMet1/+1hft0WoPjP9xNZhvSOe9MmV
koDkSNBgpBePD5GLQkzR7ExMk0hKwhVBNEWBrpqivs/yqq3CzeaAznsH1dhqT8jE
aRScFSCSS2W4oJ3idaoqUe4RnbfOJqg2Kulh9OfY3hd41mnGoEYXzSRGl3uFpXvo
R9YGFGbmWFbDDr1FiTHI53UzE8H8QjA0klzxIoZTbtCB2HRS55GwV3YEyaJjqQFk
jyp/gVl8VVdotFTG/NU3qajkdqOZ8BNxP3X7KySjBEFK35ljK/Dh8KM+QenRHdaD
qczBC6eFphH06cVmTCv2AhPQpr09xI7wjk5W+nTtBTrFUNL/HafN3Q2pCiuAIlM+
vnuWJEcsF8OrgOWAe6Dkq2tnqNFpvLnYak6b3qyAlQPt9yh6HxuuFwMej1hyOxEe
JXV9Isv1pdwld3xx/Uufpz4cB5anQTDmjok9M1OYticJNiAXXcuABErQWmeEAjgi
uTjdLSpPmukcwqETCJtYLK7IB7aF96qauk8rDn6b8tP6gwBP/eUSDfPGUMFhy5zM
0myiiPGIUebPiNPj6yByB86vU6RYwEBtjFP95D8ClSg99GbDnzpzb8zq2btyRb++
Q5LRQlNdrUkO4nn4fe24KE9ysF+ABaELCjBwHqgLbEPMKDASoX3d9C0lwC+5RSAZ
V1emT/OoycnjLWrbC4TvhcUdN8BHNerzCgcZHSuaTsxjTtaW2LHA/sfLRAe44rLy
3Sl5sCu8z1G8MKAr715gUPSdzOlrdP8qa0lB/tmQ1naTAUAbkm59xggtyTx9gck5
CT3va06o/d4hA8iA0e4o54ALnqkucK7SmjhF7o1vPajoBSjm0mgme3WV/VK1d0mn
purXWL2Cvn1wUJyPjz80vlm+EZJV6rskTX7lV4O4tVIrb8JTNyWSIbgDEKswClII
7MVFW0AS9TXjkBPjCq3A3YacSy5WuMpm1squ+JlcR55Sw1vx84v/RCZZiJ9Khbag
gImgpBeZ95xC4r4RoGSdoxutKuuej0s9QBB9dH7xrc4SOTw+d4ZU1Zmuf10hWNUV
MdbdxxCZD6v1+bzMXqQ+2MZgUN+iPUGb4fU/M5MXR2BuLC2+v6hrif+yQmjLwADZ
3SdgZo2LMDiiYd+J2gDgy1UoU5W2HfvDCMwCCWpJu4If0fSrj5ahWoFsymL687Fh
hq/GRgv6h5K2v05hnFubURM80OydFbWM2OmXQP3NRzxChu7neIpaYTnoiT+DCJ+t
1oT3BPvHPqy258JBM398c4IYqBR4VZkqeGmFO1nhDxsgigSZzvkveHYqaJhu2VYa
GkRMisg4UzK9nBdeVOBpDHZDqIV4orRUIol5tg+Bc9gqrW2hyIsOOGES8gPCyeuM
kDlL9wC9jlioXrKvSKcNCpURQ9iYDsfkDqzARFQvC0D8zJepzTclr9Wfgh+spr/i
R2+aVSsm026pDlrzgznApBlUQjNRvqL53vfzPMvIIcv9DR5Pu0HonDU0BiCKhQoR
f/Hu7xf6X6vtH63whrEPP8v/ENtg7QMCUNhCmN05gkamHwEbWJL60GfyrNeV3U0N
KPYxdgfENqdsEkDx3Mii8iyaNRozQ6NeGBfXfx39iDEO4NQKt+4+FrIEF59Dasgj
z58E1rnp9DKsCNPBqQ5Le25OXdDesh/h6K0bo9fNxZOed8TZuGQMVe4U5G317Uff
D/mnoT4yVdeHcSPwKSheLuUV8VYuuwS1dlGnBmh/u5tC1jyCV+2LsW6wmBOJ0bhf
FP6tncfQwC7cbL+ViwC/zB7jQJwxNtyWAuPWhPYsGUN34z/fwmDhigLPxmV4hWuh
GJKWekLMJ/E2yOxEetkrTE7OCbVbe4RezlMWtEhP7g93jKvn1//sQjdWufTGf7Qb
Epo1OVUMtvMpu1mXfo0ZOIRJhortPJuoBrvO5cJaXPrNqeAU9GPtlMo6UY7C4QnH
ZfezLKnVioIg3EsC8vEPAmfJG2cTz1T4cFFJ7mNYZCIbYTTIU/8PqfY0UQH9RZX8
Q6u/CJu2BfA7+bj60WzU0rSml7vs5WLZD6D1qzrDyAz60XPGGOmYbg00tzMelokn
j9stGNcR/Taplv5yMb8NxX6t3/Rh1MRp8CCBjsUECMT8w309O3LwyUMUDwSDRc5U
nAGWz6x7HNrZV9+SELmrT/S4daTRXFQlCYcxe1ZNu7BGb+4EhwH+comoIvnp2ks2
93BpVfmCz6cGhvvspRFPaCNOlv9avK2GME9vZXpcl6KhYq7v671K7JfYwmblsdnO
6tDbYDQkWz2ygD/fuiwYOiXEhqywbiZaJr1L2Ahtvqf9p+/vTzAL83YhcnjaAA/j
1ZwT4lS9GokPMbgcdX8JqCR63rtKollmrYIUrK1kKr/RBFDHmbRy09yjAhpR5GHO
MWnQ4ApbokqQhVnp1cYFA01P0FBT0ikpsk5i516HzpbfoH/llhVZChFYaLz3CTj+
1HyIMgeJEtvck4ygVl64kzPqsgpBDNQrxeirbnVk1PTmnLuXWLtP7Wcbg7/R40Rt
PYLIYdo6TqdlFTYXD5vnS1e+wy1WkNkNLJa72MVxhWLAwqWt5I83+uH2MHv9Z4cw
vZoR7dekQoA+7IhZKav9wiGa5JrjTlx8rFQIG0AvEtj4n/wnXrie66lw8C3XFQ/z
rRnwUJueMpxMGUu9aiqTwZ90K8S03gZybPGgXgvE9QRYHXx94ecRGFdGGw8rU2tt
B8TmKZGmaqcU/YcJKr6XiZ5tPZd5FZG5VhCzC5of+xl+/rsiGN8sbbpBF7GJt9QL
N5gZg5hotG5NyLQ9TiGPBJpkCBdd8mw6qCPr3OsZFZ30b3DTzEdrDZjRE4uKat7A
eIYfMlP4EA+4T7yotbyIHjy1ZZ5q0ThFis48/lLQemcOjH7MYWEmCe1+hJ+eUMiD
bnaKdIPMRGp2pNQQCRQKtaw4nDFkTjab/nvwUEEOblFAOxRN11BDqYak7ZW93r+X
E0Fe0aqzzgMYlpRtwbiQXdyOnpgdReFUC3RoOM9n9FkVRNMtW/wtNTjYQpuFgEhF
ycUYbwM/ex/WX9283EH9MgbUiHyKXY2i1C5RxMwjMynUnEiCx2nA9Xq4umwemh1Z
9sKvaBCLT1Qm2fF3zfYIkxOk/CY3pyivAbTHi71wMHbZy2aPoMpIFYwUiJ4oz3Aw
7JVixehAF4FwxyBNVg3PgoWYKLS6Yygv0+Ll7OknqZJXJ1IhJcaRdtLKxJbZ43vU
4g299HeHklxzSMhghOJKRUT2Tzz1dEV4YkVVjpZBcBB/OAWYSkSh6U4U263NnmA2
i7kWJo/T7bFYfumJ1NSG5ufXpQBOM0FHrVldGFf8Z3rNtHBwJEXXj4ccq/D1PDn0
h8Hk1S0Lu3YUQfNX2g2IcL537gA0I2vxyfPuLJOUEaSSKA4CleiYZUVOSmUWF71F
HhFo7IQ+xunwL/SsRv5kk37MX91p+mD6QQCpCKNmZjZbuZN/ArCW78N/4ZV7KSu+
gZDgdps4hJvBIarNOCjw0coGoV2W++3qbz6Ftk2e4aQ7UHFE8f6EXGd5sm951RKz
7dfrY8c4t6lBrsdd+UyMuEbZ+2RfqCeHcsagHTKnEfxWHsMEPUNM/JS3pICZbIMg
liyI+GybALxAySN9zZqjjNRrSwnNAIarUF9ts6ayGsnHAFIpLJEiR9LZUMZpa3zU
Iugz/M9IqjL/VgQiEd5eznLdEroE9QCJ/4P2H4/q47kvxpYZW67IpyX19uvov6bA
6BdjXP+63t+700n/MmLFPDXNS3WgHe3i0DAos1Hemng5uo3EHrau6R6mRXiKvHGl
8hq0VSv21/8vYM/tPxnYt01KlmgX/QPZfKtv1l8QT1kUKifZTw3oEoFGKsQK2h1A
Cse5qpOB18iafqzGobRzBv1YvH/5i90EOPMugMKuNgbEbLBcQMotiRspyLvUNRrb
+/mqWvbOVNG7zM5KD4x9rNM5kqtaljsRqECrI33MbovP87JkgqvKK09s/mj2Dbk5
R+xw1z47lwavIxlZZpHTYMl+4H7K/B6UsLFCJcyDyF/+YNqKOSAJFfMQMT/4wJ3t
uXFP2HAotWG3rTu9A6QHZ1FSa/aRifp+VQaZ/MTvuK8MYLDg+cHUGAiPBXe4+gI8
E94zRob025Wp+R4BIIWE9Nl3NS5Cd1Ds8dVzV21x9tyDluOL9fKdxiAkH0CMZ4Dv
g629TIxsGcxKta1u/QmtlAfyQnLyKUq+ddaJ1ftfDQB8UGXFCvkOlfRikP7uWdnY
oWGFiLY7PEnFH6PiwdJKeM/LcaT35/Qfd2b5pazzZzcZhAktqVaOMKTv26Ss5/ZN
A/gqCWeStY1ah88ZZm3KErSG69lp2QR29nYwBQcS9pLsnaSElLWweAThmaVKonyL
+Fn1Pa4Vq/fbVgEK6ix/nzfB0GaW4+plNYmGFUPGI3c11tMKK6nL4xHULoEOZ2vE
waHbTM1u9lnsQxza0hd0dqOt8ZVeYaI5Qc6hObWyeXtHxxT5Qhr4YAA+sgWI2IIp
W+XXCNPGm/m1Sp4eRdOj1pg3StRdkEh+AoRlPAf6sJ8mN4TwCR9iT2gdrgeBwJDQ
ADIdjtUabTDn9wZDe6wBaDwt058GZsPzNHxoqnlcPwHZ7HuCot1aFoGpt691f872
1UcU0S4UrXxD4Tf34/g5+vtyVJ3+uMdQ9MNLjvZgmorsoavdb58xXBlMzI6LE//x
zBOSKbzpl2u1du+yrP+FHVhS8XeMXjIBT9WgRtf5qNHORCEz0EkvKUgEzYG0KgnP
FjGPB54ysLDgP7FFxrfv0PWcSuPy4NVai45WR83LC6rzF2lICOVdGVPKnrls/1iE
56VEiuLjtPXCTSxotZKOjxlPsn1HYrdop3+406qmpXys3SjzJ839HlbvK0Rxx8fM
dQWZuSSAPYvSyg7FYPUwTbDvmvx2b1Eifl1ybGY0rCUAt5sk1u1P35xH01rpMSKF
pQNu4lTZxxBV+dGNC4qq+quvnUlwSt9fAISvcNqRoJJj4VdTb+RoCbWMxtpWpUf5
ML5Ll+NdQyVvF4EJ8Qo1FD9d73DAkV8I5M0/D/LKHXuKgVOluxjya8JLIq9LnT75
w1qbE7QAfOoW+z7Q4kYdFku/JODwF60ojM8IpdwCJ+Nozd/UrClrsAIQtqYLv/F2
NlEycZCVEj4JejIaJ3GXIa+iqkB+YQcTMQ63dx5GKJPQCTaIaSo3qjV5QPe1qOGz
dvbVBb7g+yA6S8svpykPFNrBkV3a01hrvA8sK4OktPPyYdjd1wFoFweUBVFqxLz6
521n2LrX+Eu+ZoabGJmOg9oUFYU3T4v2Z5lLpXPq2d4fs15C9aSFcEjP6I4GLwfI
Efae7jGLXBNtISnf+GiIIXs9wdle+G+16ZexlsYzC2DkytvsRGO1dCLBBBwTvAb0
e646oLRn+KxTpu8VI58/NuRN3AU3sSULduWd+O30Ln1rkP6ajCMLQw2Y/dBWOyaW
iOZFj8Z3NjVXSFitbxWvmL3u+uJI/2hv46PYL3MLRfRpNAjUAttxx7hz9c9Uz9ER
Z/chr0r1HrHO0aH9C9a1JOYJg9dIRxnPPsx4FqMHpYo8j8s2Ks6TVcviP7OqiKd6
4Sk3oLZp+kDA1mJEWTY8YTFLjn/OS8AHcS5LCN+48d0E/3TCtfIaXXcfoe2Rwttp
QcLcVN2DaccIHm9/qOVcmJDANdRHPuHtsphbp1PXM8eIrMJv9s/6yx+rrZHPCA5I
YwgLSEP2p+8l1sa68Yk07RhwYVpU5rBzIXu8/KQ5MzW5Ozy+N5kJTEbToeST0jeV
au083RCbCS7Yj9xvvBSJmqHO3Jpdbz3E9pXhKl9+8GUqsMNMU8axXYF/CZB2ifZf
iluC4kdWT3FbzZk4PvKsrm0kGel5NOCuoiQgIjFxhF0mId8hhDoCnKvWZmNw5CHV
nV8vUgddbF6lHGFZPoVZ93Qrj1NklIXlUmpsz/t2Zp7IHQO5GQuAQAdYJxvToiZr
HKXcas3Upmcse/oTV+IrT7HxmKcm+GSKupeenk04RSsWt7GgFAiKNLjS32CuukKA
lx0v4TeQn+SYbUY8jn/j7BtMVgUHAopgMdyhzXR0aSGugKGBh/SEy5Ds00DI27aH
DFsRrmNI4s5BE3eXKMlzw6kqdEjBw//hF3sR8KUtfGvvLt7YY5QP50xKogaIWWDa
2qCm60JT8xVk+cJqrrRHWga4qlCJ/CW6nRdkhy+iUEfcKTY414OusWhFa+WzwvY/
mUh2VteMQG9IMPWkYWecjSKgSonUXswkL5840exjav64Z1TOPzM/0mrsEqwn8qHP
saTrvSlQxxUqwHnLqLBJUg0eFFscyW2u6Pqi3YiHXp03USfxYcqi/TYdbtanX4yc
PtbXB0eoBES6MM+xpj2viAdp+c1u0B/etxWATzi446dvaio1yPCvtrTkouwhfBQa
F8Vsm6G0WHhAy2biVZsGM5vwhHS8kUmCV4zIV3bAN1QkpG/p4SX/P9L1LBvmgBM1
xZPMBF+oGD2err4GTfP/65PRRHAfa/PSI7THumjBJacGyaLuO/4SPlGXuU+TpY5E
PVFM9CZawtZWkB59L5S2QlGi7/xXrpt72kpXPmbebYJ6FyZpL2bc49GFJlW9VBKV
osMOp27tHDD0K1HvDCop09XbF6Z6W8CvqH23TdlFOGRRGJHf63irbRycchTp+jsm
HD3FEfIaQbihQELCUDSnJauuMpnXx4CI29TcRMyOYMYYDB7Nf1tIH/zJNrbXCQgy
aXzqLANglspwGOh1yeWW4yxMtqjaXdJc4ZQFQ2nNyr82XwDzn0WgqnyUMmAMU2Ot
iEk/XfcIqfT1DbshAbz5ycDvUhWU/tUdRyPGNqVJtVMqup4n54Ds1aB/XwjFwCb9
C2w9Zpvx/OJmcZ+zA+y8tRVnmm9JzkmdH200WsEOYkSzZBtFKc9EWZiGr1eDf5QA
Bdzvt775++A1Ztl3jE3sRJ9IPPHsctyxHTh6yZH71lRnuT38WJzWrKTvsidZcfUg
8sDblcVE4546Yg6Q03B4I1UvRKCDHCCd1pOVcDVmLXeFMh67up9OkukjzGU+UcrH
9U4ATgT40tLDYrRRmDqIq3lx6FzaiEEQXkHp6EHFNLT6A5HfUW1PuS628jWzmLMp
PRal69Aq4k//wNyvopw89Ty5xC4eyoOzaJO+XT+oEI+jDJtpKvX0fX0ZGaO8AnNm
CzbM4iujsHH//hbLpeoqw6dATgUE266koU4UtRgvvRDMtnIdXhQUMnzEEAjH1oYs
6ZujAKnGshLlamZvq19lyoqQ8RkyPgk4yW5bct6zekiiuUUSthpcXIiWsZuAga+R
nxvXxf5Z9oRPYHOFcOYl1dUh9B4MFC1pglYWkSTOlAqsaVrl0A3zF+7zwcJk1BKj
jxqbd3pHb3iD7QsgGC9Itncx/IzxFKO04hTa+DmnDX5Ub5DF/NBt733NQpuqPKiE
2JHsCS/aPKpQXcvV4ALMjFZJ74/ff4w0DBBvePR3G+M0R480Tq6vlo2yO9fIA6G6
OnUh8xZgnkLvU3gbyMvUpd+LUC7eWW7mZofrr36uXjcrgfF0uWz/Fu7FsKl9vNWr
H30WxZbhV3b/IqhVOw7oW3QkfytdMw9wdShCiIAddDxByLnuhO7S/mQcUr7i1CtG
LiYQCF9oYLCE2xvMZSUzrAzDxaPZCP/tOmgTcFA3Igj4Ey7uvBETtkWyxyCAA9ua
NrB77bCuf0DyqK2RNB7Xvy6hGUAb8YeukNW9nJA7wwGG0MaIFN1+KDJzzvV9HjMw
Tyr9aty95M1RQTAwE/7RQXGvAW7xj90WpSu/bXXerWpDk8EMeTyHbkeibfyXvYyg
D1hP+DPkA7IJ7dpO8wnjYRQ5C4bQ6AiNlSKqHDvQdYVFLkMhE7DEQ0RYuAihSOdU
9ptai+DIL5QwDbzecnGMKPjcfzVKghuLwmE5Yn51qdtwDXMhAw+5WkxmM3nSfPpr
AIg5Q2SG9WoH/oX4JdB/pUOvT3w0SXkzc/YnpZOpBsnSGkcKOYkY1kTiZHSpUFgD
DL5TVPTJmwb1eAoaQo51Q5rM0Vpn3V2SNVuAsDKrLuEzVrX9Z7vDRA7ozPwdPjF7
pJZuzFJVEznZ5i9oyKfBGj6FgODD7ON6AG16Yko93LLxdU/Q6OdGqDucuUGxOKn6
T2zLO/LuNOeRRM8WKRBb0LXSbOo8TNmf/7IKJAE4NHLN9YjsOvdcfWrw6te4XLii
AIw/HdGTfmZxQg9pUUB+s6e3uUmjt6LeVn3U92vLJhtuo3X4VDnIOPyv8sL3EOAB
lPC4rselIPhGuHxwFdworBZFI9SCVO8ApepHCsIECWGH7/0qisB4LCikCTjjuCG9
xYmBeMstC6ibfoOCCf3dJ3XkTjwRuDB8Bbzi5h9YahYQzIP7wlvV+NFROkwwC2QX
tT7B+xh2qfGQQTOkPMMuVM3Hi10WL46PKMvCRugr0APxVM7YIm5GwCxgiS7Urr92
lszoZ9izPHXVYIqHFm3MqfwC97TkSAGkA8juv43ZeVVmuIj03GTtiXnmab1aqImz
F3g+2SyhegTxh/Mcn/8rnJawwz5L/yn3rLYs7NKgk1dQLE9qE883yuMkT4WVaupX
/43ogaN07XxcIU3t1HyVdGQgfjV37gzDtLdZ7HalL2ildO5CfqYwEPcYsPWDyjWf
XTKKHeHiCnPci0g3L8VIaokrXoV2cm6EN+PgkDrhAf2wTxTtMHGFa/CLAAkP2WVY
fDazJbf4tLl0E9ULRZKxiIkW/iKKt941qFP1MZGhnojpQoo9uD6apH2sDbWT4bg8
6I9Tg+laPSseWVPMTjMc5FIo6IauBI3EYLJ+IT1GWHVimYj4Xr7r6E2pFVB0F3SZ
2qeyN0QUVc+8lwnrxzGt5HsU1sR+0Q8AHOYfiPSMq9Sz4q6t6jYwjB/ML1P3A6aN
zJp5D5i77LmmuuC1Ciz5NBrwRVuBFwbH+Oxt2ocH/ie8EpP52rBwlCEows50KoF7
FWf6KFL2vzAuAGsTDQMRECoMQtwYCl9ytpNHC45byuEaQu9JbqOv1153sWGKS9PZ
sk7TWxyIuyv/sQ/sTg31clIbOK4zl/Q5ljCTmW741eizXcKo3T10c0XrtQT7Hgcb
q4JWJnxkCQeEyHDPQ+tqxpNNwmgemRO5b5hLV+WV6WPmjQdCv4QT66A2KIawaGiY
Ax7o2lDfQ8vHMZg5yc5WuQKSApf5D3uOsAc3MUQ+W4bLAd98b3u3/GDS57V+hAKn
2eSlh7IvNS30PwPo8uIPXgrq04Sez9aKGu0kHe4SOf4MSgBaMsaAjFCS8wM45nFi
8dHxhjI305VGMRfIKIUD7qN5kqFnxYHsjUl70Chpq1+ibgGhxkVncEpvbVOFOR2i
v4wupzUAh79/rlRHKbkdTA83ATBRIu3uFoZkKdpLo1wT25kemj2cGz5rx+2sglvp
+RmJrMW+oe8foFm6kPJ7aCfLSuutT/RIi8iWGOaJwShrxnU5ImhUXBtOtnr23m2G
dmJLkhAILLhHiJ3ZcIlNSwDkLIkHiKlvUDT500HSJBvHbbuVy+MGkiY57Wyt0ZS2
ZijFB0yPGdmTe6OhrU/oFFsSW1pJb3UbTbaLb0hf9x08IC6HjpAtmSKOQ2/30IlB
MmbwPwpDXD7VSKPpudQJGC2FaK02QDp6qJWyohuQPJUDQBO+vX8Vl7usLIGR8NFH
pRak+JP39cXf2biOuycGGuunkqK6oqnC1m+rDbuZkS+YtJSSBZNyAoB3sI5wxICM
c0+zKkhpYBg2hQjZN3x6NVtRABOJuH0/193yJqZ/E8YeQjN6yyastOZC2V7IZPB/
+LYKwu6wcHPuIxuzrpym9j+yvG6NwZ9mTsURe5pIUkJc1P1NNkX+L0EYgVNRB6fj
WuQCXncFLR6hqGNcv6APbxF2SPQqQC4oocQeUgrQiBDta/0zgPIrQmGe1ZlK4PmQ
gq5WTkDXvOiN1n+DFj3hCykuzSVOmxbfRG3HJvCBk83wO89S7yHiCiyazLSuWn7t
T1i+i/imItW9tXUr9C+kdL/NlRpkXzEqfVHdFf6N3WKsdlXIIgW7PaU0bnoK7zKT
V3mzpPUMLyE8xRVzt9H/ZHf7bcclgDYWIC+iNskrtlexLbKnRQsRfnESaJ9j0zX4
JBkEpDvycdJMISl64rsTTMU+Hv7ZzsfY0hTNALnWhLd8AUhWvZD8/12NNiE8UhrO
3e+9zhrw3MAUB4fcdnd56ClqBIvLw35eUeAIpkvrbnROQme+YneSU6Q+yfUudgcv
AMG5qaZoFSfvlkYyPT9KNBMVw8zd9HE20oRDxitKt6OG6MXhpmjy0XJVQaou9OSA
F1XdToADInHsWOeoTilx04YKOOhvHP46TWX+HjZr5Y3///qF7TtwNShastTIyjLY
fuPSqnzEeWigPpUX2l5EW7cNcCdqljbYOvOy7/9m4dwgKnT1rZdjTHadQd/sUopz
8qgvYqrHp28XWO7q5rAVm3N8XW0Aj0xI+6ZhM3rc7dsnoHR3wxAiZgbT8h0I0Iwl
kiM0PjXlgwZSYe+SwZU6ax6ncGUjpp2pYR8zu/2ikEpqyAHU47UrjGQsbTAunioq
vPBxwCBJLxu0yJs85JrWjonCBr7wSx/aF1hJNkrqREQpetvTeOU/hWFK3+RfSf8d
V+m++XyOrUxzlpzVq4B4sMQKDvdng2PGVwrNNUSK33vE9C9W+qWOKKWjy+7Menbl
2s6aNLvyV3mSJkW6ShORvwDWSE11qfq6PQk3+e1KJhuwQkYSfAX/nwPIneUGSVF5
whHgSacN02eG2T6xP/5YlMAEDH3XWPzeKGwlJwtvm9bAvdJWWrJdXPoPHcYf/mjj
oFKzRm6270Ixqp2qHhZgetlhtb0Kjk6Olo0r20sND2V9sSSHv5H13o79vXa16gGR
V3ZeGJgk9HMHeO+iaMZfxgmCpDUY9RqjuxLlHQdxD/Ra1thpJObxkpNfVUdaPvCB
mkBn1ahK4U1uNuMmPAxK1gtOh464XbsyeGCn2mOT1+6MnaY5kRpcWBAzuXOArpqa
Qi8JIPeDhneCblQ5ovgLJbDHuvpkNqwsVa0Gw0O8YR+Jt9GzEWoqD5Q/J9KCRM1S
jrBy2xEmWeWcqzLHZDg5LSUOLyYBmP6qaTPET0oKhGr4SXA0OMj50wHEk3dMgOIW
WqxiY3gC7GLJ5mFc4bZL+PabXtCTtXWtDZGWh+Th+0o3yg6VJz72Inu559d2N5E6
WVS34SOyGMLv0XZOvL+SAvFqubH67b13nj2lXzHgrQvR9cZmauKJEdCx0Au3Y9da
xFsKSE7PNmvzXE9LxwifuwAZzduzn3i6TrBArxKF4LWxHC4wf4MxjT2NpQ9sf1JQ
ALbFFSAZkSI2xFjeuWWku5ds1aOkhIs8A5gEPFilCNK19T8CEq3nfV0ItMv36+6X
zYC2A3/re3V8G7cQoBiEeuzXOm0BQbM3Jpw+ffxFOvtMSaxJnzvdUPxgOmfuoyAN
Qfd2Z5aao08sVl/HT05Vxuibs8cw//cli/tLdnQEnE7KVC4eTsvsjSq1f5qora2u
Pf3UYMcU3JFRaYC1m9EOOvUV+ZqRmKoC0j8JL5JUgGTqHfpMZve8FNay5Ie7tXTR
nzyYQAQVJZk4y/7ZrOwXjBUoV3QGwKXKmWWJ8Z+7zlpMX0ktT6sQKBMWxe1VRrWJ
lf3we0MwO8z6B2bgFvemVIEyM8RosT7TUtI76U9rTQmQ5aTuCSuJijc+71xnLrsY
NsjhK7LuUDHFFltPi7GEHaGyvuAfEqL6+id4wsASwXWfA5f8/7bIfnWtTuJe8weO
jKW8oSfGhBdOacnl8tiTBjXROsN5sc4d19MxgMjCbJoDQmq5TSyQLQxxYsbe8IH0
xPkVE0o106f1PeEK+pWUpw0sFAHe0S/G1v/des5eurrEUgABpAU0QcKHdjMczPuc
vvYShQjLe++E422q5uq2XC/WHpJPZiW2jvEpvyyhFX4dM0hYHopimS37mNsdtGfE
l9OMUBB9BWXDCqtMhnu3ImnZ3l29NdHowWfTeHSQ6Pzr+J/lfk+JvSYKDWVZZ7IB
f8UVWrdRGNHo3Qr3Mu29hj6++s4sqWLSutkW0KuHl5Ml0yJRdRdT9xjlcVSCsfVx
h196i/SMs7C3T6M9BkM13wnEH7rge8u7527o7S1m+e3dNTNj5v287MCt6z8SZYBl
T0GyD9W0OA0YO5ieX/t+n0Nm3uE/tCBk7M9W9kaG5FOHPbMLocfu1VI7hdE+Csv7
sz7lR4/X+7f+77MR4pmvisoMcuVkpEEl8EVplqLtNu0Wc9LWxvoSmMIA8zQWPfzc
6Jn8IK2tVMF/0rgT+HDPvqqUnq1emPLkwr59GOmi1fEwr0efxDebL7u6iFqkUxr2
ftJNq+CnyG34t4n6+IpWEYtZKkjfQhLT4N0432aOEU1RmyG+k4tY2vfVlexR5AR/
U315iVZU1tVGRYtz24X1fB/N3XI2KGqiMbUPOeHn9eWYuoTZ6Pc/MIfWordqrWim
TflINWrhd1oseK2Wo06M4SSCJ9M5qKg9kTzqI9RsqYW4Xv4HxjrY1zE8c0tFb7Gs
fEJSshHAfgBbnjchsrckH1GIQpAP3ryi6W333LSzyyvjbgS0rHtPELdCfsUpS3Z6
5qLE1ezJlZxncD06w26AfPIGS46A8BBR8QEaO0ukCfm8uRVh1dyypCwl1JHMLIoX
g4S+Aw7ob65y/7xiHWZVE5DA1H0ATWTEwwZurwTch422/XgJU31E/iZ3kMvE/D3Y
w4ihSONrITNKZFFa3VRcI2cmpstMiEMGSJyYXj3A25ZZAfg3mgZohpX88J0il0X0
VVOGCAxy/+67K+VXP2Ss+9atFRZx/z1qw5g/7bc6y+aEyLhEU7RR0T8Iri90acOJ
HVmA3VFq10PLS27hml7PzzrJNdne9N7/vc+KN/vPkY3BGmjIv8F8CEG6mEuh1XGe
Yl7RjXviczTHJeOCknfxN6a3fdVRPFZrkt8NaxAkm5eqqIoVOSZJ0NmEwL3eVxlm
qzDjbA4C71EU1iZ+fL6AEKc8X0pHyKQPzkcm43BFpkIJ2TuUai7L4ihI5XrAwSug
Vmmx+Ga6StaUJb+cfuInWPYRKqS1K5bC0aCdRGIctOEx6U8WNItyxqPyacHKFn7v
YwPijqH6Hwzsf8vvP1mpqBtvrxE6bnhDE2NyHE0Y7BHclIeqY9dR6xiy2bLeOeIr
3bfkXsiYwRSsCUdTrjpTEOWTyV9yDqrTM/QnB2ElYloNNodeZIbFEVT0pMAo6xMe
WffdvXnXwPzyCBJUUuXNcURBJXpDJxNVjvjKX0v9RvBqlaT4wgaem3IoxR+tTV9w
QN49QrCUSBYekolUw89ILOJiZS7I9VeHObma7xmOxK2PCz4+xOU9f7Nj2pKWdbpS
8tEupq6HwKaMWo/tXkFu4PJl29CvUk3MtSc4AAKmMswikpMDkrnbgZb02b/Gp1Zh
+RhOY97KX2KBAaTblLpbRNp2ctG83LUkFdEieAC5giwtq+Pt5H5GYW4jiKYJSlX5
xPc118UKntZChUTOKCfTiRGBgSAp5WVX6C/xmiJe0u7PXrDpWQMlwAeuQbbDbsj8
XZpct3QXbltxJ6oAsW8W30lQDcBdgtqnWYeW0oRP4lxBtoTe3Xyt1KNyOWk2ASWX
gBb+A0QdfYKJ+HfJ/FANEbQwn8TfJ7xjY7z2Lln4wAchx+Nm92kI5rMpaEkoj1Bq
OGtB/d1VbUg7YAElP6MsMMTKYiUXTOk1Ru5vLH/yDPzTtRPUkvO4LqWfW6AlKLtW
3go971ZTrRry+jJj3+/nqOi4TLSi3YibgGgCFxLLrpeCavhLWuYrtjFVMlIzd+Uo
6vAK303+Y1SfDhXI1CRvCufe1UgScZWGJ/hZNpu+HwbV+W9JhOSc5MFfB2efYWM8
fZ2XHOeMJZ7gcb8oi/jmk7/SnZcyDZrnl40X9lfgpFX9HOfmolnqB5Y5B5iZbBX8
VIIqET8wnH9HgZF71JUmyy3bG9swH7u66lNF9b60A2FzFtAn5zwME09GpJSgaACi
vJ5z+NNxpjNslNnARLSPaligbIvUg6aWbyjD2AAvfotyWxt4wTfaZUwWtofLjo4v
AWyLXMz1Q0oeOARRgXE/QrniKK7u1AX1XFNQBeyW67UoAys4inI6AneEeIcmTEfs
yTpZ080TQdCyzfZdMjlLLb5LfXanKGFVrJ4wzg6WGHhlL5khvfdvc7UIK7QMNqCP
uvv9BNdSEB8/8CrO19xcTrudM/RCJwcGyCLnRgM4p//XVjKRZyprspLHBvWkJibc
WF405/wUhiFDrTZk+tWMf8v2e13CGBzFkXaF1j+EIzbgzID6tDV7FRimQby03HbP
W1aF/TYISxpAJfrdJlorpRh3KC6TQZwTR7kpXKwQFOt09aYVTd+U7NuMTDo8dvEe
gk2jmCWryAKA9IbZM6ocNi4PkPnoClEHGzOjaI4Da+NatTLkdNya/X0JKokriL+X
gT5CE/cyuxcA9pxYdcpgcig3U3JzwW9X5tW3D1B3wC2akV5cmWA8rQybZkyITz5U
gxg5NFIFB12fr7fTG9mLW6bqWojLjQm2k+xWUp+ouG8l+dMpVuatm8T2repgC7Zr
OmfTejZdphDvHmC60o451d99ADHOAbHErmuyiO+gME5jhji1xhdiNnA0P7DiLcS8
Y7bInHAtnBmz7JNCHkQdt8mwVBynI9LOa2+BaMlYhvgEBfUXy5Nj1E0Pg6M6Sk+r
EQ4K1icTxx/U1+/mHmluDcGS+3Y2kDGyt51v3gf3ikxMGU1YWETXgODA/Gj+wLI+
+FaBCl7/x82SfdafDQ4JjTkcl33J/mQn348PA7CGRIJ/LxrnXyEsJUXb/2kCm98i
jbWLQfMJZN1Z9UuUarV7ZXSs3+MGiGPUJaSwPIO6GfblOMhO/0CA1BAQdFJoDfdI
qL/tg8/amyFtwkd/BRSBGscrTxwfnvPj52dQ2UYlJq7PflUHoj/qkpLfY1sP5UTg
6nHiY/I/EcIQ441fYaEWFsTiP8T1KHdfyOq3iYdfin+NXRW9XPxswDjb+NVZUNFU
CmUd7PLd/yaHgPyH+0W90W2VoNWGXiFlLk3Wfy5InKJ+u8pj2xjkLWlHKyoOmsYi
YEJfld5U8y9r4AhJsTsh0Lup1kvWwmChJrXxuVideI1ECfSp8UrSWFFCaNsPVvIz
0naQ+9krzUBHyo9p/vF2Q2PaGvb1MpS3gxtL/Y4xu3EuqHDVxOzAYC3MG1AVDV2J
G8dHrRMDVphnkWD3JCCNf4QYSRBXOoKyEDNuXgzSRcHgww4yy2yY46nxHoI5L+Kc
cxt5uwrqMc/e2PMSqOKwLapjdFUw+e9bNLBY+q5tofD1YhEYQi+45DtguQTxY0b8
2iz9ls32Og6rgY11yuHPyDDiPULsdSqguHXggIrDYHQekXyGbX3nLH8SDLKNoRIT
yDVq/5ZUyZiC9uMtydwXSSFMDh7PQfiveGCh++E9DApbGDQbMDH6VdG48PRV9NGw
n589wKs4KAmaHnBQLBTSZjDlHYiHVsvfc2oXxPIKa4LuxjDbS2FSgMaCkwxJP/5B
4wOZjc4h++3jTnhz/pr16PTXGnPxIKtokHuaj/lNZYGujC1KEccVID3oAkSeqzj5
QECcyAO3GmBgfxrz4zXP7+4zBrxe2sbKj1MGdOvPrYDIhSPE1iZu6jSmsZ9c8+aV
1Cuo1f0iz1LIfLzbDDk2fcyIGxkGJESvfkc1nOrECaNCk9UTBZ2sIsf1AhmaFc9a
iPsOeQiMBCwIxgZbw9T1VWHyrfRl/8ba+K7u2ss0lqxPhvpOKQwAZhssepkYpqLp
uJqXeXBPWzWwR0Nr2MWZOYrMiJjEyTdpt6MH2ODC8hBZndV0FGXEiUREz9x7NhTm
ZSx9lRy6k5F7RdDYI4XEnBVFdCHvI12R8ib5OWflim139AdJ1pEULx3oUhvgst/a
MimYfTcHfRhWMSQofFJzu6mECIlRgy2RqOHqSaREGHw/qtsJjvSxRqPid7ruUeVE
dg1h+WI6AO31c7z/uyO29j20fv2xSbdCZeLRYwhUu4Gg0Svw6EETny4VhrXaIuyX
1B6h0mRNjrfgZO7erPBN6+3z2BYEr/nYwk/QcTP7trsM8Ol9rw+wZTT3B/eI4CUN
AEAtWp+7bSLO5Tfha+/kXjoboBr58jXN4RIhbXBJ4v3enre7ZiYYvzk1u7LlA4Nn
lvbd8vVgihcqED1zZkacjOW5Una58isvqwjYB30es4SPtNS14wtfyMpoVYaVP1Sy
W/+tOgtvIJkMxyzaJd6LVoC87xai+lBj7nHdlFhZfKmO+KZ5irMznBrqSLrSyf1J
aWde24LoYzJeHGvmazcUZFTG+fhCMV5biNWw3301IQeKK+7is/cO685QcScG3zMt
3O0j1lSZyAa3cHbxnD/C2V54CjKxjaa8JLzCjLM0KjeVuLRCf2BJkdMT5DA3oUx7
GcpyaTabDGAGp7UETdOre0GXwxKDK7QP89bDtBtKGd30JzQwjYJsXm+osMKN2llB
lF8w42DOQsmoDM2odGxq3eF8Y4de1aVlR8lU/OQ7TK87ZDmnHZnhnP6Ln9A9F7um
SO9T9pCHlOR8Xk8168MWsmSRhSixOU7kInUPW2nsWxfd4F44lI3u6gZK6sLxdKtz
DWBXq0Yvgc02T2xIxVI0AmS+JaQj9pUOXhIp0INlxrkR5swwd0OZiY3q6Q8EdyVP
6MfV/Qo5hCkxO017NcpCCpeLqZEA2PIk8zRRYXY7d9OUsAS4VjqWRbH1WTaJz625
75O6HAKus6aryWUWcdRthHu1UIwjxKO7gI4n7pVPLUIKBAZwYYFED0OR4QAmDhZR
9jBVsD33bRMQj9prukkK1dRkaMUH3R4uRxpJwiuq1eQEYsInyWIZOXoziAMx3eQP
ASGm9CIf6BGJAk7mnqmagVfbsTXpd2xqiBnLCFt4IALFK1RmPZMCLbInhJX4zEvC
dRl9fnsbokgAB36Hk5b4mHcTmXeQKbPJsQtyDlDqjV/6KaE8AUWKhBnnxCC3JrhO
ifI48gk6yEuVweaWQiphzDGGJUcPeS/MpBf78J/aLrBAyWov7KQfg6AlrEBYWwlL
WtkZ7MXIwdSQOkvUlhpOCCJJ8YMMkqqWfuZNGiLjn3qdvOVuRxUKglw1/lCN8KQq
g25NtCkSn2wY7ssiVjt9MBsTTQuOcos80+xWklXSsTkQl3GfxAddhzlM3n0Rg7oA
3cuYDHd25tAG5VRi94WdVLo8bDlGVuDj5RQn3NzEw2Z0mgTz9Jjw9WS/aqaH3CvG
b51m+SLcWivMR9U1Ce4CKdW/avkFDFzixSi9wWhS6TVZJ6PA9VpDP5Q+psg3I6EE
MJBsgJRwhXhjADWUlE1P02NUnVoNdV2oeUNC/5mHuJLhVf1+6YtvVaov7xJJvc31
iRr9PNWKhDT93Se8cu+2MJ/3MybbzazbvvR6ULnjEFvxsE2QOoJ1UFLLCCV8+Khr
Jf4CoQz57OyDXHZzxs2Zf8FNWo1b8Ej3a8O9zrhap/eJKQPWUXB3PMYWx/ZkBPZ6
sQXDI5F+orxpGe7pLsmi2Gi5epL3+GmUXKrzb6gDprhEAc8HSwajphTJifgWB670
+eZX4BTGz113dkoZd0gNWck7Kn/imfcKM+LWuJ2CjD62tq1V/VfO5k9xFaBnqbmG
65xyInk59pVdtA2vW+75iKRSJw4YQAuxSi1b5LoCqZ8MnVx5YjtjAWJOevnF59Sb
Hli76MfW2tnFbib0KgZaJi0cE3sOfXvBZDBokCgFaR8s4KpWSYYWLtnKVP3lXgop
yBd0zrxiYe9DnGcKDXDCK6+vnmzHtEoC/Tj/yxr/bCRwb/sE9cibowANiENfcER6
NM6VO7PwsVsI0IrlbcEeOvTeBGlW69YDn/JHtMgpcPCc9THuh54Fao3g8iFQ8wFR
15KXVQu/4/h3rce+fqyOo5PfrMmBPDL4pYhmjWBI6NdE8pD4sSM07x3WFBmPRxOV
OgyXV7fvbo0A7RTkupKZMLdeOoZHBmn2EP+XBpta9U1zUsbCzsdUYF+Z0vpw5CWn
NeyjVkveUliyq0QDXAj23dsjU5xE2zRr2IAl3m0A1BI2rTtO6G6pYPZ1npL6Vs5T
NKwSelFGltAg//lWOq4kaMfagaLorBXDJug9AqDpMpGqpTnVP290gnGDMfgid2K6
VNAQ9VLs6UxQdQSeeFfWXVxFgehL4gY+iUT4a4r76363f9TUnS2tCfbAUXkHilV4
69Nn/jpp9ELDLVeGp4S7KGcVccEHcEZ5CW9e78PpzBIsznX9QiSoeJn8Uag9udR0
QlIstzcVJao36jMMDFqDmzj/GfnwBeeBKYZZRf8gTuOdkQ8zgyyPzXRDiqk3Ve+7
mwDSiQTDEifzmbiwDClgiFf4LUECEz8BP7knY0ULAoi9UvSLUCdInhpSE8Gurz0R
i27Z6VPKFMsCaKbG8De2w8JW3QVdNA5XiNjpG5Ags2eTDsRf6szZINLR+avu2Nkh
18MWu65yHblKLOJBnUIK1UN3sRpYlEvFq7gVBxJLvVGFYXsOyl23scUK49A/mAeK
C8ICs29tfwhs7F3/1bR2TyS/4+U3Rkzkf5D84fa0Rkj87dz0HWcplw6y+eYwvt52
FNSZPO9ft3Uh+cC9rp0ShGUfv960vocBbYU+U0ODHWgkM9nkJIpX8rWq/CeP+Qdv
GabNAbuuFIxJH1gkojJAG/3R9LnI4D7c90FkC3if49ad3wZu3w8BORcxGJs4sDKA
ZdIhm0JUaSULdhOpbkQCc0D3rTa8ymuVCrJLeRCQ0KXDJuY0QNAkpRizv5HjQmsB
6h0qwGMguO0pMavDkFMsqm6dIyzILoad2LKLiro3uOhmDAvIp1pRvTBK3+jNWsQT
uMW8ChnmsjM5IxKlg9A2RM8pjjycktMcyJF+WjUW3rGjrKBdSym+59G7ke6PUt6o
kBbV5vMmyMz+Zbx9Kz6BvLOWc3SpGUzcAb4feew1AaumeJXdahV/ZHaTy+Kw0lss
7bLOPcnF3rqCSgcs7aRCLon6DUabjD1ss+Iyn+VXKgsgNH+gLpluKAv+dwrl7Pxv
2HXD6+JcKfWXSbNR2l/9DOcVCKoCxavAjFS6axMcDj/bgU+T+HF5nqL3WaKZut+I
d0NyiwEva0kDgmuLk4k5khoKU00th/czHwLl90dnh51iYED/YOolReV+zKTVj+pf
xI/3cxOcx2aTXzk7dA9xJD4YGRQnjZRHhSwksnf2Wru+fwFyqutbKHnDgHoD1Abs
L7V9O72NqoshrpJbK49cT6Njj3B2gB127OmRqs+tSa4pDg/LQ4f7zDtthTKJg3kt
iLlRmiDz09zkQhRgyPPiKqqqo4SYjEeb/ucaZMu74cWH4fo6cQQN74ZTT+LTqjTN
YyYB1VPqQbZVpJpWsR89PWin/0q10UsjO8FCLwQeVY09US2xQemQsNF7p6MjD1Mt
N2BDFNuGaP6qqmvNg0mkWnFhNZ9N9UdxO3QP6Tx2bQVZWFae9J2ugU2ouh8gf/Pe
wZwwG5DhxQ2zXV/oIkhA4A1pMem/xxHvJjY/FZtzgRxsmyO/+f+uFbfUVf9o2ZAn
aBgRmvAO2JpPiiySZaPf+Jk1nK0YG7ypfTzoypD+VqC+EuNHMriT95bcxNQdYzg+
jlRyJ0xrSiv9BUyRvRsW3gRd8e6yFc2r1T6/NnxQfsjHPrui7eDfbBUZtDR7xews
IpNV4do4nnN/jVDiu3Y0Z8dpGiNnTKhfm7vGcE8GZreKbpZsmVGFLXfEZK6f73wZ
krQatioBvvalmoyHMy0eQTAkuC3IXAhkbsBut7BsASjWUHvbDCjga3KPytfOaL36
TWBlhsoyT5OW16omhO7MTR4pwVhY8TpUI44KJEQSUnatvvxm4sE8S1ERuDjBcSXd
/wDQH6tvxqol1eUSqY1EKQR4dNnZORylXFIz4clCWarJw61dej+RNc2PrN9qCOPz
Si2eXNKLol5ris/0KpnKS2f0npiqtLxMJlikCZkmBJGsJ/Abn+pl1YN0ZY9uzumu
uHJs3ydXaq1cYkHXS6adCBt7Wo1Uo8YfIGO9YPSUsPprYApAC7qAOsX7HaKgaAHA
yV4wv7aesa8yx3N8OoLTXjsZe8lypPLudlYW5hFgfieJN5+BPOi9iux/vDUWwqto
1aFhl+gdzk+mvRwEtn6Y7UIr8k01wrJaGzRJC4ayfYIBLdwnVOi+pXC2SfH+3k3P
+JIIRlwnzbWHin8qiYRTBsItCf2r9KXv2bxhDvgaUaWd79FKx1WxmiWb2E6itFr+
B/dRmhjxxko73y9AOD6u3YPWpBASHigSJoz7HqnMdKpriMvhP1CKflYv/UJD9HoD
VAGQvmEkHSLS3aArq2QETmyRfbmO3MtsBibckCc0Kc5vZdvFrzXfuakePQ0y5tGQ
sWLZ4QKF67y7cpHT+xc3GGay2nh/UDBSXi59uHqbagnjQ02zPHsDrD/9yyLm/0ll
o1fidLKxu8IUt+sfIqEpitLqhSVc2Udq0igVuA7h8rSBijqKkE8izK3oHMzQBGQw
IOgbsGS6zQ8886QBknynMbDjVUt8/BJNcImcS/6FUvcooOJlbwZDJVe1QMVeUx2M
cy36Mc54EzvxvrBeIEbk/AT2e4G8f5d7l6r/TZLox0+p1AObgD698M5RYmIUnfoG
0S2ze0z+OBe/6SvTHDs+Jft9W18pCaaw6aHeRkzx1Dk/CtIzOL7HyMiYqhBBaksm
vCrbrUQ+N0AfLsUM2CSCx3PcqzZkGyLdAljV/iLS7gx/pKKXrxx4nADYw25GuVFQ
3nx6ySagQcyWwDOIdazGtXyCZC+cFnLqus7xROCRthJXX/CVLQr292Hn1b4Z8kIS
3kVB0k0lrseASK5aQyLhw9n63lp+M3LwTWQfGEx89axjzDbqiW2lkPQsFqGj+ZNc
EdFOVzqwYXDBFbLQVmmV5PUmPasg26XTQT7u76TS1Np17JtTJ3V88gmy00Plz5AJ
UXtcWis1LBuj8GjijjJf8n/sAdObmDSUdonZv4Vgnm7hWRdskXFa9kIh9x3/kTds
YzY1OGpKQqv7VPJNgKek+Cu7+79bnqmmIVYHbBRQQjVvn0uOewpPFUFTKNAcpZnB
KGNffuBGyUm1TNcKI92dLSZqQo4/WstIxZkI8qdqe6jPZLj2KORxbIVoRloAMPgP
q1gEa7Z71CwwgBMo3KUCSH6qX6EMbvDUIu7ZnEZ+CJLfMVLwl4uY382H4A+SK1l/
HD/kLnnW6jFoyRSl1k/8nFIWcRE4FcjGctACg1KbH3hj2tiCsCcxqkF1z+6BvsAz
qa/ZSeAP40fonTGVf35ZwGr8TLTxJRVsnViD9547bxziCYk07c564W0J6Pt+/+Fm
19iuy5jvf+k+XeveZMPMBTLmIMLBJp+F53XItOc6nfvKF0Xz6OI2d76CxRQHm26V
FRy7tB+mpc1Bmwsu65HCEr2OSa1bspyu/Ru9HNo018EUb1LN8j764cMcBA0iQH9p
nqLDHRwkP0AW5BKNPHYEUck9dom8mnBs7KdjX2kBZbyRoCCQeruaZChoqOCjmXhh
iNLEBWdDY/ZOb6sLjyb1NM+EiBb7FVK2bzMfaQOXijei2IQVtTgzlLaC9zNRMO7z
TtE4/YXilIq8h4PFjMr+2Qjip/6DPAm82Mi32MeENzhf36VzrP9WZ1yaO8Cm6e8x
lXFynTow7jYtW7MyITnXkIY+WXCLn78cEHdZQfVmTbkM73riYySsLlsVabdji8aE
1lqEf3BsJciMpww3cvagHLfwJgcvk5DHdfEq/qZhh3iD/hTy8Q5xrj78ulh+31F5
VjjXJQNYrPsnEPq7EOdSR9qOC3M8sIgJOUlu7SZMlOv1h/9lSB/3mcb1wvQj4SOt
HKwx1b/KEL4h+o0cz1uap2piyRITGz/Nh4Nml8O+6/ySeEdJi6sEdfKo7fEolizt
nz4KjOz9qyqrjVf2Pp9ZCPex40k4dFUHKKBpM5NGqLA7WIGgVKjipdP8z3GfmHcJ
mZY9mmHdFlSKeLkMmMNZQUqr9bTsD0JXqS+/6fVk2xvs0kQWgtSKxAHnYWqHRGJA
tUpp9P4lrwY6CFKzhf/dqCaxSxRsa8kmlJTaeyEln21vAUsATIXNslbGZRgzzDXL
0gBgrsmcmO7XNqM3utHCA3uzWxHxhs/LjZmwa04uPtJ1jzXnyv/nawS3mdYYtjRW
kiTVp0j6SgFvCsa5NUsvr0UbvtCV1QTiA6Da+17VzuR4ihpvtHQ+uFuQzriK5jDs
t0l3TsY6mPoOJyG0bl8N/MOxMObw7au4RrWjm91JETUhmnigtKbqMqXmBXzsLyWV
eJ1zlDynMMyxSxve8fQegbZarh+h9PE5PvQsiE5szYeqAKSDxaMnZ/+BHAEZLfRn
encocLDITVOaBx/LeAjH5xZ30ecT+gBiqlW2izdAI2hrdGMllWmYMK1MAVeotOAR
ToFUzEs4gRAv/nUC8bjaspBE1agyeoLM2xRl0M2ehMaB9vrfQXpyiQaGczPLBFmK
zNN5wHZHptWTbvbj94U2EMj/lXF7a5ZzX9TZngPQQHTrv62NWB/EAJgCv3q5hZWa
TzNYHmjJZfeQO3LtlxRDdWefNdiJxs21Xx+GIxz2cZS2hLOKxWBOzdBqcL0yHeH/
N2W/IrnxRB+xC9N3XlrN2UAmXRcXrNv3Xn/7geXKbY8ui1quSzvwQ5Rz2Ouc8LfG
/3WpLwzlbpn3oKb/MkireATDqGeFnszKReMzbVWeNy//MYYSbeMBQcc9hAJalCRG
c6umxk7gZN7rYWmG96kqqbzJoKDtXa7kIztTZ3k03OUpIavbNAxeFjIl3RGtYlj8
+zWQWmN1xSwHizkbxaeXtVfPMoeQmK4vvAoHVmsykTze+p5l0QKbQ+8UF/VH5esT
2tnXeYY6T2UJIAnhXSoSOO79DanQdGPkM64p3waeVx9ouXsxBgBr48TegAurtRR1
CPTl+LuYBUEJAr0yy+CdEFtFrMZXskoleDrxMDpeE3d5pK6tFxDvw23PHZPtSkB7
6eACZFvUlud4v6Vf/W47kfCdqIVpsTqhpMzoscwlBr5Vq6+nJpZySCaN785SpTWD
QLUfWvSludMdIJAueqnzH1S6FtI25lWfgKiqkqVM/dSk8cXfc8teOivfOoTdhXPf
BRzsRSfUaW1gds/H/LPMWTj+lftZwNXvBhIaMopkPq7wBaNEyKAK2IcbRU3o2+LA
iRYJb85tYgZ4+gl0zP3FiPnRUBw4mRrDQKZw/Y3UhFLmDli6HOAc8x8Q2jkYjkKA
4CTVT+AJlOeLbjME1RTLMEBr8/FwzOWLYcxB5nIPwldgFf3EUBVFISVr133KC1Jt
viNjgkDDtbMLRFcIfQgWpuAdATzIr/3T+Fi2hlC4Fv/kBtv1dAr11ReySM12Zn5p
gw/mAT1jWi4ruF+S1LM9ecDsRQjE4dZcvNdIqnPrdHvPpMY125GyggDJ3I4ZD3VV
7xn8R5DIH454KKo4Fp8hjrua2o57GPC76tbF9wcfhRGjjEqaEmn+XSf/yr47EoXZ
IqU5PBS2+g4NX7c4RvkmuPkalhTmRLSv/RbMqkWX4KT+7NyE/gNsm1JbJ5Iw2cZP
W+wejc+XpkUt2OnqcOIDUBMuDsIYMLdLYOMhpVvJY5CWByP02oiJEu2ZCjqIs0e2
ZFqcjb6T9ZO+HyuXdcSKg6631jf+Ux+keNAW5g7euX9epRZBOqCmwCO0D8gR6ffI
Ytu5c194hFBtB6uniWV56oIjSI7jzTQlWQtpCNwU1wAHj0LP/RE2L5Mfb7Mq60BZ
MJ0wUXDERw5pVuZH4GPPYzhKLlSi6NocgFmiKMVBWhN766+o3WIETny2nB3yGESP
kwIKjX8LZbb97SkejdH/DxssbqmmHQZR4dbrpSsXvHkoP78MJjH17kj9eAgui6c9
Mp0S3XJc3elSN4JUdIKrjXKN5niku+kxkSN5fXfb+uQrjIW53jxCjctnjDlHvRUu
tzkSnom15NEDT/XK3uiclumf/6+WcwAvyqeiEsd/c820FT54000pNiv5zz77i+jY
WDnwssgs9ksaCllLeDYlzCnFhUYkX3QHFmIr3bhauU9L6OeJmW7SFULHTeNDKZpA
UDZHc8/5xTPIRAMQ3H8YLCO3qlbjgI9eJLfHkBpWnojzQeYjQRIaNMWjx2PF2O3U
kL2qAAJfUkZgcW5RJ/7GMIppG1iXEV5e3F/BkGcjpEXDo+F0e4fUxEjxZz/HNcgk
dKZ9romaAzKlnQ94Ds/Z8C+VTOV6VshoYPtbOTuw7TrudN0b3IAtHlg8R6oEbzRf
Fkv4qTE8G1yQK12s4e1AXhJlormtPZW5fyeAEh5W4ErLIvtr687himEDhtf3vluh
lQjDoJfjARQfD2lvWFTZrbnXRYt3Vv4TvJCvw+h0mnkypSoR9QZQJKTPkGvTNUs+
RW1eIS2YDsyDdAiQsypcoBL75PHkF0pLv+zT4sP/vRW1dM7wQpUR3jUaLPNl1lfQ
3GrgJU+5Y4huMVzH6ffYjdCkzT1LtrjjmVr1HlE/VYif2qQIv4eUt9ThH8wz2Qmy
cEG4hFzl5kgbqlzrbEPmboBVmOU9cjcGPNge/9jO1DaGZKNpMqpAhgWvlSn20xCy
mMiEhjTcO7RQrsGPdwipsi1Ab81QNKavcEw50+EAhSwoW9vHn0p5AK+F2c2AKSul
8dKo6jnDo72Wdw1KwE3rklkrNxv7MN+ZnvB6RBlFAgmNPnqnx3RxjgxmH9MKlR5s
81pZol9jSNjWxqDKOsYB6X8I+A2dZ/f3YwbEDD6bzf+DNHhBTZIwi7pZxOwjyoqW
z6AIxuMCtCnUVzyx1jK+crglVL4/0iVJDLbyeh6oiCEGf0W+ODTETRHPIHvQZAJi
a9Dy36Kl8xdb9mJaaR9YRaiCizKR3bCItgG3MwKHDccXh9qCItz4kIeWf6WrwgwG
V3uoDfhH7Iv5Co5nZwoFNHlUp04IoSYko5XUWdjzncOxWn5j9qS7a9K8x3cxqlsB
qS/gnO+3dfvBRJlgETBs4dKiijwbJo/NTZk+n/xW3m8J0DzS6d8Qj45KLmhWJklh
IrTiMbTEChg34ZQs5a42JFjBoLHnzx/aOu3ndh/PgmUf3tbmPpueT3vaPAEzbkcr
Vugq7afAaxRM6iYcauJ+5P11M3ygYos7iEhFM8GtaPDaHeoxymfeLXYAwFeglWpb
7PjDur9TaBIW3z3mHYSh72wup1r7iUYq4gp93cwoaI9+FmfkeJNdUtcPfM+oeVPi
h1KZ3ZB4UbH2R4BRn9YxxuV2gA+0SIl9NUTgi+Rk9Mt2Dv5ZrEBzqxpY+N7W0oQe
IfL8CCM4ZkKz00HaTSqeKxUOh55Dx+YVM9IVhZrCodqMIHDc9SMtjp3r8sfsB+YK
a5jAN8JfmTK8HawVA3q9dg4Qnj8UsC/QrXAqktSleiPMfMNpy7hYlIV1YpZhEZvx
KDfEBl4r/KthT3xRSwQL1h7Z7xgBv3ivWmuvpz33X5IKZVSXe8PirNNGRVa3sCBk
j09qpzUalqez+8oprwHequPfhb9z3nnfYp3qXYc2R82sfgQKXoMOV+IpJG5b8yhE
sqTyF8VIY1gykhyaqHCpMQf0ldGjo1MlSsVk1BTlnWDgba6GSboza1LE51ebmZ67
tHb+vXsg1VJXSvgM+e0ZrJ9YF0t9QGbcBjLAZua/MEcEo5jctuVoELxEarowdfqh
V47ZVZ8NqeNR1HhZTepLkuG/KSKE8COhUbJYhgWZg2FjWS5AwtGzIeRXsv1yZVXQ
V+h3cCimHHlNXSPr2vxSrC9Gm3B9D2Nq0JSJMB0r7Vi5Q99pjpLK5qGywS4Xkt2v
T7Z4x8aOVVJLqzEIWhXqGTMDsNdSWAjWtNOFny1BDYm0DN1v4xNQLgBeEkjNlpP3
gRD+s9fIPLVCQKnYdoP90d3EOuo2+POm2/GrAuYfgbCpji9cGfeyG/ivrIiaFFjo
LmT7mbllxn9uluB7NM2N4BEbka0iLg+D+osqLPi4BYUvfOcqs5wWvTp7geND7WgD
pTpwwrJpcLOerfLWNgaeNkVgTM0XBvyrYoXAwyJ4VOT4Yr6qPAiz+JxbLHRmZI3B
rryO+gRt45xw/O0jLloetqCUiWlws/SVYgi9OKFpvqJmxDYm8pHV+d10W9BAE+KJ
POOQk+uewjKltkgoyskfbjCyzkJLMTDTtak8Sh+mAA8uADrMqi/wx+z9XdxChsWr
7/bcf4soB4pibkxLUM02IEASJ51u6h7jHb5nezuplJKEFYFAhvBx9ZLwbRoHymBA
mdC/VFM8twUEC7wmgkorXtHzW+KU46CvMN6VrM7rl68ILn/JDNZISBfbCgMQTQko
jPjoUtq/Ma9thL4B8OxDnoD5FdZPHgcS80bCrJGl2u0WNbQtzFga6zXBcFog6gHP
SCnNJJue+veuaFNS5JQvN6a5csUqhQMBqz02J6K80WLlhvx6UVa4uiDqL/TJDARV
QSqv2uDWaV5ojkBM91O9NfwzuW67CU8WAKFSv6KZSWov9vC9WT7RpvvkzlU5cWCf
fdkzSntC90IrNdrBsOkaVWTSQVTxLVjTyWLk9Dwaj4lRxhxmfnwAD2LId98Qn5gC
fk0VyEYh4LJ2YAVbf5O57E/QWox5Pak37pIjV1dTjukzXvUZRHrWsRq+Il8bT4Ac
7yrpgBsWcBT6XDGZoS5w+6Yzio0PnpGox58WLYgpyPAsFVC6JSnApBwNn8XeW9G/
w1vQ6Z+AMMug452lDPEV5FoItcASdbA+MnnL+XLrqtkmeasmIRHJUrjnWrANc9Ic
YBD6ZuP7YDa6JWHgJuUhyRv0GYBoRzpzgd1GDfQQYZTqOyS8mPx/jLZLz8XDAfN5
xcwF+lGK/ac1t2/EqfqHk6ovYUcGhp1jP8Elodjz8W2bb0yQqLnipMD6eduB3fm7
zHJGnQgFfaHMHC580w0vaF7aqNSsRiVx0mHkKR1ZDhWAnqZCjh1lR/IifKC6Ed+c
ZPtZRd15CFpSHwb1FBA7YaXLUracyipj+5DMnCQJ521lx3ZBg+OA1WvkTFa7Xco6
Ilq86dZ8RKZqvG+JR7Gx61FuZKIquCNsW5gpkh/8+YOzJJN9VoZ/Kvugu9MgxEdM
3DGXbOpXv0sH6l4QLuwjZ/NkoJg1nU6K055u0owPZKskI9fPRaETDTnp+7lfbcOV
lPEEIgVg5HakK59L+Zct9xMfiiiBZOCS2SP38CyJ9YkP9zjOpi3k2E/81qd0Vw+t
uXeQqe/vHmv6UjCbLSEl6Ij1q2X2PpgZxHU5pvHq345znXGIfqGo+myFUAmgjKgo
lJ365D9/alLQ7E2AaWBwFhv9Jxk5lAt+naR3Wt61R08xNQ/t1UTj95qsdWnsUHmV
IsP7lKLSEZflB/zyfn2ZFu0QX2KnGO8iKsRfSiA02yofhs8/9OmCjkLhHD9iVc8+
0fK5RYgoxdnkPC0cYi9Ui5XOE3vTS9W25eO1suGpE4p4TbYMjAIIp4TxNZjZoEHa
1QwEZX4/cZkdK1TfQAnFkB8M56meHWAn5kf0mkLaOyMRbKq9Y+9hnwgEpxMsf3i/
adMG+JEPjzBFuUPkxDjd9ELNs8VlXsx/KkMfMRZcykC386A8NjpOIB5IkX8jfd6S
RLhB/KLH6oEowsCtCDGKG4vxrZBao7bDGc1Rl+IM5Dq9jtbRsuXV+NZa7PGzw8x7
5mc5VoGiWrl0EwQS/7/juJQJHEjMzgYWAlUxDD8XJC1q4yEvgKgBctEvh5RfjeO/
FdLsxRCFpryhWx8HPfAfaS8QY3xSycTS3kcE4lgV/RyrJJdbGaaf4x76owhN3i6h
oOoHIVvYLZS4aq3QWw3vK/E/1xRMbyzz959g9ZlicazRe0IwSpR/0izqfzHGB51M
ZMLgvii6IIYmNgpKsVsATtg5JKw9a/YjbPCYy1IbMtLpvcOkSBMb9vQVxUDG3XXR
fQMwR/pC/wOE5RBHKHhEdrYifC+YYAP6ukX9Hg1N7lsHyER9D5CYIRYdrVBHXhx2
oMPD548aJdQJEQJOAop6ubJX7Jmls9jUAjATDuw6sY5aSGLejw7HezpAAhb+7vu8
IpLydUujI9RYxMkk/uwkNfa13wd27ZyXFw5aIBwZwZj8rYw6ubgeofYFHSkj2n/f
KycCODA6+DaZMQfEqTEdrKeMAWHer+CO1wRP+jpXi473Hb1dpJGKUjG4eBSMV0oC
qXWSo4GAC90wJn2gi/ZTYex53oUXpSGx8ia5mhAA9jVmd3oUtjaycHboCO4RWPwC
CgG3m8wiVHWKkxgfjoCiwTrOFrfzmhGOS1I3CgjPWPLqMpX+dDMSJCNc8gi6L5XX
K6dzXktDZBnJ91xv617ccXJdw5gWG9WqdmBzApVbStinXgAmBgE7Fr32RKJMcCiR
+3LD9i0KL9Ia0haAbig4pRz2S1p6xiWIlnPy6j/l03he4DZSsv043Rgm76zQzuoi
XoFu8lzEjWz+Z5xUQgvwfTniRujmhrxDs8bxdo5GZT3kxSvxEYJS6LxIiWkgBLaM
l7rm26bVAyhn/r9S5nUjuwqC5NKsADmUf0NV7hZnvDU/BDtxytlMPw/ULMhLUcwE
85KEU/KxBqLaFwdNLblNO3Fi4nIpySkRkk27FTWKIqqHaJ8okO3vVFmdpmju5f3Z
HUVTozzeWtTQG8FzPdkx3gMhhEprnp84VhzBnagptsbUnETsB2gKjo140Y+pH9dD
TPnjTcr4/fMxz926fRicrQtXvvLSQyUOok/5j9ovoRHmzH81lt2U6iyikLHI0k26
4wI8DIrFH57qUvtLnvUKlwbtGAeQzZOhpj4jk+gtK7DrdptebNtVOqTkJBsRMbjy
ar9cl4DrZQLf1w9znsimMoHkLtkkwqTEnFi2VJ1jmYXOAcX/LJwWKYOOA+qCuZsS
oUWPNdg/Y8PD98mC61GVTFj0f+aRK+Bp7Iqld0KKG//FHZ3sCl2JYogS5tSEKxFY
K0QiKCWkgjOWmzOGH6d+Qb4PXJzJRHVZMIDKhv2FAJc59DBABNdsQxW+U1LlCbda
69kic00eHpcbz3swgKhLVmCIaxdPIAO6Wr3UG8RqNj8D8NzGhLN4N3AOJS7QOxJX
y/2qFBHXyRcnlmHCSrgwm8S8/VKbCUlGk60R3Q/3AtdgWetqyK6QMMKWcM94Qc2L
k/T3mfct19a2ma2TEEb3OxEVyp08uPDxV3OggY6DXY34ABHYIP9FBLARkzxKCHX+
4W1HUHuQICyf7mOy9neyLZgIpw23YnV4LLeKaTg2ADjj0eedzkbHeSRrPUh8dUN4
wXye7g3zeST3B6kU3cuDH8tJTg4JVnR7Qoeb/6rh+yOI01Xohnf/KEIPs20l/1fN
59FyicDDoDZHrv5ep0vRunPxuM40hKIXjdeE0yh3TiXHp0QHISPYSYC1zFPU/av+
nfhNV/CIpbaWmhTMAX55HUKaQrpyWnE9WkySDx29Q9lZj3eT83rbDLttc4EUClNS
mw5amY/2cs9Eullh/N+hiVDR1/N9lz7TNoJB5MkR6Cgm+r/zj8oj0tbbsZv/33C3
8AA4HAzI5nj7ZLaXrd1NMO6NsxdeV6g6MKIWl0vfkwyCMJnzxDsiPebTF6nTDXnR
lI7qB32iKustzeIUG9X7xoj49T36ZtUbMQzL8GzhhB37NaknsoMRlfmrVU+77fcq
VqU48AtKLKWWGjCzCLdyCC8yZuMGBgE6AgcBPCm8viwMSJ8Ns/w4YM+YAGCnz8LG
HpMLIFWvDRJQIHZJxJ2ia5IBvMUEY2+9xteAruRoxMH5dJdosNAg19MUgqNWR6er
2wTcX4BYqL043M6/nT1f6k1Zrzmq818Duk0xf1kxrhaB9T/xKdfSD+aS7kTTNrjk
6wJzS+ZNI1tyceFvWwGoz+9BaUwZioNG/Exfo/RaqeMjizlNzk+BypQUyPE/BEB+
XE3Yj7L6n7QwREZ6T7C6ib1mU/f5H0j06EWv/taPud4R6YQS37Hvw92upjiHf0TK
kyODR5XCbVgKxFdawncprOblR6dMIga56PPjAoPhkW8Y+6gNRxgXJuQlqUSIEfWX
1Rz7dvF/QLF/xj2PLi67Rn2tcczb/cSNXNYVLfXiaDtOVArU9/7bSebuCQ9tYZTe
Bt6qn8bYPAxfADQ/7Yg72BNfjoFZnnuVgTMJ/65vGqw0E89OA0C6zsYzLje+lK0P
/pac2An8zhOvFnKZhXV7VoFtIeFp6/fY+GtGKw2FJAYTmXZNsn6T6wU0X1syqyVk
mzNqVkFmGDi8jFezTzO3rRuWWTJ86PfdTfKrrZyMjWYreil8x4x3kpsH05DIH1tG
0JkHtUZsieSS9NBKVz0uIKHvfJ3Nbdab/jcFq8UxKc9Ng2aECbuiVD9Rw/cqXX2Y
pYm+k3O9FHwJgd1TWLiQan73Zy1eU1k4rQSjfh5DR8fe1gA8h5RoswQBcmTQNU5b
Ob2RBjjglZTK8Omz3LNCoBSRweIDAVTLWBY9vCOsfAxrBpZY/5IHGoGPgsuu9bL+
fa1bPTRX4ZMDINe/1nG9kpoSBxg0R2qUz8nVupsF93Tg9whzGkKUfNBZlADn2JzH
PS0oI+zRY7/MljtcXy9VT0JFGtVyOjbojV2nX0wSvBbBw1jQak6iwNZC2WUs4crA
MeDZV9OL9+ck4nbGmx72rGx7By52ZWggXRrt1vxQL0WGZrt3H/erJOSxcWf0UcEx
dBasBvpIbJKDkJf9Ke0vs1+NuJKYT/Q15ggy2npBz7KprzfcrS+V423EpSpynQue
coiGiri9RLx1KFqznykZS0SiNXRhokJ5XiAton35qu4/fGHmj7DIHTfaQ8qeNniy
aXXR5uh9GmIw7Iiemi5ui6S/MC9VFfiXYzUxOf/3A7Xn8pcdr/bR4GfuK7Iadhee
uSafMMAnhSqOTl8xdm+GlDRa+HSC+Pqbb3dzFfg5vWkHb6PhDyaRR/mDcoJxGDgT
MP3+X0gZZWg1apAA90b0qCNOzwim53hBpZp3ep48JSF63Sn97f5sEx4Lh+H808GL
mpdy3dPY+X5RbDkRsvOyxidHth9y3xFGEjPZL+Tf7+TqSFkh9d/4zUiDQ4i81gHX
PhjZpZZUG+mU9h200ADfER+qCh0ZlMgk2dFvMTucZfRPemYhXlVi/Xw7Fw2pb8lL
KmUPfDztLcY2NkfYUMHBKgGNuWqCgIRrIHkdExLiBeOyhnBI/5BWqdau468ROMVE
ftrlJT9DnHMnpYu/fGFksYxwJTz0+9H05AxnVfo5qnVW0WUUda4zrkYntNL2zhf5
aD/tOPH07u+IcTBCziu9q4bihrUsBtMCUWNSf0bCwB4IfCU3giWLN32qq6qmkrn3
W0h3szr+qcooYv4hP3WTSSzzkei3N/3t47O0Mwv3O8CkYsKTBU0ORZMdOiczM05a
EZMGmHXPfjjlqNcSsWaVTA7kFBP8w0NmRx94lNqhKyMtXnRY0cFr4Gb/x3Gev56y
6ckiP6lJrqfmT2UaCLsCu1GiwTlHsP9Tdfb9ncaBTlXigNNvNUh/WkMb0mdK5evb
/P3f45yb6H95uXzgKOWU7O1/XYpjTPjZG9vQUofQ0ep7jRCPMHc1W7v3O4MY2HcD
pyurSMLzpiMVr26sep8Esm9+FWcRyJm9gYDHljz9pANn3CmZ7IofvTuBM0UiJowg
ct4OHcHmUGXbiZY0LD3lyHM+WWdU6ilfxntVo+9v5lI/ENHfDWRr8nqfpVlfNv2P
/Y0QWC8JU0gLQgS6kcg8uMe28jzQGdAeijDjNN5pmzJJ28b7MdgJpv8qWH3fBEPi
egxgFzqwF7SJQdXP7f17N/fLyVV1CLz8VmFUrRRnxTgeNrWsnKYi8AbMr/n0mgMc
/NlHrhq1P+bHW0FN6L/WFEwgGQ3EE9yiqfJWLpadSQzkAXqp0+7izzZnCb8BeIpA
Va6ed6p++czIuR5Vr32f1Wx8c3bCzcZiJGcqb2pMgrW/H3m8o8ok+XFL7VTYATor
DrgqsqhaSzoh9l7+qRrPkEnDwIcN5ucK6e0Uy+O6D9Y4BmakVLfbomYJYTv0pkaY
qc7LtakGJ1M32oeRlizHLJZk1qAws4Js/BasrXh42BUfhJJWHAKiM8SpWYk7Ag7N
gFnV6P5LlwlZgdEW2pitrU2FGAzOUEXyNbdHftc9ZsLXwjjj2OS9jWi4r44NBhp7
0BhVj7U/KlLpxmfxLmd9gp+Glo23hFPlLnEdpJKDpSTrTuPPl5z8eG5FUJqszhyh
KTLtVJ0rtHj3OrDG5UGZ/cCVNRUtSk6H3K4/qb/WlOhYHKr6dU/UuhlbCU9TqBxE
p5lyDU0g1QziDFkfh290/Df3u9v7iH2wJQrmzNHI7cnzXvvtMfsKYnm1juwusY+U
Qx+hcx5e86k/Npy4UeGEBxSpolV4oaN2lIX4AzAQasPff6o+DfCvlQMk0TaijKKa
Ip/n9ySSzyaBxAFyPmefnyLhaG6LMlk3YQJWLNmPjXduUkQhq+9pyqJPe6YiXr2b
a7nCXvOO65/Sd4qmtidqr4BEc+Kp8f7Yeajq1kzxCp3TG7XQLr3voeAgmL8SmJDr
kc4zYI+2V+Q0foazCpNCqaDeoG05Xej92jREv4N+AKUL60lvcoEmvtnVzqOirBwe
qC0KDyFwUEFG1FvIMSW8vL3qVW06pvWHXoVH7Qo6l9yLYG0fTfW5Hg2qh3C70Bqe
WQkUlOMSP/EoCS4b7V4Wp7KtmxR0ibajws/093iM42eq0Q4pnK971vmoctGGKCPd
S+wHtNPF4PDEHckhneNAbr2WqneBQOKj/nCOJBZDKsXACfuECglEIP725X9wy2cd
X7demIklMxzNHPmrbnX8cSxJEwNj2QaZmEfE1sFGVneLuvtWOST7tE6Xv9LC9W/a
yNcfoJO+8CWx5XZiSafSwLxsi+fdDIyofSxupK5G5F9BLGFnH8KTbrLbtgFD4z6p
NXs3SK8rCs62L0vlL++naCJoWBovn9RCLfg7+Kl+4sV2AcYOUQ5pWVWKVL1xNYe4
tVSoC80B0l8HvNRv8MC3U4U3dCVKPRvIX3dw29um4DjFH74qr3ILdbaiUlWg6MJm
sbUg3Q+ijGWzU7ztF/x5FrVjHqv45aOfosIJ1tr5hqLY5h+BmiiJUfGpfLqVYQeW
YbSdBny9tHBdm4hy95m/BKw2UTtYrc2WXkjjmX7HlHmKHRU4huI5I+M1j/aNzE/+
sl/Xrnw1FOSa37982cUTHwB1rHS7AjGhZqwIJqt0yqnbMUUmOFW/ZkumPzR8CJQb
8gvtnxjuL74klLaIvNNuR3WuVszIvW5Z+9HpKjUP6R1VREX4sqA0Dam4e8tJht86
IJSO6HblpdDLl1JyTmGBWCWeiTcp7Zq3pj6oO2H8flTJ6EwHs44XaUGq8YPt41nX
igz7m8nEKj4GsDUBU7ItXs3KseHBWqX2B/ALs8sydHFA4IFYmd+TDr9yrzcM6RK+
uqkG768FfdUmG/YubjYoCDDFz60Nm3kMDH0B2DFAyDdedHlvULqgqh9DHsg1/0Dq
WKZsaumULQSQkEmcmVYdB+3Q5wnS5gr7QF7s0tDC27sv9Hg92Hbc8dlCEYREofNL
YT55tJLd542PduiVnrO7uC2MYdv6AOce1LtsOMDSXXNkfEBlezURTJNZfOW09AfI
OkqcyCE9gUXFxUWFytJiWS0jbKEUQgUXjvipY6H4BVNsw/w/GpasOi3PdHl77TqO
RfMMSA8FMl8b43SPMy+JwMjoNWUfMQdyb1A6AlZ7OIQEI2w6QkVvqBhxPv0ypRtj
X581oUBa0Wm7ABAPHyVZr9SSoctIri8hH4N3gdweoo+mzqumXh5+LMV9swtN58UA
4aPABq2dSWGjDpDaAPk/AJn7rVycZ2IYoN2n6Ub5hzkRn+moj24j5RMCMq/STL/B
66tSWyhbDUg0wTnEu8jeMustZ03NDZRCiVmrCdDdk1s4ulZExTOODtk9AMGMzti1
DIUHJHrfDt9u13pI4HEKp0xwysA5dWo+q6qAN9h6IFK09YVVFf89AEdhHOp305ww
RRi1wtb3xZQPyNovgmbWlIQE+uwvqhSkTiRt2FRx8Q2+eTtBXwnrdW/az35aXjEu
m0PGY1QtQ/NwIzz7L5eYLzmigMYyCFvTlCl2NXFJE5ECQZkq6flJEQMEDS1nOwaF
H33BCP9sullqKe/R+vA0GWQ8ywA1vLUtIlq9/2Hjmyd6kR09GUEx9ZCiB4c2OCp5
djPiLBJTdA2c3vlNMuzaMVkC6aJQnruZGwzfagiSmSVgZ1fftM/NEYeOgf4cIGWM
Sj6cBH8DZSsCFwfVvdgK//D5Pj03nL6KZeFKsHilRBqmpiSDD1hkZENj9TrL0wr6
HpM4YJLSunJZbOzSpHOYTDKCxtr8Q8+qKdJ4tHn/9KVN0neelZWWnT5U14wxpwPA
exLyEklyo3bEXeuo91UVpka4LTY6Xhxo5/H9IzJwaFG/LMorMChIFfiZrEGSXhLG
V5aPdY5arsmKUMUYO8c7QClWNkJzBIeWuGT0DQvX2gkbnmHHej3d9jZuA9uRA1ub
sA2fQPxWXUOzw3pymHR4hjrPa6dYdL+0QbjDDVaWw07AR1phCViMR9hZhtQN/CdJ
vnZScME9drkY++E6ojLxphmsQVbRyZCXlWwboHeHxMNhY9oXp6J1+dYdCi7FjHw3
EuoO54uhwfKv/fQU2CI3ATBWl/Chpzc2JeamGviKgb1xsn/wiRZdVbcNjLF7L9xp
Kv8B5YlIi3izcUaBoSklQJarIiZ7woTNyNJ86XWErgvP8Gvve5EHKpOl529Hz9Vy
CwTddS0yacZOwtI1SN6vmGcIfcjR1WqwI5/mBQ8IG3FOp/x5d2SWGxre96nIVbDx
W8EQWO+VKbgjoXthDa8K0yC8bDr0krsFX3AVA5nd8OEPPqefieJGWGGI2QUOt8r0
hUUt8jBvk5gmeZA4BtS9cCWyqBfCAoeaDlHtYoDe78sabzIAqG4U5MIKX7r0a3+D
B1uCTGpViMKgJ93sMMTak04K/NMPmgRiFBX8OJsIs8GNxk4aGoc39QRPSqyH1mUh
Pq6aASVCbEaRMhzC9zxytRcWPdqrsfbi7pw08i7lkw7EKi26CLcU1z4pHa3rKdoP
U84V0/blzHgqv8OJ9iSy+OMqZuMru7lJt0ImVPuzBZa64/Hhf60ep+Jg3QDajaEg
VinGn6iNb4ZPn7ax7xFwHRWgzVSlVcfs4V2HPvHB1hkbPqG+Dzd62Z2QZE6ON9YW
J2e7UnT7Lssg9pxQGRBCwpC0jDwn2uRR8qsy2Xq0NHHVvw6YEwHtPFbMoSsLy22E
zYcWvsC7oFYfyfIr24YUOP1ELftZbDIwYSixRT9D20CoG9YloMvw9PleQIkA0W3J
/dlJRuX7GuFrgzC+VCGAVlxK5HReGtQdip5290B04iVBYBFFw8tEo80gz+D/3iyB
dCz+68SxFwm/E1ssetQjoLClm5rWvUNwApOYVCXoKIyLa36/0CXcBmwJyuBRkjcR
pN5mBcl+U+rHthVkn2zmmX9a2B9/luFG6GumGxy03onZMno+oscr3Zi1G/aJCQn3
S/7WObF5njZ8wJj3Wmq7GKjsbsKrBme6cNcx2oUHdAcQoaXa5IgwJ4lGL1qAMloq
DQrN+kEZcnMwRJ/e+hE2YXo4JgH0nKbjAXNcwQN6mZe5EosE9Vd2HK0EYr4UTr7a
q/INJOA3O+LFabREz4Ht7Z6gJOOp677Gre1/PFrB3jnkga1RAkLNu1kGA0gP5/R+
KSoPDCnypRmpS7vfVN+s+RaUHUfw0iXibPhV/myQc/1w0/YOqnBIWnlGn5iOL3vz
KhocIBG75NLgjtUlb7dOtEP8gnhdMvE2uuHzA5/GdbcDeNn0AqLWdssrRiqEpHFe
01Vu2agCEw5Wcy81WTYVdjegRjppQ70iAca4m7c8sVeNg8HsoB2nUYknGkwWKWwW
dAOqNVbjrc+N2ybxWUqUTiVRhrHFBksIumxBmrTrXvte6gxlz4t2GKsiADGabG1j
NZ650jmKsM4zjOdZDTs1n4LkAvI6MAWRl8ku8/xTIO1fJqHDKsRPKTz9WmbQj0xW
uM++Lw3516Kvtz+Jd4cIaUdK1/zGl3gAiXMXkdeaVneru5bwP6j5mjABri+74KyD
S70W2hU91u3BnC1PZqGTmEyDPeqnDHiC+VfnaEoWDa2jItB+76/f9MoovhdRB7+N
HG+EtD2ZmLk/wfIMcvjPJKyUjWNsc5elmNLl2xTqWMjqsCZQhyiTZGp3qJamhFpY
W0iiAhjW4cdKxGc6Ma45NRarWendF8EG6M7urHw86GTnj6syss+xJIrVOd/OARpo
8Bo9kzT/FiOh95Tk00gpPjV4cfERUtY6oUxlM0Km3DLcAlvbiytnJDiw8VPdoFA1
hpyZsJ8WomTQRHgrfMUZVA8QfhKiDPwjO77ehgeA0/aKyF1vBlfGM57/qlH6yvbR
BIjhc2FY/pZHOe5bmt1Vzuz0ZczcICypI6KX2ZEHtrkVWm3NaUA6RPY33ObWBhLq
w6hEKSC0uXFpZebW7/LOGie0m8ZNM28ldBmIZIuiuFZE+HZ5eUE4y6djGFcfQ/WJ
vAzaqTX9mNkPVkCNQlWVTg0FZjqj5e5zfAvKWCcy4IOkwjTYypOrkdChvf+nEaip
jmupGesA9nzPeWxdCjBHQP53gUHNA88eW1IOIikpfXGG4pHc9Xs3VIpEknmx6+s7
9e6YYhR1UKLIJ52Iguhzgtzqi8YgeYQIqrdoaRFIj3Vc9cAvJTGid0C2tqT2OjY7
EyxkFMLr7gfB+1LpmA9B5mWp44orjccNjn2X/zLawlUj1yw5waSa2sKs6BvwOYXZ
xuOObElg2RL8DwiYYX5mgpLQFGNuVuD2SaUdaskxC3fzwfeJxmAmIUbyEaui6k3n
LUXS0pCg37Ywce9SVALAbw2qSqgcTJ82DihGET534lzBBHXEzKbBd7Y/bzoGqRvj
10da+yxeX3bT9HjnSeQXwrezP+xgcClIE5O/rfQiQhFBuAo8wk0yUxHcHpw+JQSl
DOHDplh07p5HHaxSUhbeeNWNICFjZs5ND4q+cBA1aKDDkOywEHeeJXfsCKLu07WE
n4lCdjqrbMFyPfMqPaE7lLk93+zueLAvBdZvMU/ztlxMqz7vTRkCRK/xr7dLL7Us
TYRunQoZzedeXpVOlPp/xFebN51/gI2/yGh3F2wFYnWYl4vWKwGnD1/Z8D7A9exx
fl9QiYh+tIcBPbEiCctoWTEekMlQyDxXmXlGCM3L5Dzqbpx9xecuW/y436caOe4Z
DgT4TYCDmXpm5ACcmg09dNYB4V5vZ/MTMO6JB22KqJkvn7zGsgi03hM3w7GlONmV
uHiZEYkKffg7LlYvr7dJ9Lzm3xllbax//GUMeJMxr7BNVXzKnt00r+r72d2b6pwK
xeWD4Rq21woyJ/jERGt3hNj5YJGccamtw2BlmmgzS/JUhBRP2JpRfk1Z/Qh0NUAU
KgL60k18ed175PZrVuaUUueehWuTPHWeJXwtksGRYZW0YpWWesBe5h3SRY5chNqH
LjbNQAKeHU///FICqRdy95aWANX1aXlDR4f0xRsDXissuFatOEjR5w3G3c99Wr/L
d/zwcO6hXYYHv8H0KzMWqo7YXiok4RK309k+M2K08b8VV/GD1xKVLstF35I2FfKa
da+3fThTp0DGOMeaK8JLDi73aifTNWJpOV8dNNDcvY4IkZyZgUmBEtD8eRY/BhIa
PNd0R2q0VE3SwC+MSX+e47dzOaxOroYzXTYcLzSdHqq03G55aEk1f+Jx6MpnS19B
NDQOPzFU4iaFzWlZ3f9NPtALX6V3ybPn2Gc2zsLoOWqhB1HLl0Khrl5CTYsBB/ta
MPzh/6lVe9fHzpMMNpM588otQpmVRoOy5wRCrH3XFE/M3bLT4cBlLTyQ7+16Z2/Q
G9TpXMVPZAJt/dEdjNQCBExr9NSdttA0hu17k68tisWGPA4JSxb+uUlroiCULgi3
iAu8YZVJGSmwlEdTZ3rPcLcMNvfiopYicAM96VDxK7LdUjr2qVkIOx3WEh41ZLSR
o01CWIG1OzN0P8OoJf69Pn6amO6fYIy+Q9bO5jyCAcIoKvObXoDAMMfpnzFz6aCN
xSU0UlkL5CUQif9XFCBljx2ctmxY3YlhhtSiofV3TEBH7vN4vgOxhvLn6pZptSaG
9RA5S7dHExPkGpTSfGBj1JNh0HXzyFgNQZ/sJg2Ocodsbs9HVJKsZ+8xiIWKsTxw
ThiyCl4OAtPHDv4wOtL3Z/f2TnfENsYZj6HBh27WyFD3m5mMauPxb3OxJOxC0zN7
B5079qgSi8UcSDXcbRDriNUiam2H3DR3R+BQ6y7NzNpRDplWU4Hkj6Bet8dXbNU9
MyKBN+VQ5Pg3yi5nFqlcfcgUZPvIQ4jnmMTU5X2pCN7rP9ue8CDqdntSrnboZSBF
bHeeA01DOUQnrSrrC5vgiXVkzG081874YLikmQ627BIPBBIqu0SFyAiaX53RxGPO
paoC1wP73OJDddIN0QxZMjMRpVvsh+HrcQdjWeYgQY68kto/7MSOpPqxuIGk59SU
UgD0sx2Vt6wuji+Lu3Hiu5ILmaVOc1vrzMe4NRMTj0c1c1PSHxZlhYBC1uzeDgc2
ioccO/7EMDrGVOvKpu19tJ1LleYOb7pr4NcgsS+tafoTe2dxcDZ4D6Ti+U7nmFbi
9t5MNh0+xb263bMwB64cmM6rFPW9ZNSY9aNfYI7AY6ElrP8XaUUt+P60flC3CSGJ
4p5ISNhJT7tBH0XCxE+3Zj1jV6Iwsht+d5X584fQQ6PB5fHPrkkw1/c5SAaOmxHt
vqFvCvxF1/2mvEM2asx1Cs6F5Q45jb48Oy8lnzSR/PIaRfjE941jIS0E2GumaQWE
czFVJVT9KAEWPE7Eb+biEvpAdeulZbwvAbwq2pfwBMpky0hmrd0Ih1J3wHBmBjpz
hGzZqlziHPD/78mnE1zomCd6T2KAvkGCigtggF3Tfl7h+744ph0HwvjqAEQKg8Ty
wLhSfKZiIVp0KsCYgtqtO8pXcGpTRa45/YXtHhErYiExDTyaJMkrRK/XyeCOrlne
qOtR9S0Z/nQGywR2GiFtCzeXgwfUvojAQvRreDPjwlza0j0i4MXxW4lQi7ic0EjL
M7m+cmHAN/N+rvjTjF8dzKhxFmcEZrkcotuJ/SItL+TiHH5jNgVS9niL5xO/I34t
0hjt0A9lBqp287kHvhOHm8/DPrzDYdznNNWENmln6YGh7O+K6JQIWnlrBivry+7F
hqXckctznZzwzTbpHmzAcv2MVogAe9hVoKISCAILCxCx8SFV7VUkHJduKo2hxJt3
J/XUeTtYBNpPWv95QhRg21dc7ux2BQv2HTXwfHIl/n4a27rxBrCfg1EzbTaqgmVu
95szXfnV1GD0aFd01CWEJmv5QpHde+sULGCs2WcK4cQl+Xipy4II9RhmMuMsQBDE
WjNzHlC3NnHIu47aXeQrF4htmrcTdTn+q1BsJN/Nb8FCbmrARKXHr2IZXwo26/f7
so+EP52+rD/4R/v01P1SptK9PLYFbTNLF0iez8gX+C8wbwvT3m3ep1elP99ecPdG
GroxiVGxGH+vkDVkF5iFojkFym9xSVLeqYEsiTM81iNQ0qjRkjbKd0sxT3hY3Hus
D35RSDaZMKS32Amr0mQJI+oH4E5Q8d6DEwvFGuHnMsNXpGH2jyVaeBN1R3mMhpoI
1DfI2+4/dNeG3L4wwiDpO9kRew+hNTmQM5qS1EEKYq8cyXZxIRVr1dSWGtUj1MAB
GvOU1Pmg6Igiu5nI/QcVuW48acgskdr/cj2poEx9ZG+uivsq64agW8q0mHN/alma
toyD3COAHV4S+dLqtR0rvG/h4HNBXgNFQJP68zwN8CKecvrDrsfeBJgMdd0FXZ5n
YuZwwy5nMZunYaOrGQT/OhqYRvZaAjPY0hkJVBXH6On351pV90ApkadvBl0AYz2Q
3cMGLGuGzVOMWDLi7nurNLoTdcaJKKyXnJjQI0i5gV1IuqkaQh8WKdNKWCg+6vE1
Ed8QX/geCENeiMI1Rx6Ra6Fd6xmLAAuUujU2UekOVlQIwx3QxdMNYXRYkBVk2fal
SkVB+0bfu9e8gZyIrZOXe6f67tKJYn8QpNySajDbmTKPDi8a4EwCNYpRWwB/+F4f
qHFzdjYe4e5JLTCuVh0zmL8GkKoICA1Napo4kEBrsSVAGJENOgTUnsoKRhEu3/Ip
xCa/D/GucNTX9uHpqqm2z/kbOBtWDjDr3LjSZI6FNrflhUjEfLKOuT41uLEcAHMO
iIE+zP+lJ/kBMbGvyK4YNfcnGxiC9J66iQVEtKTni89ADEtjxars9Zs/WoJKnS6s
y3H6UnEZMiE5H+hIpVc4+hm2UEy40bWgoRhwFRSy6lCbjy2Zur1+aIEb5oh1+dBB
FrDTsTGSamQRE0d+wRL9r+MPy9DuCp3MwiGvJekOi7AGHWrzmlEbW5Nm79CCUqx7
Stf+aaMN1PRbqMtpRkiG5hbEe0NLZQSy1N5Y8GpEpd6dhLSo9lW5BqvL24N6tZSI
nO4+xOt1wj0m5jZb6eOJnKgVZPOWleGPKpEYyHCUKHA0cxUNEuXZiFiZXZyp2ddH
w+ca26qpq9wivIkXEJe3mOIXSwqQ2Eg2mhjXDvq0l7ZA7IgKYLQeMog6Qc0KWaDi
dASTOICL9POFc0Pq8H8OxDjvbvegZlithsHU4GXvkSnkR3iYICcKZa1pEetwUDgZ
vumglq3P+H7VvIXhV0Kuyuw0amWP/9ijJncx0ZrvdCJGxF2XTyzCLg1GHH0CKSea
TKPK9MF0v/wA2v9qnLvj+cN2XZ+XWvKzUMDvqkVb3V6bBneUmRAXxFEOpjS6Xk/z
PTC2qzjVm/Jz+4TdpuRVF3DttYZT15knN2MGM0O0xRzwwVtK7L/l7RdwI0Gfun1c
OrCHao3j9lq+81kEI2LG8Eepxiqzj3JPqU5Bo01Le+M3lVrQEoV6t/2Jy2TU1nw7
lGVGum3hLQjC+Rnpu1QnW5pQ6rFe4VS3l4BRPMBNPADoGeDJdSWk3zMRw8gDjK6z
F/BGNG6ep9johZikLe9gqlDhC45itAiOVOs2VgFpuM0BJeZtX0G1KIiDygXMZdsz
8FKOfCXThl8cFTrE6J2ivKYeR+YnTmfdC/eLFeIIohcKLlVzM07sBgJm6zMlDYCP
jKqF0KZy+irlcx9xxqtMG3N47gRdAjsjYDFmOgQ2yrohc6JkkMUy9HksbnqcRVA7
SuzizHSlSExM8ODCaWOQm048AYL6TI+vFnfxQeJIPGELBsEi64F1x1wVL/AKoPEu
AG+dvzzB6sGR5VtH8XW/bkbDg82W7LB8Bojsy6rla6f0h/ube0WWKhW/xRoItMk/
nLZqUc/mJ3HUH9jV/2Is8D0Atc6eIZC7A5WQmR9lX7Wik78d8ypm06WVlQ5j2KWe
xZX6/V/2XKbmsG+iOUjDGHlbnqff1FekErXe4zt9zGkph1aQv+yUR7LdsD0/Ajh3
l/O5d5Xva4hkJ70eOgw0buFCX/yuxk7Gyy+GZaCQF80czb78MLSuCufvqaPfc0T1
be0Fzk1wGV2vlTd4+4+kuFPOvLDG/+RvJ6ybmTXt/zB18DzuHSSSi3uIrgnzyHzl
Q64EL3n/be401FP+80lr3BS9DSjH0eMWAeUJVALxBX/KGwO2CV/b41ySHmcwmo7w
Tm5kc1Aeaf8y4niFi+i0WZpowdl4VgtMS420dZjpxCIF+FkoucDHzNyAfwVcUtDX
4f3fQmTq+K3I4dPEU4asX2jqAYeK7kKRi8kA6bH04SpEWpOD/HlEHwiknw/yBFRx
zYZHWztjGqIRCdq2UbLAQ3vwL8K4y9rmQV7pkC64THGL4PtstilXUrPaMZX/NiJf
lTmsjY6XtJFFVRBUqnb6peAF1EgrykDbH6gY6kbSJDPyaEHB0XJ9jBj6MCNorTnH
elik1wm654X5SROiYE3Wz3njLpmlRblrB8j85UBpe3rZUsGTTdYA1dNnP9O/V14W
WEO51q4KlRr24rA/yvJ3PZUPBvQaHylzSlKhfEjZyF31Gh3UiA1Ka2x4hAb6vP/f
4vVWgfJqDtZvzRX9dutwq8+3kx/vQdmfwiBgAfqbp2y++iM3MfgYBkKRamCnHy1y
IEnTCvKy6s9/6fFKrCVOeck+hMS2oRuZMO5iVqYoVxb8TCFGT40S9bw4PQ2ymeE+
Ggg1EGuVdGTeQ5yfrLMKj3dCRMLy0DVrvUa5tUYOLwTyIRAO4Q/48S233Put2aGQ
2gfivfwExyzDRsaHbpGBQOQE/NJ0cxhA2Ee65kqc6Pk+YDCy6Fr5SCASRzZgK4Ol
wQD7z9RAEzEQWXjL2la1dfQTXY7iORzFyq0MnkULdRmgJUHG/ZDGLW0/d7/R6qiA
21OGT1q2f6ac8ieGiJojv++qkfZag/DjIIdAZaDaWmZWtD8m58SGxWtnnOW2zRPF
yI6eB2t+L/J6p97FGA9ilvv/nsGam7kxPf4DcVL/CFw8EcYOYz2e5uNDRkzMfZ2E
6TbK4+RMmhqC0/twtfQXn1YxyPsL3pu8sI2zXC9QkqGEYzjOl1MsydlPrAT0sdj2
SLHGlUdppfcRkstAbpRs97jGHyJuz7obHstHLPThfDG4E9wI3z2FosNCps8H9Kqe
plqRqLMceh8iT/W410U9kqHT5UYqOzz5+NJ3bVAWtwuKDbq735ND7LlZbU8oIsqD
BEJq/cU/FZs2VA4JU/k4bW3SeqzCKnse9s6mqoqEaGmtovP5VsdYPqa8Kcj/ckYQ
u47hBqnAO2QLoHatiMqFhi7maSw+M+2CQdzMSGpZl8aETUNOj+IdWklZ/Y91LM3S
e6YAs7mfYhjgLzWpgMCMcCmWOog+HtXo8P4EoY0ABVpp7hzIQZs0s4z2eJgTKHfL
Rrj1S/Y206AV1o70/SYCt2xIlk2UL+59PzX2shoMt8aVEsslv/vIucGZ3EzBkJE9
14KE2YbXOudbQllHSsQ62pgHA6MotJI/4hGaQoAhcyKqLzC/v/OLf4b0g8Jvu/NM
3kkNaxuYu8j2bY/vpDXAmSqjE2uupnbLF8+KX/YKTYvdGWVAckXyW4Ex4gsOpQAS
lUa88mEiVxnhA56Pl7uB+08a9DOclodcREE/d5l7vpiLoJxzjJW9k4DWolycCx6C
ZCNgzji20xo7XBck/qnZGn5ZLrIrrbcsbjva4w4e0x0L5jmBroc9/cfyAzR3+09M
qi/5ILja59J51Gojf9IOpZnWeDhzeGoFnWVFTDdH6rg2sMDlYF4he88SWeci2Q/t
DRkw7LqQf5uaLZcBpKIkR3iHj2SkkU2jQNmAxY9Yu7Qe0kf8JLoYnErJa3pdQMkm
2B0gL9aUBmuCa5kk7MCtx4zkalrZwW32OstFw2SBp3l10TFMVJibqJ+4TE8owxFb
bULJJy9/w7TieN/GB/mQ0iwCvOb5AFGKuwRY7H15OcuSwDeDdBIQoVWhRSWW9ojB
aDDd4gRjjnPRaeHBhnwREU/cph+IpbLcwP+9qAsOmRUCgELnYDK6JLR1uBZo0Hf5
LVnsLoftt083kcn+/A6BTmYWovQWYiEpXv2r7LxMOgF97bEE9rW3XVytCvZXzZ5K
JGlvaBkPUZjCG89wLFhWPdRmi4+Pr/+uvJoW8avCJanrZTpvAnCfrHtiDdS3Wxo+
T3WdAtut4wdsYpnwhBjyk3hWHQkwnr0hUKx6q/z3e50wCD6H538iOvSLv/HSUqk6
ZOQufNrISxPQ2FvLo04Af8JGhgNhfCy/C4SGTboLCR5/M+dZFE5sFYRj+s4T4gf2
yRUweCDEirO4WiUU3/p9ayluehk/B/xgO3AgnRBDRDSEcLNVdj9lUUA5mxVQYea6
6aqrGGpaQuCwYxeYL2Moyss7rS35BRgCv/Q6PUXAx4ICr9m8m/2yLYpYtmUYfRE2
lkfMSTpZZP026zVqnjiaBCct6aqWJ6ZsemXljJAIoY5QiVgLQ0mragjgjvHaAoK0
Ox2sms/aQkZa0CrIA9l3ADCwwUn5BL02s4u9+ziJn6Z/xKkO06AXfgtz1EmhetpG
pCWP6qV6ecszNdfnnwVnbqHUnRX04ek/vuKEfWXqBDMsBF3+Mhh3SqImC/IioOfI
pM26QYMsudoqd5wW/9owknBT2dUlR9uUW7Ddb4r9AP87Z0kW1RINV3YbFjfF/pm+
D2Ot+mIU0X+r9zwwTqIvD9uTgJLe6X9R5K4CYDJhMYjXJE3iWRkiKaVOkHocqECh
nZCh5d+SUZOQF2P/kfrfHADm5se8Yrw34kTZIdyMqwjHf8y7gcXfGdJhMfPoultb
si/3Z8jLVZtERUXWgOmQJZZvr6Zsz3hyNVevYfnLkIj4//5G5w00PxyKKlNqQRmZ
fv468XV+XNm8SRESZ2tv8vtn7v0254UD2QeUTOn4aurU//cumQCsjiRXKI5GwpRj
BTz/wWv2Po/+L6w7ajB6iIdJ9fnsBVXdJPSQugw9S5QgyR5pLwRwDWV4D6g/rNMH
zDvFOCJmjC1oKsYkqExEn1jntV5hVv7xtDBCjTG5qy9UX1H+hgmfr8QsArGAhWl+
v/72u75JDxZ7lUMZWiZjdYlHf2POfIjVVcdQro6pJ95Lq6xdKOPYpD4ssDV8DygZ
jvlfNsyPjz5oHwL6XuCepJM07PNrYaew+9M3GzSYkEGIcW0uaNz2ZjXWQKT12HDw
XIPA8ei7OpiXpqSst/ducHzZfX91CiGkDyyaO+C6c1+rZsi1Prhzr5Sh7ptIYPyQ
mb4LpV+WV6GfkGUVd2e+HH+8RH8N/N7l0awFFuLTJobL/6z2V9KerexRxl8oouIr
XLXDCB5Ki4uw/81aVzhLDCGyB62GUN/xkFtgLe5tU2uP5CxgFWfIRcOXOvSpNMt1
L5Nc2GLG1tmHTBpahrZzMqKXXuGlfwdBtTbzXTK42lWQPdQSC05CnBwAyTSwMoG4
wNnrendTVZ4w+fEtLsEBumQ/NyrEbBtweSMeXSklOoVGJG9smC0kwxRzY1ygyXwc
klL54leP+120a5LF0XQoA0f4Qs3JuC/Yz8uO/6aYbWqlGa5j7EMNsApuRmKUKjUR
PTGmYEbBsmpS7wSXaEsMRyz9miLJSMd5dukpJez/6AlZlSlUxiczd1D0HXDB6ca+
629GNekFR4anEEwYRo/Xqq/gi4cgSXEpJnHi10J8vxLJVrCM9nnMu3o1jmaLRHA5
MRh2FaHof7rWqMLycE1+9dbPy3k7/anW0/SA5GzGFnFgf2KaVVt/gzf4mmKcO+wB
E1mb7NWna2TVvxb4vPT5oXu15Ly18c9cv6cr/BWvuMQ9cVpftMKutafgdgkEkmXX
eJaJCE4P/ig5VZYiqgwENbByiKZBcHPLco2N/OfA6dNo800z4jc5pEDPvPEpdWmJ
LKDxcgc1ChSXNOU16DW8h2VxxdqaUWICPI26mNMGFSZ/OBEIP1oamEG+x+Wk6t50
c2uZn2GWpxqqC0a0cj29H4A4BafdsNG/JbO/QZHZR3M6LYvHkPixnrQTDZnoPLP6
MDsLHCRhqMPCBp4LfPc98xmduGbWCn+VYKg8qC96dslRkgTceTbylXd8l1wQEDzk
8YQRApfB6LTS7P+esr1lHCWCTMERU+U/jQEEW/WvFtx9m44NA7D+gZ0+V4qYIXTf
xudez1RXwzB27epSsA3d7KPu3K0S+S2LJKtyRfCL/VZelA9NmF5TiY+fNxy9Uvfw
UNIeDWtYYou+sNBENIi1eLbs2EUwnFc6BBfh3s1PG3KVYVHqB7WXEGQeQfyubyfq
fI+F5j3gq+vk6Wcb8kuxllOsN7mZDV2Ww+yG0PcqgK5DGG+WqfmgP3N7h2uS5oVs
SiCrOWdEp2S/eoPvdXPVOwLTP+EPLb0LInpeJyEIF5X4MJO4Zjm07ZLCh9Vsh6iK
kfX/ZO4siWSdAmt6T+gHDnKzbbFRjS/MjM1OXb9i0G2igPTkfsx4rCQ9w2hLSFIy
DmGiQJXjD+xlZmW5ew2TetjLLQwMLeVeaCNFtVc8p9C2PEzUoH83mX50wf4ndezI
EJ+MYwSwEQvPVQHOsGsEJGi0yLGV/v5idSVcP4t/tB6xbEWpqqmM45dPb9VKd33O
mMQLP/unitf4t6ObX53pGziqS1tfprSP9PvXO+cwjQ8MTfW6DtrcGioEZ1wNIH/y
p2HoOVIlaH7eEBRpqLuTzHEySXqQBx7dv9k6NTLEK0pto8VcC3CSNY51em1+9+iJ
h+frKe/ijmdXts07jTdDzGVzcBtd9U8ZXDxnvP4Ib8AzPi9v3NocyQK5iX9eSrQt
yFPhKcAuMXDWgFmBESApSFo0I7wVMeONyUfXy2yLt22QkuCvHula9HWGNOH8hsZb
1Jj8pTtY0WvW2BRC13pq1Z6+VmizE4gvJQ5XfomFI7KW1/SS3xXRCL5Z3OleG8Rx
xP1LWJMbXehq6crO5a1U2dainxudBjoqRlJa+YNkbVux8I4kijq9Lz90aOopqn63
rTK7TXiR6JS5m8pFTsKmWox0SRSMTD7vFIurTN3ja1XrQ0i9hZ5kV+Oy8hh3t3l+
LC+MG0gN6YZxtMTvG8JDk7bzPyE4uqk/SL42czsTMMVgOq947pmVqOUrw+s8bnR7
ZNEO2NdbupEnIo4EZyR4aSl/N8MQvJuknLAoApP2saY/A9e20Kzt+xDTYO/lghct
Goz4vEJtZNGCzfw1yHVJAyVj12HQPa4vJUjwX5EcEGV39bwauHKJU1bxqnpk6bWE
bCr7T7U4vqMN8vAfS0CEG6TVPuK0d8Vj/WI9gVRv/d9LKGg9OWd6DF+V1aj1bODy
Yr0j+NEu/4Ud/QdV4nFjqT0rFBqddiF4hmWZDpent9PlAl20XVLHhPVr3CpMTv3l
4gY1+pBUgiJx6syj4MYgzl/3p0mERUOWUeP1kemgXSMLMEVHzJ8cjHdHTEzms7D0
E/JU2oRHC1juI79DPCRbC24tFdhJrfqFRzXHI/t25fz0tpgQbToy0R6n+eB+Hlyl
SpC7xNbJFboOGTpLZIVh03ZJPCGAUS2kyhmp/1P/0vVIi2146GGlSHuE0/VeGOJn
wBY301Yt7hHLHWGkX7Q8NYnhgH0FhClrcKCTFXNeobXnOXeI2ITyJSSH0L8y+Sqm
eMuuI98YgtXaPl9nEXwghnZeh2U57mEIqrBpvsUlpugxcHLMhjJdaNVRVTgukP33
goeZiLvCLVaP5yKnIZUEylgbiP/g3OO8HJP5/X6Yahebk50h0fI0h9OyB8okQAer
Q4rlO3OiIRAqEobqZ6RTMYRUW5zpVDG4LevILz+32uAbP95VfQSGiYlrnnqLu32F
F4qhAH88Z5S3aNp/N5BZ9Z6pkGF2Okk2ppA+Xu4VaLc1M6xHF+sYBCs3lKNL76Pc
hqa21ju4nULCYWqbCIPnnhsbBuGy+pCM/4Ai/7aWqIdxJbcBUvSWPWu5oYM8c+cn
5Z6dZ+ljHR2EijwAufnzyV4APmES9cVDIhz8vhUHqbKZtVPehWQPUPDM8BC4I4bS
l/hv43UNztM9Y7BZxRgcjI+jObS13XLGBmV1Tbiyqk/kExi2lVhaIuaz0pmrsjHr
hbkNwTPdrHtBzOB5qySMMUyPDae+3hMkXmGnIYHPKgGuuEmRqdI/QtFgo5MS9MCq
B8yno4xZD5JSKC6yrHscfz1N5CvvuMg3N100wGB0NykXJUGtFp1eKIDhchHcZLaN
K/jsDnMT1dTy1ADps/QsCUjnmezqT8dEUHJwftF7SOMZuemKowdpUtxlaGRhe16g
7gJQ5LIK+lkbsYbZB+j6XjwKLsZR5EARfKLOaVzOmNREC0Gvv2xJlwJawTlhbiJ7
1VA5T3FpHJCZ59cipYOv9JtPp+nLE9qGWPNcTF6TCYY8tgJYC8XkVG7TLXOcTNsH
knR+jfpyk+2WvRr3MozaT6c1p2wdpRGKY/Cpgpnb42YrL7eKRYeiJXVThuc/cL8D
bcdQ2FuggO0qUc0mw33O8x/SLmPkBZOMhgiGwX3d3KXp11B7adr8e+DZ5K0xPeIz
RgrEkpTx9vhXanJmUZ4uY7WsIR070AYh+kpgK1/ume62z1YqUP6PGStFChY7UvNC
s7PLq5ceQNrXNBPSoJb+OHRO9Gl3csXORVSgf0Et7+IOLXt4rK8t+bq8SfmtTQeT
MBwmxoXlUSPth0qrbdIwJ1fx1nTLtrhHZO21PYCUjmirqpZ8rhllzvzevF3YyDWG
i2QZI1Z0IdG/M/3uGB4Kd+s+E1CX1hpDR9Tup/MnS2IfHJO45w+9cC0pETqcjOzI
SGVlv9yiwG8924IbtBpuYzGVrOw1JrtEZ+jMvRs7mMLIvkKCjm0GXuVksfX03u3T
FPvAv0QkisVB+7AiR5j1ik3ivzpMzXHFPzq0E/0B1sqbIa/zP9nA1ydebzKIY/UF
4P4OfuRJzGdSrKCXbqvFTeDfcZg89OR8q6wvmSXMABWUouf1xdSRiBc8UcK2J07N
hm+7/lxvLY9myCuTnYLFCHX8TijqZoT00KGMc+VYNPTc3t+YpndeQCUov6aloBvV
co6BHFZOrkoz5V7Kl/ELs+EFCoKEEQPrL3MJqYdUuggfyydbGzPsDpY9oM1u9ESQ
EfVT6E5HCkeH7xqCd1HeqFRsQxgOL9N6TNeFBMsx+drlamcw5XCRg70gRjpL5gG4
8WxCnXmxaR13Kaa/ODo8te9JZlZaKuSzjG1I5jzbulZ4BYxkLmfXfOEAmp0tpctx
Pv7mHQtnLpLsESWD1NVxnlcvtY2jaqSNm8JL2s2HVTe6tmGS30dVkEGcm81/bzcF
F8fZP06CSc60+i0xivWj5WYwEmAzPftBr/K0EYOc3KRqyve6z722/vgWkLqvn93l
hmIx+7GmArcb70t/aaElFEmtFkMiEtYOt9opy0dlJNZ5X0cpaqJ3av48eijM4J8+
fYgvB8bOBLns9mGWSIDCPx7qZL5xEGwFz7iKehd5VDJ9WhGgugVjupBfMNFqVLbJ
ycYe8n2ZSiE+GLj0Pqcf7/HTePuClNLp+rsydNEDa7qiVlPyCG2walz8+It+8OEw
ljo3/yKTL1lzR308w5FXRS6VTwn8udCAhuOgQPa6wSJcha1zWW6VVEdQpelSheL/
yvpYg1HnUCGuDuisPLccRgsp+oRjS1cJihtVcjiAXI0iDFYTsLJnqPKvQ954hbdR
X9bbMxjDQQIP+oA/a/U4BELeWg/yDnqyDLLyShzxMCJaMe1cl2IOJ8s6e70Yltu5
7rit3Kf8h2G7L8fyTP/11kxUZAi9l2iZDLGmxC1rRZrR0zrlNz2vj/fhShMeS/Le
fni6qdF02E43vrwfXw+Jv4gl5YAkKHmIj2bSYCEZND3jN54Yr9OvnQ2bpVs6ZBto
3fQV/Rjve4jAc72SK+h9vpooyA0xpk6v9CXunD3ndeJ9h5qSZsgXxvgJM3zjK1yI
SfJsANUStXYPB8zr/J+JjhOzUfJam6y1PsPC3VHowxidKL3PK33cpLj5AFaDtwv0
nUpJRTiV2707cRPYhD7ie9OTit7PFRlGfR9iZAFTTK/VrwGXsTwpsdBDlKuaTf2M
fqTWu+Ay0n7NbbBE6ZC14iJefEKr/zFnI1XMMaNXnkM7KkU+m9abUSxUpmrFbxx0
aNHRL9H6OhCmhKMJ1BOvEkz6IwgiQc7YM8s1azb6fzMQqqgDA0AflYYqqaVpFxBi
IbjUSsevebLc37ZzO2GIFy2w3K0itvTtHOkj1PqDpC0qIHOlT2h7gpVmez9FbJC3
oPo4AoFdsAdIIvm4xogMANixerU/R48jQELSpG4UTVVpJESBLsnicyxYZLI7bkys
DVqy3Cd7a11JO7NIgeNmEnGvjJNIVS3pgrh5ZrrFTK+daxrpFPHrrizSURDESx6U
0p9KFJglQ/ctS0GPXdw++Brkl5iHJ24s8LLmFuYqHoHeOnial4N2ziaa7wqvFhSu
WDsejXMcgBUDLhmdEwM6XmsBFH/jWPYIGpV0jGA84OmLcwWRck0BkCiaMya7tzd7
2/WdOgSmJLRYLn0FxSAtgrkQNStOU2+3h2d9r5Ey0cIUoo5EpqeCabRQ0+E3oIeS
tYFOwS+GuTViql0yH7qdloYogO/hhIISXTgjwZfqU1UmGMwyA3NaNSBWm87twJ1S
B+9Xd9eMrT/aXDsEQwIfaoCrB0xz/tty4AgHWB/xGbtJvH/8dcESs5+/lGhVCwBw
5nhOLcXrFvgW/S3W0xyWZDTICQcdyJNouBeYBChdB/K/txP1bKc4m9vl7EGZZfr3
5VlNub0DxhTdBvmmrhRMzeVINkxn1MwAPnyKGhWXFuSlEHHAge7I4uuv+bTB22RB
nN71SLXP6W/N8wYXtgBF09Tid7iEP4rzUXx7LVSFvFVXD1aqDz0orRnCuUP/HCQz
g6VWsB0QRozLGJG20RGOkjXn8MvG2508LYVa6V1DBThqOT3uC7hsRCbYoydtngyv
d9NHg5PaNaVwBgrPGrJLV2NZPGQ+sdpOkeJUZjjnPU1aX/O8lQ+jCYvWTWG8Plr/
ZTeNqrY87rD5ym0ayZOJBvMH57vmBANJGT4IbPxnUTosR614rjpXE/PREdSnJbxM
bf1CuiRcJ6f4QvahNNFmZ4T8HKwVJlpP3xpAEXCo6H0DKbz0Rsn8S65M6XazJSFP
cTZq1DCewWncotKNAWTHATS85+GgcHKNGx/Xjauw0//EQTd5v9nrcU9felnCZkCl
u9AaQhdt/B0iOPHkadaT+kg/op2mTmhkkOBbW0Y74rqRYuiZbncNISMvVtZk6oOl
WJKIfDSfU+kpgafEy4hGt3hf+TQiE9eQRgm6fBgVo7PW1L1nk8vQolkMFUfIW/DY
ZQVS1+1xZHJt7V6uR73ZbPrJD77ljWfwSxaZWpLxx8HFVbBvl1XBBsHHrJ2+KrE5
jc5XMaIizYJavxPuF4nWmHf4ttilJVqKCQF4JeqIKig4nVTwu5ROSjAUsZL9bVMn
Qco5OHbBpsvFhLOtG+0wgUUIGwk3odnmqJQ39FXBrcHjBReLAY29Ke5imiHxh6Fo
1xFu2FxoSrb3pfadSuPZ9G2kfDip/u68gIA4pqb0i0RTb0Se6swdMXJsG65p5wW+
O5y0VjzRlZp/tpac5RT3kAQsh51A7CV/U7hzlLVhaBG+fnG2PY8VRwT2OQ1YVMgZ
l5W7+r+gchlARYSr4IGrHwA2px2Iwb+oW9qYuZKAH7nWBQFqlzJiWYhvbQ2vMrLY
0GOcaB8tjhdhskUgGIbvHseqB4HqBVkVP2P1VflgS4qWDfnzNtBBZiODsrwltfRK
XZt8Qv2Q9ve3s5lYkz8jSxx9obsJvjXAqr8F4IGpzNCxEq4iBDsaItTSJK+k5Rp2
IaT42ZFUMQ72PRSeK0X7ml2Deblbq12BBiBGw0zk46HEm3D5YlOsJXw6tcz/GJN3
MW3fonPciAnJiS9uH4CBc6bW7X1HLOzIbQ5Vdwhn/tVD4AjLscnnO/17bopsPa2J
j5W2ejSDC4XOrPkCdO3TUy00h34JkRTMjwmOHB/bujYOhNuCrse7CwdcvSGBejXt
+wCDhp7d8MXThm/d8kru40syD5h1vKbxDuWk/exqjKUpAYpMbJnsE/aERP9nhKZT
SiRGadl/v/RrwDgAKmlI4s3gTxAqT1XXJIbZiJg4epG3Y+NEyFnniIs/x9JWIFOq
NMlh2z7G2Ew1mK4Hd8k8ATn19VU33h758nGo/V0NcVyreXAO2e3Ip+OejvK/Dz4q
f+njzHQWUzA3+7IOtK+8Q0n/oq0aI6xwOJfJXtTHSjLfKS8Ajl3HBPORHQ3B/6W+
+OJYzO+mFglyniBeb/mVFF2qPGOCLOm0vImWTmeCJY4sjiQZdHA6DVeBzDVVCcm4
jbtxsVuzKipbkJkwlF6bZA889J/NxJ6B3ifzpUqzAIt2B6fvLZ4RNsdqZfrxcsbQ
3GZb35sMT6L5J3Ubby3+9Ain+fM9cSS/FtgQ5o+zPhz6ATZizlUQ0BwtBbIRluis
24HuwfhEnCIJXXtTDLE6n2j17k+MtqQct6pSWn1KmNBtBe5YMr0GTdVjipPr0FQq
U3m549R9pJagRjhIuNPaQwSftSlmobougvZA78coIdjK6LaXxvJqkc6KCoc9GJH6
4UahH27OSd0LHJhyjNUV6Wcht4E+6aSqKoqIU7NLQKMLZBVUJQRaDxdT4t4ZgGNi
Brt8d+6LWeLWFpJ9L07dxYxTBivNgTZkn0FpPsD6FkFNJiQiWi3UBX+jLcNYF0Wf
pBTFM16zQcFNsUtz+MFBZjciZkAPJlncgo2hb4VDZp1Ks+bNEDBzb66gbJy8Sy/d
voeXe9MHHPN7vRwLRMiK9yUn85ztYoFyFk05RA8SoMyqEltwLFssOt/OiHh3U7C+
AP8z/wq7KUDdTw31ZtbgAzXz1IzFAv170dbn1dza69OjSfIIXkDSzDhxwFI6ulLt
DFpmt5tU5SGanzS1WWAUwpPNdVyZmEevMVCQqpzNhWrf0L0ANB8CP+iGp8se4kbx
Bf3yCPRPtafJhbu/JSKV/Y9oGpn8IwXHdy7rnq+nRyrBNzN1FegHNij1Kd0l7DvT
7VoxyTziGVTq3Wi6++gLbTB9Tw95Oa3Fi6P3Fd5hHw5PWhVD614cx3wlTKmcd+Rh
vzMoO/i0hOaqiKCmm+N9p06FdBSJJjUjzzR5vVLO5XBSFRQiyda5CtlC9VzsuYev
if2rY32HiKIFMVLaghX7IbU5JPtSQbkeV31lsZw902AKO+kSQC7lZ3cVJF5qzA+j
7ywZ22POV/HXl+pzKXNbRheSqYgYuZjpjRUZ5X/10N68KviPbnyvTIPUdf3hjTCF
7dfCmJtWBcFDFU+pPcZSiPdHNhJavJf7P1vdYIVPyuTnYcQz7nX8ecMWqre0/DZj
BjilPpI2gw6wYDyGl9MInbt7lD5DDslIgX5pW72E3XScsRa1/AFgk0XJDHGh19JC
ELCyr2pObdgw1CjTnomLQHxYX6lv/ihiKamPYxEybULjV4WgFsqSwnfdf+qkXPZC
dj2JGMx1kYfv/tLW68rQL4YKxCn3D8IAdtReZHFclSYx+6Pzniv3MyB+7XE9K9wH
kddCm2/bKEMQ5WeMcI3RAxaOwfqHunIClslX5h1z8Tr7RSuolVzFiuoAF/ZsquqN
j4jE4Yt5SuaumrrT4tnCK2ATM/EkZnP9AlxhJzV2WlXizh1AbAR758fV4Agbjy90
euJdF02pqBFauKP0cjP+i/7YHBaniiq0+bwgjLHcHojaaBWrDLPeqY0GHKgfRPhA
OdUJv34LcWH/OEHnYmBFdZ6jjJx4eBH7Wnyxqlflv4r5gZ8TwDUKHPaTlU79SuKs
bWrDz5+U46W0W3Fe2m1Zjtqh6eM5ZG/Dp1VWSvzftdF6EnbuviXzkaEBe5J2d0Sp
LxCBNIdyzNFmotkBrsRQsvZJigptwNQrfDq78AmlGxdzx1WTPb3fA3q6PNeYaKCa
czeZHGYe8DFSgtEwxcpY6ro5BCYneHzCIekwDiTrI4wtzckmdJRAFmQ+xUOwI2oq
d5TX97rDFM6zr6vYJvh6agXRtXX0tmLfKgnAq+pV9MBSgcYwXJuutvk8fn05fJDA
0g7qOmbeYZBNOPXuHM0eVJl4C+nrATSbFZ95QTrRlpn6zd4maedDj8VIoJvbd9l5
kFKjPqOUsRuJf8xdhqRd2aZqqsyrid/vU2YqZn5kVl6z0WrF+6ZP+C9sjVLMTLbu
RH9cJQAwkgdOCdHt/5teff9I3DYq9dTTElE34Kf2/xLe2LwfHqjKpOuo/4fX2svX
z1M63HCk1h2uKv3ATM8VVvo4Eh7PxXrXG9/b+lfFyd6sj876IvKhpfyRJFHpmxJ3
g6Ij7n2nCXP4xjlpvvEBPiTaKFIPoR3/m6WFrwboVHhd18zBGzSl64eVnJiue4Zh
oMxwYrfT9Cs573Aa4/zP3MI0K8iQ5kvMAgo3U4ZrPfzHVTNCIKjKAbPY75TkvB1s
JFYSBsgJ/QgYHmIw+RQBrUgq+QP6SCkZwq9S3sfhyJdit5bKyrRueeSPogxINevb
Z5KVH5kRxWyC3TIJzFZu8pGqjQ2ix5G4Z/i3uiACVcsFHF8HWjqPNdkcFTET5aST
yD7m5Z1ji4PNJXeq7+xhD38Of66JljCbNarQLNrtjYM88muRy6RZ9ee2C3BRm0fs
mWWCNsrWnsvxrcvdTEQs8g+W6synNJPzFIM2utWUIDIJa4OhSg+w5qZtQitcL19g
5o2VaUpUB7WXHjZnki0B4aJlT9iFBJ8HZH8kQEC+19ta2pcW4M8PNgEMBobMJ3jK
W0R0NK4iBjeHCALKMdeTVAcYbSW77Qu2gy5rjIypTLbW+XB7XC1asgdmjPEdkbUD
m42oHtQK26VzXtPahquA+WVIaf5HYVzzJT+TxRx3LJCyDEnx0aUpOXFTFk2GU+RL
EUrlTkLOoF2Gn05l+urf8VAE8qVW5cQi01AdacwfIyYgFakT/60t5SkzpZDu3nDl
ZyH1ocUkYv8DTIsIvtCMPbLOY39Q7/TlbpnfKTe/KJ+HfZETbNJq1BzcGSGDzZZb
Fxg2AIZdM2KU97xBrDk5oAiF/AK7xQDQuEPRRKaRTxyAVZ1vRddCmL6X2Iah1EKd
JePjOvAUUQwrFY0SsKNt1/+E4gtHZQzyzzy/17ta7C53i5zRcWBI0J0scAjVWc7g
ufxwndZuMAqOsQnaf0jtbwNYtm9TwflJ4VniB2iZIQfPiQo6QQPBcIe3nhxfEk88
Olg9qvY+DNm4GRtOhC98vvPg1A/dOt2rbe6soiuXO1Cghd2mO3VRkQMyriZ45wTr
UU23661uJWmijGbKD2OAKDCbFGLXFSHiAVPYPJ9p3arEPJuHvt666UgQt4gWTemT
NxofTuikcblnNVAz/oCX3An6Dez5U65ISd661KXVdz+PDUmpnTDuwa+tMPCIBaIp
MdoHCMNi1WbkBYg5LanxtBQia2R2rsmzozuMueSdd/agn1lxUf6W1YMpUkLYCmt7
N1Uf6JxKl3+3BntJa/TmnBYKM36kWBDBvuhyyOr8/9XZWXGD0hZpzCILEq7zo5bO
jGsoLP3XMpe6tXpA7wc7Ukda1WtrLCUWN6Uk0qM8b0Xo7wK4/NhsVL4fw6H249BE
7ToeIcLHh3pxs6b5CdPudODLq0+jQn1wJmMMjG7yumFw8hU+wh9VezlJEcsyMKt7
yjUefXdbMlCAnrZW3YShcH3ppYUFaW3V87MaNL2IuBmfwMp+azowLfG4lol/Rq6O
tr6tJs82CSXtUBMwHzs4ksioDmlh16d0LM3m7JEEipmgifuzrZsvZqCHSJQvNAri
tNpjus8DvRDt7jAnH3dah+3K6gYRp6pmvXV2Ye3T2ZbaIRuIFoK57JBtP0FfWv5L
v++9HUjkpXOcXcoySP8AW8V/YvT0Sqw3pUFPjqo1E+/Brc/HJWSeulsXfnTZ5o/6
jsDZS+5nKnqZSz6kUVG+6ppfzY44hi6QVpby10ZLn7GWVwRem8nu0QiiXsEu/VPQ
RHdjDSQr1I3NxyVxEg5Dbv4EknelMlfgoHUPoHJ6mDpsjxITQbBs/oUCofQD9g9h
SB35E2UMfNSQ8izBVDsuzCKv3zuQAKygs3i4XYs++jdliGJ7mHUG2VGx68+q+iHS
t3pPh6vteL2ptnCjQ3vi2CBB/1pnXtJZ37HIKydDPBs+UIudQ42OJdxB23Hrdi+v
DTl1K6S9yh4DKlnFyFbP2W3keP120e5v+3op3r9MU04XWs4FetCCFAljOt6GXqTS
kDJ2ix+0hfu9Gy4fZTGGghBZ/6SI2SPLpXgQYOr/m5ezkwj8aRkX3IJgvR5JeiXd
VvkEkjl8rXI6l6Fhp0MNnEpQ0A4FLJW+3OAyWdJyNY1kfzmtnr92UY4g/qYP+oG3
hZTR7CkbEy3g71ws5gtTGBgrwGFGaqilOgHNr24X9PlTcrkpTtc5C6JRr5ubovy2
J41/Q6A1FqlHu58jYvaXs0dlwFnmOFjjjt2aOfGbuJvdRWp+LcpMbRxBdN1LSyx+
vHX82ue/RscBkGW1PSYaFSzxmoJiWl9EhbOu2CwVsuAFpvXA/G61qzj7QUCBRWAf
v3lK2b6F7/WsA6qtFtSxawnpc9g6Us7KVYU993KN7bsANb+yBPFY2qhCaxZsvsc1
arS4I83LUPYjSt+jWEzAgmHLe4F6csDbNOo/SyxhYbtt/1H9D7qccalDAB+jpcEw
CBc5ByXiKUFwQUCGzVAqxHrbpI+YnqIkmIlieRB3+Zs6q+cZXVcJHdHPqGnlZbME
8pHjQ3MLjpntHCY0X/4KWA47hXpAIScwrP0R+wt+XBRCCVYH5b7uvf/L758iLwfm
HVGB4zekNJ4XuRavduYfAuHmLARM4nd6d6/eYGYeuq+Y2HZ+KdmoXKulHeoc5UvY
IgMg0E0JAGCCaW1OldSMIxapRPAN4OSfbok5SPGwXKhyWeZSJnHVFM4KXw9L3ZGW
5GsYs5uIlN5LiWeaJ+tS3szF/IoyLXht4cLrziD0LczbC0MYcV2uvz/nVMO8O3vY
lkQweQQozoV5sc+vHiPVuvn02HCXMjfUEH5iBnnBbBvA5jd7frZei/l0yTpc5x77
1gLFyi4lQF5BNlcw5KrVG53NS8pq6V/s4+2CxJiBmKQJdveRvP7s24QPL88ROm3U
mJEr7hJYBpFcDQhsnAYF4YWgrjN+4QEQdJtFwFbbT2yhlEVAl3hFKod28OHhg8eX
17B3mk54pDCukIJ29m2QTtDqFI3rhSnBWmCHYOFAI/UkmCJ0UARpBUQigPyCs+7R
a/hIAtjvr9sY/GGAwiBSzhkjprPQhJJqW+KORfj/C8z9Wo3sz+Iu7XSJ10JljLJA
QH0oFkBBjHH25PFElQd3pSp1Ej7c2O+u3LB8h9eSNqf0xEy4GSl3TTignauGq6Pg
zmnOiJYbigDAIaRtU8d0FrQkPT7COntoo6GWfn0Hz+7Ur4tKDJEHoHvUP+U1zRJ1
jINvPwJFF6xX0krp8hO4SSoJJV5IR6evT2TCXfePmhMoBQi/naVIp1+EqKVycBTE
vbfXWTbNJhGgpEz1uZmI+Nr/1kXtl8w9tMDxHOCwHzZOhQv2EC9ueeRKnWUMGcd3
b0jTTyLBSZxqKRYdLDMlbf9DzRYPIJhlUja/bHFuEl4lBTaojLkGYjrZsbO8WBDX
JRpNEZmvTvEenUzP+T/iJnGmPJQfqOs/BtmQKFNR4AtLfBV7BpyXvzL22ScfZ9VR
PQ+7k7GFl4SfbJmknO07BRp3O6Rrn+cIeCIsMKCZY6LNqkSXgT2FaPX8t2rjepye
Y+cqaZaKsyGBd8u0SkZ7FYj2urDDHryhfxchx4pV73I66vfwx2MQ8mQtmVymUp52
G94abvYG+/dX3UuMgSEdBG4wXnwIkm5BnUJ1ryTXr4ghpuGlnZKGs1XxwQgCvXDO
oz2+9rHZgNmse+UnXA1/5uR7BbAB1EfZF0sWDk2RJC7dwXPr2FOmoYC0FPFJWrq6
O2/aml2md0cE6knpbPUWDZEsg8Ba8n3TKo5/znpiKzySZSjOcvxGy0IJu4PE9PBZ
wAMEmAZjC5Kb86Oh4BqOYhZYmZcTfPUQ5SNdJbGPCUC8YMMWMUsNjL/CARhdd0Jw
M5qjRg3dDJlPI8EIs2zYThfeZzkcRCcrDsomIZnXeUXWljFyRa7gvGFjZW1oLR9Q
u9Wkg5D7xnSPydbVLMmfvhQmRxXRSVYeDtFA2OwkJhaJpdkb7x0xkZ8uuOB4xIvN
wf4zZiBNXeAVm4ZAyAPsTbW/Son3iNh9VV5S4HDDP+mZ4BmTd2tAUkaDyoT9BgWC
SIzCL+zgl4AaXK4U9OCf2q1HQZLEDvOhEiNE5Ph6ALdHdYK+pkW7G5hkr/cFh7V3
DdCDrVCL7X4xisIaLRKDaXe5roe6xMbsXdBm7CBl1PL/JVX6TvOWkDoft+mAe/4f
ZVJ1/dbACNr8GHdTeZu49v2JxDE2Wdnt9jFl+ZPaKybeB7XRH/cvWDcRVU3f1rf7
HAuLh0d4nnBfXLEMJ9FLLJ8RTrRSqHwGmxGWiT5h/qwtnhlPuElOu4X9KFnGICFR
tCSKuSEosv7MaFjyiLtM5iYA2vCHn2aHLXdTje1fdRGWjoH6n4/fVSr6rDGW0C7V
9ij2jze9YMJehCjGXTKwWPPXC+ud+wrnpd+NgxxYXObiMEhjaz+Up4zAChdJyXIL
FE29/FZwdyS2Rd3lv3Ll5sDjMdD9M17uOUQ3WE+h3y7VoEiSDpDCws6OEVhhnOXi
5B5V5373mJDIDUhY1QIk5gH/c2KA900GdaTUvrSTGRYtHDtLQqswSd2fkQJVQ00a
ELxSXAHOO6T3vvgjaOYLUXZTWVelN33Nm1/dPpSu8vav8wuMIUoCv+pcooJ3+ecu
cvCVEp6bjp8uIW1V0HnpgH2mllSXsqG8HgnesNSOdA1IBCtYnFeOjZEWffMXgXka
cDFp+lYliz7WzftA/jsNWU+nrlKh1OUl0O3XI7z/Vu9InMqJGcGvXxUlwWWGyxff
wOqPGNWTAZ/2cO2KKNGN6tzMLYB3LLh1fWCpyiJXyOfICzAdFiSCXPmtp7oMYdo6
wmPVaIZLeLPrAj3bGE44ifsLzN/qSepcu+un7QAZpBkSOS95z04ZBM2BZdgOH66/
Bjf5Efg+wUs4bLc7unNZJu6BBRQ9ff35L1FHnI+LQwXoZ/37UKa53QgTWLYoNlOm
vx18oXBl6Y1s7W/3sKAhTUhOp+TzMxoIswzTPnLiztl2fxO05eFyLDkx5ljkiGvF
Uj8szcbFI2SDA4N6UBC3TmO2WJ4nzXnVoz+NVZEpXJbK9C2dQB6N9JF3mv02Y5Vs
gj1hBKOBX8CopjsfZbNAFeey13EUMzhBEy1a+I5CDCiblXjQyoMY+m+B4dHBa66j
GbE1A87sxM2d/hbuByAXv5g9IqjPu3htN2Dou3uo3iUJ9P5aW9RUnlAEhF+wZsD5
jklGrUQ/eWD9EXci+BRW3UiINsowSjnHyGPu4kOkRhruiqp0u1yQYVvHKNYaZHem
Yjek+nAFQsjHfvTKL52R2D8K01WFL7R+B0xrs9YsmGngTSCvG0qJVzVlJ3/ey9mF
o7HVC7twGmBJxf9SujbogLZELYIUqshQZiemtb5xuBBQzcTxPRdGAkBcVEt3hCCr
3xXfKMK+LVvWjEweQcWZJEK3fYgjIr6Bxub3ZIw72yS0d5rY4X5DEgeh0g4EwvcB
ArKe0AkK0oB34U0iakGxIsh2HvVCDdgiOsQ/tcT/HZuVVJzWXJAg8jgwwQWITcbM
pFNSAYE7jRij5LLbRipp5iyHdOBX5c4owOcNxdvdXCE3IfZiSw/ZJMBEODZ19na4
vNhQV9mqLoLBVVfNsJbbuAs1cJcrk9ZDYc7SBKMFUFMoTsbMO89q8a1ouuX+3i4Z
vgaWfC721zPe+kpv3opptm69lrqMJiLHAwAsUaKx5Wz6172nKNik10TkP6qowr4V
lIFFTeF5AYX3WKwhCWZtUUXUE6WJZOy1e/8Eyt0IdLSQWmL1asXYnQqkt+jnRvI4
WEc00ZLhPXy7FXpqeI0cMGgO4QY43KzTRNgzvY+taq2bf6zPTDNdgcZrjBFE4Avk
vCcamCREAvR2Lrpryt/54KEvLnpqyx5CQuV7Jk1zrDKmABfdiPZW/GUjlRybcmAz
VO5/yMNRH0h/xqG5gWNoQs74WpXQrspEIrFVHXeB1CBWsnIiLWw/wu7CCda8NWAo
Muv+xzToOiA7cysSdv05D/nqg4VDXAIxwGaYQYkRB4BJAQuU/HkzT7wKn/nwXTeV
jaHNJMSfYBk6xvTRorCO9l/y1DRNvY3zcti99jaZe/cNC5dkgk1lNIqFFvP7odZd
O/aGYPwuABGzqZVVAQurFhORI1Un2UFAfSBVNBqy36vy2bO7tRHm6CZ5Ro/borax
oei1zwB1vgcdbbzBT81GYKYucU9U7i/8LjKx6gexymv7cggn3U8OZxMJk+In7Dv6
6SLQB54cIaD9Gp4K9JnHN8B/kBJ02Qy50EZfZOpkaasO+jp4H+zSgrEMrBV+hml7
e8v73Mfxxlc9XDXiDJraG97DpsIcmlbhObv9NnFDaDJjv5iX0y3+T961TGhwR4KW
91zXl5ndC56cIj+QDWoJlNuofNkTzkwUvBszbX8t43AWIiGyEb72Nq0tGG5ZruHH
ExXfCzdM6tip4axQz3gTuIf+FyFt6oEc6AMbVaBjgkEGH4x/UNVl6pxotUFfY7J+
8nJTu1uHpjhxd/2obse7AnqNykyHUEhoAUmaByl53DFhUXqlpZJ7GBi1orDmZFlv
riZj6uIwLFRMbQZVI5JGPcvQJK/iXDJsE73Gl5IMm4ep+va1vk8TqNEp+B77DHqv
AQnXFnA3a4dYGvTJJht++70W5sWiQe2FkDnDI7wLMJGBBk0ZMCeCfcYnuIJ6yBFG
LPpIIAkdjGh91t3I1SmlBUeZF6SrYLwaBD5yjmn6GKfgAZ0jw5KlgpvDOt8pMCiQ
yQYPlb3quRe52cGtQKFQzjFgLiS3qn2Ynbds3l5W2WAkzaHowo7EYXTUxRwC5nWE
xzajLfBGTSIa8GHiSBtlh9ZYx4zD0iFMEEky9LVhyGhBTfCOvFwUYpj7vR16QyDo
TD2FBmJAAL6EXhLYve8GIn8FEyAPMY+gFB4mS4bjud/PZqvV0Y3aK08TpOj9Qwuy
ueO48R2Qvyc3WvkOCHspbsfmSywvUbPixtxT2OJdCmbH5/HoAJxyi4uuiqIuzSmO
YZkqGJy3fQ7BweSfEPNQhlwAtOe51/SOV2kn9C99kisKaMC2w6hU3yv+2VxAtio9
TqW+87zM5KFG1OzQao10srGqPl/KjD7HmzbXFduDbS5z6pm+3nZYLGDwL1lg3+wo
E7GzTAcp/Eneiz4OtDxGJ4N0CttntzitIxhfIpbW2c9pd50D+00/jwV9uf+4gUEn
BZ7rC/HK9r6NGyv+Mr0US+TAAZip5AVgXI9Y7gx06lHGW7Nh934GTBSFZl9MDQdl
pUIHYvudOobXKFBqmGCtXx4szrHXH3EDVjtiiwOAp8syGhaWbzzh3njPz2xqyBVk
i2KK1O4LA9eE2yzk7I+iqd6w84AWttx7IRJb7z7TEyrMpotW1JEJlW7mly8rln+c
RYGv8pFGSHnXNpbzLBXUPikxsEmwXlZt9fT9aJwNFfkmbd0batEyim0wqxedGOiE
b1uOeQ3A7feV2cpQtXiXyzNYFZplnl6GZif08XkRtSsbfSt73U0ZW0N+Us8OXB3L
J/MH7ZHji17ItJstbB1pgy4YIgvXXPnBjvQOZD2aUpCw5jcLJQWOU9il7AZc/GPn
iUe9d3QV4BuE+wxcYI6lXW+TMA8DD8rGvvMCCzbRQwpN1loY58vJM68gIzUv7Mys
C3X9Qonk9xbZxN8HlGv5CA8Fxn1cRqhhkE1wPYzbKu5tYha5IfaM6OaEI05G/aPx
0hiOzmKbbidCgAUkDeYPNOzmF8OsFZ9H23605wtMpfesDhJoPlUrxdPse0GKC/Ad
4lsu/wOuSThf+5cW5lvpeYIlfxAf2dsGSPiwKjGWomES/OkBXDd27gBP6Idl06jP
yRc1wtKGK3pqa50qMjokRFkVCoXedktL2UEwz3/km5MsN6ZXgvfXdf3eYIc0HGCM
DQQU4O44eKv6YsWidKcg/8Yp6rYWEnb3UHlocIHop1mpOnEojlPOK4kqZAyVybes
9SRqktoCIG6xU5c2eMVko0493xbCILFp3R450AT6VnccYlAF3n+GgFjJUbjqDtuC
WBDpBBiyjOJdZWn9dfIRXGi2+/+IffO6FSNT5T/O9s2gq0xFa0jt1kiYoE2Svwlu
Mui6h1adTGwqkZsy90zrcd2BVVJHbATGtFJavc04aFD1Rts+Rx+rmd6Iosbkf/Uu
LMSPU7oJiNiFeNCX22ND7uTS4y2+4I9/xgldY4YK34ScY/UAbtggW5LgEqAndeeY
nOUPLP3TVEC3tiaGvyRWJWgCUcI/SBhXaLU2+g2jZ2L8cHCEwjdzTyVfEagBD0uO
zodaFQgAlN3sYjnuUu1RwAycIFnHknWDuC0ntA68lJ2sdv6PP1D6QMjG+xrAeEpi
P7MMg1cT7R5v+GY8kHF7X2R3KZ50KTlwxkd6/3WkrIrn6x4WcGVi3OG/bJp/1wmA
3d94avX/CrhjC666PxAWBSnOOw85XsogIY2KdT95koB8lKC6CInU51DVt/w8aKn0
+6RAXmLVV00ZU9RwOlmKVVllWZ5ww2U5F9FOUfpOgs8Vk7AxEx6sZxid7inE53+G
rcaVvOMoTT8Y09CYp5ZN4p6koWObA0BS44f1d6/h9FS3upnAJ4BhdIusGXICwcPF
uvJB9K6y8fMRZiqyFUEFP3YBa/hgrUC4LMGBM6hht2mh7mKIV6k0+SgWykDlSn3U
vSnMY3lJvJhLuOnUNUaAAU3sWQQCPeVwdxQFmO+GmSElDp+WiHVbr6EbYZjVbWuX
Y4xHy/ictXy6rfaXJQGTPSXHn5lG5wGsl49fc4/b8BJlkDhThvpkR/GjpEzy96/f
lxCtbF8edMwhadUDFd7Wz23cNcR8RG45zoMpUJ1rYuah+RUiUGjE4FJGvuvWMHSl
ohywCGjuyKCRB3s7WX90KgSXzgLgQ13NGLp9vbQRscMlbiVz3OVP0RGWgNiO4YOt
YnXzd1f57Ki7S7lP4zi4zCoJgM5tXLJF4W3FgRGSGiHQMe9C9EIdHSEFAIeCMoLS
seMavDdBRv/0LxErJZELnNGAKJd7DNGRQGyskZF7nD0rg+HDJnCStWywfu4NvoMJ
r1+rLooyZCM9uDbe4syzMidXBN1rW3F70AijhRho2Uczkb+12KEDk4HyB4vV/hr8
J+7sARGA/UQ+MRkZPhFI4nR7GBtiLFokiHf1E1+nMmscI46y69/tRlS9cdhw9an2
sbg+YkxDHLBpyy9/nbRYBx6icJiyDLQOuovwI6DZ9BapBkIMjw5UR2rXUr8PP80J
qe2FfSLtUnla0HZ/2BpBVfduNhOCEfsQOUqDskUVliZrSk8XMMyv3b4IM9fJjgKR
wPPcsy97o1dXgaVWxj5YJJ6oF6bu5hWCd/vcqu50PVw5oQrj8/rooy1T9lxljJv2
ph+jvmruuEH/T6WiXaYf65TYuJRPux4sA4yVQMicMicr9tjB8hNYDRnfy1B311Ta
9VO1Ra95U1TSIAInQvO1FUFcJUiQQ1UPQmS84J3FKAxfHJYaOQdC8JhUj8WBBv0V
TnEXpejs0gD/2lzE7g4lD7DzTqJd6MGfrL0bONfTZZKUEdUqnHkYjrm+XGWO6REs
rsaFvsxhH41L1joiYoFp1tz6LcV3uv6z9ioolSKJUT6OgLirQrESNV5a4oo9qr38
1MNG7i51rzmQ7O3Ma1Bxs2uDm7VoIHTAWc2UC2jmfI4Grv09yZ/t+XPrhvjBeB5U
F8hwmVS4L+55hO31AQsrw493pYLqm0fMve0YGVaOViJClpWBgGMbZw/BUjGdkJyF
qGsvtr57HwluhbDx4jpgr4XycvLW/dT2PvESEI84gxmgrJGAg+UjvHdntk7p1JU4
RCG8QDsP8nZbL+f3R6FAZIllDSIJghpBefk3lNefaA3Uh8fIZ1M/5xegSwMxyH+E
bxdpGUuY8D+n7iLI3tKxDcI9aorlZunvpysIc2pOwCYhUK6TcEhGMOHrcz9C1nS3
GGewSOlA3EXLhtDuNhVwLmK8mjLrP2/OXbBtKivFuW/If/6EAuX80g6EPm1+WKoD
Vs3rzJXAVt0qyIWNUyUKtUKsiLfM7cn6ZXvBc92ydcDEMbQI9aSQvN/o5sePSOVq
GtWN+T2sITmVPAkEtpWqosuJStwKyVwT2r+OxEPYLSpCbf4zzH2yG3zFwcBKE0xz
PRiv91LBhLaYnimeSXFkNFazf0YRQ4cR2pQ1ngy9BuhM8ST1F/B3sPcPrawLiK56
uI0vyoWAB1eFEw26gQ4N/mAyctN+XZqbM9xocurcFzp1tDxPNxYoZCjlBbk7uSO3
IU3Hh8tfZv/kAV2j+GwSxRfzZ/mEfg//PmzPKl7eqIgyIkFmAptRTwWKpJblhYDj
lBVTRVsJlFvj3BTe9uQ70faByoz2ZUMzfU869lynAe4jR/tKrlTIxOTR+PiT8tp6
DAgy+Z/qmorqMX6qx8g/fDcW7AraRgQqIK+qvnwCNtYTEtKhrva9kgqpiyu7NlDu
4Or12Tj508tGFuauy/aN6BVi8Go4b/cf+GCeeNP2weHATNJmj2u85dV1uBlEZzw8
72PEjnGxed7bBboq/2MLNAnQ7vadidqlth78sV2h0Cf8uKyYd/AbzoygqtZZiF/B
yzn7nTOA+ZPcFLbWRcKlzT2ZUCTUtMUTlA0LpG6fNkseqGAwt4osjL9Jo/jZK4WZ
5o7af+ThTOYFxhCjzooIlFhcL1ka1HV97fbL+ltVaTXtaqdsFv8iZ9GGq9vlG+Ed
xZqHXLg7VT0+qjWuM9MKxrTPxhpsi962UfZC5rufw+w3iNMQ51NcJWaTNe0NZ6Un
HnsSRl9uE4TweQc33zrbbf6TuPekxiqpSKfK717CtBRR1h2gDzfp6hIAEyRco6nk
dpVXUvc6RUFZ2qs2bRwXQ/IliDE1HfKva7kXe65rwoUT5lfymTXvjkEeSMWQgMQn
TOVvUWkLHX9VfVlQ1VJiM7zfXq4I3N5pjBwgQhG2TlSo3Gh9O60Tl7Ugxtaf19KQ
suDmyNu6AspBiihQ1LHvAqBBR19vT/cWyIOP7yiHRWRHxcfnvAeYy9GBFrNNaToX
bp1W8LYq3jMbeFXtKAxCIpQc6spypWFZdvwHm+Q5BA20hBTyHOJlo3eFpS79kHnx
IQJafIXFUDYGiFzKZWUknBMbvhdL4q39ufoSisKrG1M2HxFkIf6xSGuchvOtuiIy
Kph9kFvetxdvnOyIe0OEy8ocsepJOxVBKNmpSm5RNpDWRHnxfYQ5ys8J0j9OnCQP
+NMtu0P4CG5NROe2pCBS2FjZtYbLZjJLSr4u7pT38jCny+MqByZXgL9+Lynp9DYe
5FMAQEMPT3r6/+h27bZZlDF9yMHciZcM0CMztBosp06LsTbs5sroq7N2lVFIoPMF
o8PZv9g/7VBxIMaw/ws/W3TQyzUuaZ064PEypEZfz7gxqtFgtfHB0wrGYwOHtQWg
OKJCHNrUbJeKnytsG+zzyjWtkSXyP+Kk+6SS4EPrglJMUQIdapbeGR55UfU4F6Zm
PBPaFxEB0sgLfdSFnaUFF+JAj3MpTi+3fCU8n55Pj13cxu/SJA2MkW1OhM+xvdWn
XX46OiNnaEswwoVFrzYkLLLj+a+7t5UIgOXclIQ+ex+OBMRK3LF13GZmnkQ2IwOn
3THy+k+k/0JyUtc3wB9yFGYV/rRLy300OMe7GLSmF5nw27w3cOGaNQA30hfY+n4K
EBoXgVFU+BUYau23c0gU3zQXnwMJJZxGZtMyLelKV0DJd4t6nRZi8QwxvGl2MmLo
OEuXNQ+caPTd5BPPWbDcee57kJrxG0UEYvxDk+KrubBkuTE+QzallMkyQp64Cl7l
Y98Hu1C7pjkckL86SmcrGmx/X2jqT2aeApBxLOBggT5jfCIrqEmBp+y7xL6or54F
IRyp6tsocWUoy8Mlszf7sJRVgHNNCNeKP3mqX6TkuQZMlmu2dis6aLmm3JNz5mEG
sfSjANIrv9jMLdySy0MeSnR77uK2yAZ7E5BFcqTfHDhokTaDd0bLuxP/4Q0vdCZW
fvpuR/3H344SLq7mg88oZC8/LU70McCe5qbdnQ3/rzSe1x6MIggG1Gb6TvuYVvVD
pgk9VkqLYHyc0iUyiZffLLf2VXZOZ+tg3hOlqRhyOWR7+hRXMzMHHPPPHh1DWDjC
DLB0lThMljGcHdjeONFT5H24tzNLihJ/iRQiLFW9BFrfPSScXNG+URBFmI/CHROS
QorxAyNawtetPTcQzLePbpl58Bsa7wywi0NiKSJ3wUEUJeBl8mmRnL4JvO2LbEp1
P2r0AaUSQtM/WbTN5CV2HCoYBWvsSBJ9Rgh5EwLnHBRbQihDEAA4sOz6hVyfcThY
E3NzexU7ZhJ6+z2bZwfR7QrX/zoDQl6BGmFjNnkdtPVrUOgGo/ljDYGuGDSTSC/1
8hm910LDieApZ0zikmPyYLHGrntzhji1jeo57njeW/mXloGvS1wzkZk9jwSf6vtR
LHVeGZ3cZaGDZ5Pae42unXQgGBNq2Tx86bsyKLvl4BRYGlBUlweuJOrPFBeIuqHz
MH2Xh3HzvU9ZS688uYoYhDMKl54sVlFRZnVcrHddgt0AL+PMCGcoaquoeEh+Es5h
/8efvn5oJjB5snUvwhgYE+z7568McF7J1doPCej2K57WcbpofjwnPTybjkFgtSDj
cRSKytUS8Pjy0litOUwdDZkDvT0t2MAQrG53fRUEWeG96B5zf6c8mQ5HADVCwdUN
ztEZpT+Ht38KWixr9RaieFwPQEnImhzMUUvR6zH0HvQxFfUXEUBk25LG+zLwiUe/
psCnsyCRNUycOC+lSmZJ62peFYgqMTkQGiNUr1eC9oH7qB0Bz2iHSH8WreQV1ROE
NKeHiaM3naHfgGDseZ7E3ipkgNaxTpkqYc03RF+VqwWv9UkfbT3sKP6vAoMBlfvF
F4HQir04Hw37JQUdJ0qx8vYLTXu8n8PSpPLG3buPDJ+AJO16JScDMCDIXpovehEG
zOQpKo92/qaua5BJc3URY99tgcJxqAP+LQY3pd/IxURaY61zsgjNs0EQhQr5jp/A
MZdxL9gySO96NuL5XtP5oX2sc3SjEz83pFvsW1zYBvicUh0pVuz91/lT73AB/DmX
7yhE3b5k4Z8kvQjykGW/zWJq7zswQ8hqI3OoYiAdhqgcWyBCmJ5L9H5CPthDnvvH
OYLlYr9g/m9pzJHs+C5aYKo7DS9NLz4gO7QxWtbsbMxNMiPrZql7Azw44NPqsMhf
kp1e3BsmaDpLzj3PZbhVHM1Y67hDCYkbVBOb5hLscWTDk3mcycU5zzMeHQkXPSdu
wUL6bxhM53wU5uza8P3a46wW26Qb2stM1gvMnd/vn7bN8Z+hHEHAaMXXChxpKfW7
AiZlHh6YYSRIZNsmQHZvDk7B0IRPP7vdFEJOMs4VTq966kwC+FXaEbCDlvcHpdjR
ipyO7ktuivPhXpMJFHEAdOYBgRQPsvyOPzMnAqrjwAj5gzwGqsVriVQgfDr22GHZ
l3UvGWxY9VKnFVwyxlVI+znvxZAmKQmMg/I4ZcH+4vHn8W1YlzE5jX36oyNQggIv
WKr/8hO31ALo029PLotx6ceWbTn9JSZ+s6npXDwOzBgGfhEqySQqU0R/6qJypUJC
T+pHtWRt8j5f5rkR4QLBqZoewzQ105CVlFGG/lCRpKab+7KXf6OeIS2a40WuewhG
gFKwJ1yCpU1mszVt1iyt7arQ4B7sRhJbfFNNJAmFUh0RCJnx6SinyAzPTYdM2D1E
83mYWNRQwKko1mv/ehoXQz8QMGSTdUi67zHunmjNjat313fScNY/yC2BoH80NRWv
etm6S8GPpjZWrv6kA+RhL5fP+h699J2eeoTJub+Y8OP7uGshkaIMy/BrL+HIU+QE
tZWn8gx5XEggNO+8VYpvx9nxcxYRDnbb4VKnPKUQkYbHDdgiJGDgKNJqJb3ktm36
C5iQOk8MTCSVo6+E3ZYqDIee0KIYHmSTMaW3EySgL87afakFdupp1X7lQ998Zexg
BsWWMqkZpaAaNbf8eh4I4Uf01P8LWANgcnZAciDzoJ0v7FPNdrAzkc5vy0+3hlFK
KCICIfdH1th0UpVhuA+YQLmK0wh4qP4w/MiTBkxJmAsgDd+J4TKO80lTk/rNvfZZ
MyA8G1n5xT/kgzQI8Hn+peMJYZJTREhGvNupvAUG7LkehKFhk5BsPtZ4tpOEAgJh
m0QnFVM4wq2kc6hHM6rllPgKOJwK3/ywzSKv5APpy++9nVGY3e8Cj9lJJ8SXEHJN
SM4ebq6gXRvpRUiKBhIYehWIQjJixSfN4XxtSxTnWJdp1iBBNkXO9G8QpY1UFnwh
iDcdusSW8W665oc0Ck/m1DX/CmtfEo45q8EFlZzNr6JdRsY5ssN+AgTVxB8RiGvK
JUMjjw3OsVDLbNzgJocd1zK9Ax2FpENQK4hkDdeIfry/QYLNvaRSXbGsejnIAyy/
Iu6Byq4KLU39E6Ac+B7O7D5Qq1+OxuHjsJCt8cB3P2OJXm6ucrfZbbOPL86Ba+bl
JagUXW6eCbMBel3WLKY+WmBMf1CFc6dhAD03un79qlwRAZtdaQZx5zsHnT3z7vmH
T3IySAiFhmKmPQYLuBNs7GAYsIkSNeYTBbnH2wjY580LvvmvbS3pw7mOjr9Ezkal
tOzbQRCBn5Dh7HT7oEx0BHeNWr/81vZ7I5Qr52LeCiIY3K7Vjiax711FvLx3n2jK
bs4hTV7ztLK6m/P6lOEgrdyXIIiUmkBY6QTbka0A0zyKQsQ7wHxNKU/FDgPPcWCg
FzET3Jd560sB4C+BzJ0AeoWXFgwjHiSuyD5yTiM8vFXJL5NcO5m6+2dvqkp2KntA
zB1IM65TNxnrN9rfMh6YZPkU+XgU5bqAYb984qILOqVwDKLUyG6Ajw7T+VRet+cr
2dC//zPFdGwChAvlOHY1q/OMP9jrZu7+7kBHYEW9/AX4IotnJK8R6HpHoNIx6jwm
vKR5MIG8aYN1LlUlI2bz8nW25DUEOcVkMAs7Gphx6b2eT9ksaahJkjPtoQsV7zic
c0fmf1s5jboB7cl1oPNXkzWx9qif4oZlDpvj6jijR42+I5Puk/OBCMFYV/hTMKRs
stXDPrt4o0NdJmKy+o4Suhz8+LIy7h2EM7G6gb7uFZ5v4mj5KcFDsB5wPJ+FN3Lj
F54RYQos0ZsQYCp3RmUr+hk9tbxN8upsNc7ZWhpyFYR86O6XqSbHOX/pKZFF2vH5
de7hsHKj7Gv8PMXoW5cpKFG8MmAJLcCdKAKdDeFAwc7y4vkX1MzAUS0sNZoTnaf8
DIOXQ2GxLMQ9nuj4e0Kc7I6TtM+p1wT5Fv3reBcHFjWx9gmsXWdw7nwFEX1QALPH
vEanj5ulDC3wEgPqDnKyJ8BdMwyUw7g0xys8+e952x76QWWYtni2AIvBi7ImrcOk
byrnUwQwwzHRzjzRy7Rc3H3MrvcP8a1xo2sZEdWLw48Mi0LiMPnsKK04MXAcMp5k
pfCxYAK/Hb/ztdFfZi1y4krnXDpvvoAkh0HZ0OnYr6hwPzzCs87tIMSE9O8qhWQn
lXM9M4o5dOMJXavrgjFVAqgGP2k/ILLsiY7jxCDrHMK0WRx3XUPBou18DVydIJUv
sLCpQivlW7zjWEI2KmvbH1O/z4wq+fof8w21TdJuJJQZA09MXf/PyIDnteZzwwGc
fjpRLBhwdpqLRCKPtKvLcZIXeJByHkPHOotTXw9XJYkmYvbI+nVZoeQOybloivR2
dXfomsk6FyFoxmyOxaVEZz7TJiiEloVrHTa+Q9CHZKiiM345ISo/HgonIiU0sxBb
182iPb1xFP/PpGErFSjF0d7GAY7jwfwbF+DjgrLVeRpqsIy5MsYOFes/h9qoMFhn
2MeOSXNzZYWHoVSXBD7L4Bsd97phxQka875Y73fDFeV5tRVwaqpelxMtEdti7T5M
cy/IT18CpMtrCCp7sOUkjr4FSm+IivCVQr0iAZ68bSk3/DCjRa37HvUK+4lfoIlx
gT6xujvZCDX4eNbpPgoA/Uew+F8aTkManPpPTRsseTVGVJR+aM9LUU860kOuJV5d
YYSYl+QgEGO70mXQ/M0HNFw6qob0dSu6ngqwqRGoo1B6hhG05eTbE1q1uiXc1ncW
uY0WtGVRalx1Mzt/7WaxXnqIhYG+P5b4HVi6PyA69BgVLrLvRdRt9V/QobVGEAmd
96ZlO4KyhcZr0Lk9CYoibP18kNaRnD2cnmGSYwtVGalO4MuNhOz0zw0C9S7KpNyT
0fL7JPxkmODBMDQE5apjTMUYGoAm5+uydPOGG9V0kPPulBe9bGgZ8eHbVg9bEnnH
siAtcV0pkOK1hYyIJ6c0FgHoDfxnh2+na4DQHBSKeZq3IXydqfd0DbI4OE28nx5g
piSpb7QuxEc4Jy9XBfugQeJiarpXEcNcYKrFX53W5/KLaR2yDAqdn6gDBihuV6Bv
RfuHEN6PcXqyocI3s68Ydb65sZ56xYGlsnCE3pAK1+hlymC4kGouAXNo4Ge/6Cmz
p2udkeYOzdIFPZVo7woEqUowr12Fgk+UjcJ7Q7VetAcyNb3BWZNa/EeKTYSrYymY
Pee1imsOCVBdpVQk+NmE+RHHGGuUV1eyEK0xyZCrB0x9gG8qkHRBPRXgKXs3HzVc
1Z25rk5/iY6NZamdGg+ijbUWNmMfXZcW4HvIKmvbEOOpXg1L9CpFdIFy6IAWW21O
XYV5fcWXdu2KIZRUfFudQpCAVJ/UCngb4gZT7ehpJGLyAcPHC9arLi4/YXF+BeN7
UjlM9Y4TCltBLHkmKhWQE0NnD6QiMYSNGOD47tuPBgsWr2uhM7rZcfpuEqA4qJVU
wZ14qpOWaCF318L/0Gcj3D83wOdH23mW+k+WK9yPFkRNqM06Zyu2DNG9o0XuA4ww
KaOtIQpnV7b3XhSodmvhNM7qpS8zJEbsIforMrqgDmRlMupFUqUOg+lwKz9c5JhL
tK+qQKMAMTAi22dewUmOyIjGx8Z+ku+oc/c36HNHuP0UnhKpMwTe3aubFsHPyJZY
x+cjGgKw8pAusUYzhLHWJG+jN93Z2Lfl6daqZKzx+netvAfCEgOQel6iJC7aPk8j
F++IImIpoNr5rC04HP5JknIRaBQKK8n/MOuTPk1mTKZ8HkZsJOAZXfShqBBB2Th1
vWRaEy4pWJfXbSgXMf3VL19B9cX9BMOZFY092JFumgaWdT3e4IG1KCobYtP+hwt6
lxGLGuoVYCoi8S5DgZtwG9jrrkMq6dgiMw/BRlGAo5P1uoszC+1Q+lBrUv8plojI
zcz4yZFjRTMRUtqghETvp1C88D/c5imIbFEL6rvoQllgtBnCBgJAS5Rzg1KsBOlS
zw8mrCg/S/xRG9LFQnntNQ12hyOryXW/jPwI4Wdj1wTdyYJgr7YILUKfrYgt/8bn
xRUhoMcDs6Sfb6iFFHdXjEs7RXoNBVLgeW2Qwjwoff7Noevl8mUxvFHFcnzgJjvX
mY6uxpNOwKk5y7V/I+wd7sho+bK3yswaq6j4gWnn5tjv4T8JULJv/D9g2WZehjzv
jLWcLLL/ns+UK0n432lj9j8258TZseWBjhU3DQZKs9m53ow11h8GEzD6QCJP0kfB
tZDKkDiLzXFDHK4u/J+a5KoBWcEwDlQyVR0X0PrfyrU5yVidljpYhJde3BMQlhEu
SsGHpFsxAxgZiubNMcGKMBEATM4hfx82ISnqeHobtDxh25iDfP7FhDXK0jH4YcJI
6Sjc0aoyoGY+NmEdhYal6eYtz90cWS2c9np7zUDOZKQzsjr+FIgigPHi4V81Qik0
dwZlPRZG1K4mG4Bn1RRW8Bowed5tue2tlw9DioMRo1y6SPc6MYFJ/XwfR5aeZZ1l
LnrCfScDWRhJKH+ded+PR4fjjp8h2BaKE0HxKXH9wokdRE0Va0ojelATu+biugR2
lI15ihy8dicJNNP+MlxRlMnfY0ts/x42zwNewPFr0x2Q1NGlUBm62Zb7KvQo9AwO
DZmNCn4C/mI3UF41GjTZbET/tJxlDq0GWN3vwEj3vKjfy6ZLlKUOPfGeqtLhHSRk
o9AyEvWFA/EVAm46xXT6FFjs2ZFlYSIRBnt7dS+xErVJYPlu9v+eaPpYo/NnbcC1
fV9aveHq75Hx8mzuqF7QWWaRK/5LRcKzqEb9x4r2h0aP/wKrs+rN6eKnvRtYNo56
9uxvavxIP2dV1yE7+/qa60lXZG1v+PQL5Lcur2PPzTzly5kGv6MP/7ZdkI+HE0Kl
E5zFPyQX2V/m61wvvxK0/fZGtIQzJ+oJJTFHjacgJWCQQrfvojcsCyAi+o2BOKqY
pHqevR/y3HUR0PionQ3eFxWAUi9TSxJFvluNPOqzNh+vFnyjI9bwQBhkHPoCjGv2
xDs56U/ChTNOuQPPwgc9MU34YYc/WIvLmoAxiLTKIi+9nrunQpLWJ0d1bBBGvptC
8UOV8VWeNbYmd3rmvDNMi3PKulaE+dzreRZpXobscC6cnCZxILJNzmrC0zRGzQF5
TofyRDi9jFW2DOg8fgu4unN2gQG9KpgxZ81oF7sfma3XY0rbUo8uZ+WN9JPxLJ96
oS2ObFpHaPXTD1CD5d7S7A5Nzy9irFIyhqV5ij6gH1NSUSyAmnMe5LjzsXuS6TBb
daiIE4xaaXVi7S1JODbc75nhtxMTp4EVxxJwEpaW+2mAUg5IVrkRxR07vo2n1O5J
HlYuUWqLMgbG9712CFRAMP2m5zaNA1fXg8i3tDHRdCCZ1z1xWdZrACOionmuoxhr
PMRpOM6apAg4IbS4bXDiOUHE1vlcoJzadduhiggFp9NlyDkNgADfmKSYKEeHk7U0
8Rs/KFyvpglrC9R4gzaoyvH/3l2i3vpTbsxCF4hPPjaH100ZfXNgL7O3/9bNxyDS
wepwAjT2bHQy8Vfo7+lDbLuRmD73V8bAbEwCzOV84VGIdyL9AC/RB8omzYENxCUg
917SdWZ/oftfGshv9AXPrptFl9FjbEiG1Yx73z1+7A8mtCt7TGfpzvF+PqQjSHCa
ilDuHxos2ojlzzkU+ZiwWZtMLASLkvGvbAj1pS3nCkMDc9EAkbElnuCWkLpJpReb
0TKtIWqVMYSxOXBlHL3yTohk+Y9kiQ+ZA8mIh1aWPoXWAVRC+w1OrLSj3TO7/WlQ
ocaIBl5jJn+gYJuV88nJ9Ir5WwSU3RZn3ivvUq/tBNaV49vsSo+ly09ERgSYJybv
w1vhS6lnquXnikaPvXZj+AdzX6qsgYvGL2wMtDXMH/cPBhlsfZo9AkaAiCd+/J10
1ShkCK8JGiTRb7rssHMRY/1JZdd9qFDOS2RHG0Tyc66sC0iDX5Tn2d+GjecDP3LV
DaxBncXbmLgI3vzWRkMBJ3Ulr8sfold+VCo0beKSYygx1z0V/YqiycinQ5pgAPgh
HHSVlj70Ciaeh5kQkW2Yv+pKKofHp0dfG2jlQkJXE5ZWomi71ffkWwifHuw/wgTk
UoCxIwiB1OHYKbMFQHTMlc3/IUmaq39KwPW/r1wNEf+1doGXuqeFDB+vtHWJ7gR0
fthvCVYT15RvMbZ2ZIyLzwUsGtceMRz8lNHrGMWJTpEVKg9U9ZnryceMYVo0Obx2
n9I58VF4lWGJpL1NjeJbuXc3xCpYrhz4G6OeNKXznuJVB1Y4oPYnczpmGSkj5xbN
NUEPzM8DcvzB7y7BRIsIce0G5xYoufUCT2gYNenlPYrXLxR4U1s55lv/hl8ZyODe
JS3ni+rGcETQSKPfPhLKTHgK2R+i3JutyUiqQL6SacsLxDPZm/GtqtqeUBS1LxF9
3dv0t0zNTfjySFC5lAX29qBjIhsImuJ+CKwtDSApF94Enk0JXlArOpksINJv8xmf
m53CAFDmToN2mKPwme59VaxuxAG7oOXtZOenlJNAV9T4258ujnYFWHoZTI57RjUe
DZ1t0k607vCg3Od4naO+axUays3uop3fI283Rha6qXc5D0BqsyRNAxke1Nb53KkB
q5JPIYgHWTQtOS6KfIaoPY/SBNcLY9x6Pp0l2moFa65oxOTCxoai7Q/2l/tZaaZG
TbgV9w2urgxm4v2OqkzofKf7OaFcET4Zbh8mWHr2de+EvQFUcdU5dTyaCQSBsPKu
G7PNtLmoeK3e+AkPPbmSZHPanvmFvVVGiLUCEvmWOHLLJRVZHvsJLzetE1zV8pmr
tq7H+eevPSRAfz4EXorq2LE8J7fmLk5kqIiymRDnXtn3xTnFEVe+nhxRUjVAGt+f
DpCJ0DbbhXvzNcwtxWQk4RVnFbjVo4csfH/QFQv7E0LANdsNS/xcdJNJ/kLd5o9N
TO3AfVD+5x5utmBIZMQuzHNP0MzkTSXPOGGl+Q1USMnyo+53oNNH5Z+6feg8/gRK
B2lm4bR6D9yMOLNM5Uf5hi0F5PZnIh+uqLTdFvJkPqxkgosbEgDPqqB+QiaQLEWs
J08Ya6YXjogK4lzG8sRY/boJcaYzkHx/BiB36ooM3KcWERFFz+yeguJHF36YfHUX
2d3wB/gSzmWNrmPxV6TpdUlhc/3p2X3DyM6ZkCdklpKJv2zou5zeqV1oDhTWbiHU
WlvhILX5N9sL71ywwnIdSVfHe1B7Hm0+hwigci+jk5lenjtB0Q5gHssNGNCctg2O
iieJHfh+yr7CZj2VuS8CxChRqfGBIH4i+Hk+lMF4Ejwt027M2/St4XXJZt5wtdYr
uE1xGeXY0RazksanJhLFcfwxNReSxbGYeQV0CTCptnGCoQtwanyPERr7H+y3k499
4X+VTtwDp9uhNUCKJsDTBoVhBaVhFuDkDdk1fTvTDcHr3RKKmkpEmWRb+DNnYu34
ee/pvFQzl8ZtSpJjZir+FPrT7legtk2wtBYn9YoVZY/9/qQZjE6tsLIVsFXc8yA3
jU0weKUESsbZorHM0tqYVIDdW/LlH49o1Xt3TJ1KLpt3wzcq/kQybmvJjjUEW7Gw
4hCvCsZyccYK4Q+HKFPdHeeAniccwLV4d1hQOXxVoyxDGyPVgBY1PfrX3gbfeFj1
K2poAeizjZFre333huMTkPPRDNADbsC6pZr/iWK2z5yoQmB+wPtm4mw6EJtHbiSc
wa55ppna79Ncp5SYnVL+b4d7rRPrk++nucwvKr/SN8VOT01NSoq9S/9JYInpSBTi
+NFrDY4D+mgRhCVSiEUwL6pIyO7YAxa/ItJE/EOJsgB8UKONCenz4PB6ErgIa8no
LvTpFZ0uFWm7tLws3K8ByX6JtQZnBR6SR6iAnXo4Qm3bdL8ww4q3WRfh7JZUZIHA
1FeT/dBBqrN22T/ElXoEjbYSSeFtkydw/lXCEzRmHsTtlSqdOva9pRRT9oLxeJ1H
Q2F6j+SJuLoJwqUf7I1DfjB6uPtav5pGa4UyPVgkDB4yI61nug997MXZo4RdRWAs
uCaveSt46C79Up+D9NHDLYWHj/7Fm20/L6iut8aDnXHf2oP3da/6uRBA9Rn9hg5Q
jAiVJmE1iCwp0xnyqVKR0WGcnRBTBelbMNWYTfjpZoBP1ptDBT0HQSY4Z09lALzo
7I8JqDkvQtdt7NgvoShMCDrhuTdoGSD9hovo+kA7NNSn/9baLWvVkPnql2eeCjJv
6GwLlMykOqPMTiooWU8Bl7qGePqlQLXzXkS1TnRB/mdC98USwHJIvDT2TKgkyS4L
hRx2DcJeh1PcESuMjAQshht0Kgy1n1FGtF1c0HwsGYgnQzQHBduYIJinE6Z/Ot6P
sZ+TZJyINcqvY9d8W2g7lv3otspVMwE79zlaitRF37027vS3YohyYTgmJg65QYWP
iqWNWX9KYKiuqxiIYd2xr0FYWGWX07Tfk+Qp72oIVinkqdZAx0uellJ6+JHLEUvF
tKYHSHq+zlKPjI9vsEPSd6UzoqQ8YzbFv73W7YGJEdtCAfBCbwkXQeT79rOsKvU6
e5WFWAleHFkYqoRz6yHfwxU6/tcTAjIEdPMCqhFYkyfNV4Ro8zrfyn+Rq7nto5rS
GukBIaBuhmlIVBobtbn0AQCU9HqFJ2JGmdedx8c8PAJZO71W6l9CHn54TtMNa8vy
DTPsLDjc6KaXYU3DgDJuaMiU7tq+Q5K7yhDwDBc+SbWeGZ+hcWr+mH1VUWqvZAKI
ay3JczzfeFuJCTkCwAZbXTW9u130CVplQcUHreF7zh6/MW/PPoGXM38sgtkLvyq8
lb1GYYWXoYOOGiyBsA4wyViEyYEiamiiSm1iUrI8t+X2EfFaFMPjIV9Pu0Izjv3H
vsrGqMVJshjSA+U6JTfnmXjX9VHJPeBvwBSgviR1SSRkovLCs2luqio57umeci0/
ZWKKj7mbPCDqyqQVWg1D9+7cU2/kw4ASLJ6InRfhyiQm95FG9ABy83JYb5Wf3isW
gOfjWn/4Rcc56w+wjqkogkUQTzrg5lOwE/Efgb/SASgdKc/YEDB97HRe/4vTlin+
7Gpd7h0YeJCQp0X1SUWmK3tOMDnwmfxFkCvO/YYFsYixatKx25EM8qT9/z0uAxNN
f4pm56+ibr1CPIveznqtXNqvREEJ6ruTsfycOeIie5jYl1K4tEjIJRnhEygqKnS2
QEuSSwotz8G+DFcdW1+4ye3nMNmpqqHJMxQFScdnq5p85MwpOkz+t+r6KWvLJjvj
uwbhQHq+yhkcpdCsgH0lVtcDafIr+D+DkfKjnqMO0RmdPDgiBsIiALXH9TpyPRgL
RJhkPhf95FUyu1UokM9tjDtZ8xopj1KsNgYEZ8VijsY32FXQq/inteySmQn24ozv
j11Df+ZUBXm+ueQlvnIcI20z0rNxCeJFQLrkJ8xsaczAMGln1l3uN/5wW606XU3c
5tCQ6ZxV7vLdtyjEBNb9O7im3pOVXM0h4P8mZiyhzbRaJfepzjoPkwxiJUmwZsqa
Q/03DEZhbwxeKAn/ROXxb+/rzSKshAJhclbXYcmFadzeVdPK4qn6rGrL9I1Y0COF
zQPYEGo8xu5ozMdUzUiKSyGXAsVF7ID1V6sS9xgsfGN7+q3wfufchQuINfNObemS
Xx9fOE8JFFfzM85psPhoz2RlpMO+9HfVISiqxmb/9ghuypH8Ln4Ihml6cjCnog8B
029LfZV3mqJO81N37PFCirEjArYYnWGuV1xVBsvuPaqms6dOA+ShKXAW3UjjJUR8
cPP2sw5yZ5zV+taT2XHVfk4tenEhnk+weCe54nBk+sTo20/aqQM5IRd7U4XoEEdM
VoKV4FGNwBn0O1qz9WqrE5hNPu+zY1o9fIFBssg4fn4OFdtRbBqpc+douRUTwbac
sau+9PGBwIWu0Sa3al+mXbyFJbbFfPJQkRYcKUns5SvuaUmMCuGaitnzY7ylEIfU
HEe2skz+19LgujBF6cW8/TI+tIvmH5A/NWtwyYmsLbXX2FSPTXA8R8WXOVgbsIRm
1DE0a8+XCekILxoYcE9TaSwN4PujT9bTQPfyYzg6i0Fh/zN4TH9YF6TiQu4bJKre
jdoIaZhr2gnuW1JxlMZXjtrGiUFVCWwSJRHXQZsmkF2LklWCMV6qom/KWfc/cuOT
/gmn93YHw8rJ8wRqgsTYKqjjqfYCbcxlR3qq7DzuwNj2HxK81cdYwiUfQCEwX1h6
4CtLkrH0OoKaNbBanGBrzAHSTmAN2B+FSVg/PwEs692fdOkHGKt6YStRO3ws4zwn
EzTemWCdIpHxa/QhKIQ3KrAKCgjGwtji/AOj9nQo+ifgGfEG3T5CebHkkeIR5dxA
9EZyEErFOwto6Nh5miGFDv3QFJWepsq4ybFPgB7W25sa1u7p+MkplfCqg3pMdtHf
leeLWvRdbYIGuJCT3VCyP3SWK8bifVEjsOo0MXe9jPDJP7CeH3VaK0nZGSOfOPEB
zD+5jggwmyjiE5PJYl0H/f0E78iifFiXmhMouNpSSsFwtNAiMP8Mjzn1wyeP4OXv
tzUonFJKF2ZqLHCJficnXQ5I5NmcjIKdXpJU6rtu7elADl0BCdtULPEQyrvj4L4H
j0U6RckS6Q4mJrLSQ6g0KZVhLF00lSyddNEHNoXCx0Bg7JAG2LyEOTfFZmrXo9kM
0oUQQ9SYJQbaOgeuJalshW7nSRkCmAND6hvELdN5mwerOuM1F9o8G+3Dv4+6CnTP
DB5xJiWLuC4Ii626EHScRJv/KCldEUfTbRkfedeiFgYBS12nE+XdpmWMXQ95FfCV
IwNi4ETHM9uVhH7jmM5BthARA1DF7uOu977pdG2ssLtkoaEHOWGVXpx6ykEaXl54
cyHRtc4zg2+zLXLIoqHi1/UouJagKApXbkKrTAVfqG570GwwrAadqG5rUGl+bV4M
1IpBQrznLOBdQP2/czfDfqwS726DG3J+RtV9ZTN8c5kQgPcQE1zLdTGiTZRlWAwR
wbYyDbzOBwtglFUk8Gf7xBGGfFlilXRMvB8CyYMIC6fhvr1k4ZYDMfGQyIuwwakE
vW3A0quUUgsa8yMUJcTydfiiYqoadk7RMAg1ODYXitnw6W4L9EyFdPX/TojvY1Ip
qWx2Axx//B/yam5PP+3XSb+ANtMRypirHTqDLOhKsG2muDf1/lh62Xj6YU8JyQ9f
edNd0jFzcCYsjgKPIJKl+5/tKKoqh2WCEQwQ6I59qKfvwdz07ZZP5F9YAvj3kDXw
0YWHH7+y8m/fH0DUdXBAyH4w0Rm27DTLqx0Ao/DQL9OJGjLx5CHoj9JNNvDbr3d0
We17vxuVLu4R7zlnKwqVUqHdj2NtEFbKpTguvlA0EjDnbSuNKpolWBe5ghLAH7kc
DE4xEV0uwSo4mUfm0x3h+iMvxoVSNZYfAROSm8ovEsx7fElUO4N4CYah30z7zoS4
woU17MINe/UojrFdWuAnV6I9E5/6aGQNVkQqh1/yctBS0USJdySM6t01t/XzWw6+
W/2rrQ/BP9l6jRg9wCXVs8y8MIyCHkdKiS1OPT8PIDUrcq69Wxi0EDXSfhCaZOqq
+1mWDJIpeoeqxTzg5cQAomeFS91K6cdIbnVmOzAFVkSgu0m/YpKLo96LMiqgDA3b
f+sk/huSd99irioYTBkezJ/xxly4UTiEuA01vziGHPwYa7k01GgeB467ZxVI+UsV
4p09JjUEjccYlgWQNXC2gnW8SQEMyG7TkWRZMQ+M1mJlD38ExpQYKm+GkHPcUKBX
dinLzhL7oT0WpyLkWC3AXfvcHd0l46lLlbTi/cHgUJ4QNAKLHh+ineRK7nh7kOtx
5deU27WlZoLwYwC+Xc4u7tJ1oMgjbZmINw8pFE4Aw7W0wOjorOMcRhFvcOONJF1t
nnbwBM+hT2CopXPyoPuppxSzuPL0gJsDG7O5m4QrDpnNt8x7e2fmg8xRlbifg9FT
cSmLoasnBB2sZDyhtuWcheeSrCfeN82QWasHHcbTOoAd3PntjvGAAzJeYUCogsF8
rVqfeAP7LAYUdGgqLW9X9pZyUTD4GQarpYIVaklSMaHYzhedx2yCtodFGVwBCJDp
ygdOg9z9S1C5k/jjVcaCMT+xowg5C3eLu3j/FhNahRVUropcSvh9dC7KQwa2f1k2
ykcDUxNa1hmpB3wnWs6+iZIpEBMznktY90gmmK1pWHx4J38Tq5idO0JV6Xe4QQKv
IIb5gC+J3UMiF8Te8Gluc+3oXc3v+OH1k76Q/jCP9d42VhWg4JrtJrnfkDSz1++E
eRwS4UfdSZayY8pVQqNkMwpia3Yjbwlywj+TuXCa5qB/n1dmUDQwO0aEE4SUm42z
k67XAlO+f4KqDZ0mhMmFugdFdosB9/6wZrz78OQagOoLddmVKOjw+qFf3VHDW391
921jjveSRN9QoGVOtHmldTG7yXT71q2n3DyomIWo1QGReQgiMHA6SET5jQltEg5b
Vv2Uwl331Y68kuALHRcj8CuxYyVzTuLriFgZEq8NirbbdY752kvgs20Mw0wdwYbd
7jLmmts+kqjDj6PTebVVEVyRkt+YHsod11uTF0WskSHzufR8wK8eY7curv0Eeysg
IPttT3L96jtuo7lRLYbZZ1u58sXhchPaYl+REV8hqQCDsO7r8Xg/7+yLfYxen3ti
oGQ6YQO5IMc9PQiW6i9+QnisVF4veyc7jSAu81FSJ0CGqO2Ln2h9KGIZBBTGy0KC
HEw0h9Y4EJhQMsxCmYpz1aSbRGMeYjw3h+epABEHk+t3MdxtA8tElpgrsBDCY9L0
WcgQOQGDQlXmssluTP3yaOsXkn/njYxOuemvgIHvYgEHpA8zOtfpDoKzjRGagzrw
PDr9kBEFyrSpEQWUXLfditYtOHejtpPD/f8xvWozrajjUDduRYvKxCR9WgRLxp1p
V9CHzBI23zOrKuCaeMBb9qOAUHAvBqbiR+YAbSCJZQZAMlh0fqmMbiQceQi7YtPB
hS0oZiWr+qJN6IpsMg9DTrVah1s+1RDQsdkPQRReIKuFTzkHXKnMhTE0FMLbxsIB
Lx31Gy0cl9C+PeVJZZbMmGiP0bzo2KbIJZqkdia2dSNNgPpPsqvB1SG51pP5hfvu
N0Ekb1WR9+icU+ysqTA/MfADbBb6INaELtu8PjOVVaVyjXfLrEraq8Wk22dzHXRc
tPk5O9dDZ18L/0YRnxDIu+AebPOKmE3IR3KdbHwHkdJpUOGjaSXcAEqjjtgWA+Bk
fQgo0w3gGjBta7FHNTgGd9vxb/Ai7mP+ry7xXX0xZ4Udi8nhJ/cWsYoQZ2bW2KM+
mczpj9sTV2GJX6i8chmkzTtFPxBW9yLK0OsRfPIlUvAIglp7ZYN5qMsi5Js04ywj
I3TxEwxv3Z5XYEG4Yqb3IGtvQH0jICLOG5APu+lox783Gt9kTLTW5xB7AXW6Q8po
UEbZVI6mytZ33CvqZOyTuagL8duyEp+A/xuvReTOJL7TeOw/3ITP1mZ8gOxjxMt9
d9BsTa+fhtOwQcqcX+jAh9E8C0DSVdJWpwjUK7VowBdlgIuZSvv7pkkg3HxbHzXa
3oJezFCpUGrXsJpdD4ubTneT7axz+BdbxANVd0dbHKESpsaqpi80hhf4kyeNHEN3
dPB1jJP9wEyHf3DCCmVdBZPG9ShjXEX4aC4oD+4WBtCyJ8XXclKPaUvQ3uROxKqB
VGfOETk5mEB+ocoUGO62eUNvpptnHdK0RZNAmche0ie4IDkgomq/1QtgUrJ0MEbV
baVtU/sbf25O/k5bYbfGmC0ZU0xiZJW0W20JAJVKBjImaBrCkmxbm4kjGLLrjnGW
yxgb8gDpJaslLSqSnmCHRJpMAQmJNZGQhQ2DJyijwzj9sw8nVSzlifM10Fri/rRm
XFhIvmzGaEvX8qSGgU6X1sVd5lw4dTsiN+8FWC4WRtdefHKXrhGi9PRfN6ZygRtk
j/p3Y/qOEofkbc9ndoU8AWE1e6M1zT7Z6QcE6nhDilU8rnEYj/GwDOVfZ1woU+tA
MUoarYoMHqfjIzKAxndMI+hBftxjZDiOVnj2hIJtWtNf/DoLgSQFxwtXqzHgs1eh
Qp8DY25JFmeL0chHcObxSAfuzOxH/nNC0WPo4y5OodK4fRMNlwncG6PQvixPIWvv
wv37ygcxzQ5890KEPEfN7w7EFp2TaRvO1VJBJNV5pw67Ph6jMDwC3FPyla/oxVZf
0wVT1GZGUBEQfVufpf87nMtWwyVj5I5FtIfo0ggZY1juFb18Ynwt+txvx0K5ws2k
UERH8uznBYdF+SNzptOqpjSFIj9IGjpzc+H5+ibk0Re030cBI5QO0jnJNSo44DzO
LIAQjzIhtCs96kCsVDdnCxULemaNannkcFhHemlfbv4ScXIcihJbHiaSZTFI5TGU
zswogWDZ8mwqRbcOG23SefJM3lfUsJvpwKvFEwbws+9WmwjqldyePhD9LhPD9W4J
FP2v+053VNAPYmSC01oIFcjWDe8sW8TNQarhrOSwSk8wRcxje+M2vObiv01NaG2+
YZI7VpCSB/QI1LhI/mzofkVSYZb9uIhuCTsbKMO11YVXt1FnhOJcebx3PFfVw/TQ
WcfbJ7C5hI1ERmwrFnkvlREzDebDxPGi6M7wJzd2W1uG9Jqlk0bg4RVp5xisIIZ3
72V8nZuJuvL/3iWmCeH7nudfN4y2Wd2OZ2bK4TbR1a65c4jqPXsYSU3kdaQUQ3Zz
FNJ4g28+N9uJwFM8WOkAjMDZ5KFAbj6gPW6jR2gH759X4AxTmUCvDE+ZdPCmG4MU
MtaRDYvThTA/grenUQTV+EGQJpB6MhyX2Y9Sfr+xe1mkG39quI812Wv9B1Dy1Q2w
PZnPzXXbnhhAOBTr7tXIlaz5P6YTlRpGkpVGKjfxVYOq3VUMnWNn7AcicCqfvv0x
mFtOmH/2Hi+0DY4GDBbH+RNn1nM06QbjJjo9mlZIEw8tMucOmAsILkt2MAG+ZnH3
4q2ZQTgFs/3nfivS4pWMf8XJrpwAI8bmnvNpbYU6aJedXbNOcaUAxE83tVF3wXPB
REstfysNOXoJ2t1SvDtazg0zsepXhyyt+HLZ2Vo4O6gkfxhPIRV+jao6qK5Q+d86
eZe1yPyTn8fa3qPJqmmBFnw6dhJhZqME5qSvZicSlspNKFQnyonfqB2T8zM/jGX8
WSaX/HDMhsfoYIh7+6s6sddvqnZtU3LBfVu+54n60wMAnQpYBPQwog5nctnG215P
lBy9p/UMet7LIq7LV2ZIuKNUR9JLPFjhiO2BBL5R0atRa0o6cG5ZPSqqlRZsp22a
q7mTI4mRijpzCEbZpmlUl6QD52PnwmmPHvwHOGuCRmL0cOjnisLeMd64lRwPK6iR
DXK6Byvv1TcHSRqTSZ2ZVGgXW155SE/G6tjHhPke9k0Uf6Or3EP2vr0bnv1sVeiO
Nrp/+frB9XdzIXayrWr9chn5xyXJX3eJH5aRk1ZaOUvRE9OD3m1ymp2xYuuEY7ng
pQ4v6d3dQgrzIi1EJky1Jm/S3jqpMw80hd7Q5/vxTAwvFrJLzpfvXGK5kpGLAvY9
IImIOgnm6+3Yo/Vfm3cPqbjtCzts+Rxcz+Gl/w6Hde1RJgGSc4srabEVXi3ZUvYP
OfXGSAhVfhUlmcumlNOeVAahKNjIoPy+ZkNNL4dVi3M7lIkj/Yjn/H67z4n1OdKh
Xen1Yakvx0gF7j0c+QltfI1/r1USj5+F0MDJCFY5qSt22o0/q6pIy63q+gcBZ7Kt
C4SWYYYwENhUGFZjWrZsF3TOVVrNzRv7YctFkLF6Q2J9aAwyIkkX6KcmPXcQ1LHo
1zSW5bQJ1568jj5qUl0MD+a1y7f9lSd0EM+31UVaKy6XwTSbA563nCHGm6wCGwBq
KSELMfHWvaifyYeLOJpaCSjuk2PWQw5sGTJMW4+XWGYrH+0OAlQFXzZgZSRm0w0c
azYDEqWD5UynU+5xapDvTfvg4UbS2JQqpOANuQY14bjz8aFzM/uRJSPQTfZ3vJxg
Ja/OwyJfER20GMbIFi0In5ilvnq3i1qmpj7t/0daWaXcOf2lheu+NXRpj3T3lg8e
9Mhs0qtyFN1z2WaRInTrpLvl+LDF47npB2+BwnuvLovFB3+QiIkGU5sbuPl+/4G4
3NP2ZzQUJFn7P37CBqyX6JvX9sN34IlXbFybt594p9Ysr3NwWRwjVspykKFliHEx
BZ0cVnHnLANKSjzhReGG0s9SgEUq8q2ukFHUNMregEsMyVogxQjl8q/eT31s4lAD
28/5v/abzFZUF6U8J+obwFGuuT/nBRY54wSZVJCyBVgGw8SHGaombu0ogH3nZAV0
6j4PjV60tQthMAa7jH55Wkdc81WumNBJdXj7XuO6kT4Pv79lCcpVoViGv5+YhGa3
R//R6vAe2kOhgcY/1nHdyALlN97P4oqLzzZ7ZB3qD4pP375tVRepXSkzje0C3r0/
nv894yhGVuDtcy1dWZqEB0BACvxqXYRU8n+qkjXijphHmczM8u0pt2xw/sU+ACxo
IYaHkM5VSoubrXhwRh33pMhAB3oUGNpx1RhBiBSTnqvOAvGu0qP283lRHGMuGN48
BH6a+JLkiU3hAkXtSUcITFiCyenHAcSH6nfI7hFfnFKjvLXZ5cMQjDkGYfXNvOuP
1AXmRdyQ/NAsAUr9pwfMeOySeDk+hT3S6xXkwMLPfvbZKpiHbv3B1IYkYx840hbg
Mkw0LMamiIBOHi50yEZ8zrteHZRwncRPNLUOaRJIBCn16NXHcKte6Dg70XE8Il0l
6tmvUjvAIPybN5fXI7zUIegMKS5lPHyd6DzdB6twMfOuEFH20GqLKY7AapyC0RNT
Ih4wa5onFEPqeDDLp20QLichhgOSR/0rtuk2k8iqBAcK7m3sFCRiIQWR20TPzABk
aWskOeMkY0ao1v+zvNY+leXDI4SfJZejfabFb3ntCphy2AnvxXoYG/PR07kcqcLN
41zCumsF/7IyQ11J5yi6ABF85bB+ZcNk1MzXEIs4wKIRfCXaYRC5081HX1QCWM/x
MKT4IEsBHzivTqVfrgZMES1kiIEjbX+7Es82qGkPo06UJOQoYH5Le7/YGY37S37H
nqF/587y+qNAKbaJZ/f8DLU3QFjzwisgo75coQUbR4NRS6XeaDgOD7LsdlIrRRog
ghK18IapehcjX7uvBWop5dgr1fchhavNMXd739Eo7lYAQIkvZJkAvajnxYwWHZhg
rfBKK7jfZIEji8j/LPH5Tqz880TC8AwC25XfTx7rKx6pwwT+2RzllcD2/LrALnUu
fedtiOHNoVd2jAEUHTsT3ptSuV5iS/rV7Y8ROFrOIsZrTF1stbHQ2HWQa9Rj3JWc
l4HWNhMGLFf+erORpdlGlj5dQDH3ti7veNgU+TI/BkGPwUL0Mf5zvY1YTSslt9b8
WLvXeLco94sWCq/rZ+nwhETVYT3K6vHe/vFO6xOD1bfyUlRWResttEvZYR4d6T1A
47yVzP9s4lkviaoR0XH2WozAOUJAcJlMyoRxswndo1CtYhwntAPKEOYoWUTmqXnP
iyoIqH9qQ/b5Sz0FBV4BftoWZ8KjGgiJfYJZuvgNAIqGdQ1rsMCTfps/+qc//+XY
oqE95MeBHM8BlyktzuYwaBtNhp4oVYkJGsCkXloScEU3yQzXFOBJdaehEMz0w1gc
hYUY2bIssBt/thl41Lbmn8z6JLQD+bL5aO8MVw3SJXEB5AETIFeT5zBUvP2aaNu1
5vPH81m0D7AGBnu+i8RbtYkAC5CNgZ4INtQUDquz0aGEwHpI2sTb8qXS+/VGIH5w
kwcq04kXKL2O4aSAVmPjgoTsezIahMSp+Rgpiuo1o8RfvNWLx/HJg0nxHfo2whOf
7fJgcctLdDzJSnzGSD8hDZEQ9P/HYKRJoZ+Ac4633/dUbcweJIzvJoHYbOVBO3B/
r70Eu6GWiGhVhk7AyBoa3Xagd9jw6QAKzgZPZMtmbsKYrxNXpvfj4ZhullCA4nTd
0RovkKCTE+EwcwpFpmlCt9s7QNmTwGwgGhdlsMWebCST2WwXm2DHHhTTh+h5GesB
X1PoYjtoilCOv1zBRArLMWSTtis2ysspA1lAO1ON5Y/DiZnPN4Xr6zw6CmXg5Pe3
FfzKYDUmSLpHZVEQFVCZPpvC0YAEAbEYvYlsLDiRIGK0l9I99GCQarXCvDUSCiJw
ET9MRb2ZXM/P8xJxfuSg+UjE4nue+okEWC4/BW/32KVFldTOfIkQJug+os2NrPfF
bpQOz6ajCuHbSXDWzJ812UVEd7i/o1C4gHzAQyFnPqhg4vPfDHpIFyHNDiD7i18M
YHlGWa5xcKykx5kqypvA6jIrsxp2B4vQtt+hEa1u0V+FzzsEwKFLhtKzHRES5GaF
pO9gm5GCSVATfo9SAqvN5PJnSye9k6rCLazuGWF7BNuliRMVncIsUiJwN+rELez5
WjRvu/URKhsk8pvOWfzZqx5V393Q++ipNT1mwKvNrO2bGLOr9whv7cDVwWXAxQKh
UdAui05nZSQL6a0byQy4FIsChrceO41FgLx5e5t8Pfv5J58tZ9sN4fJjYFwzn952
kgnD88eJQla8YQP1vVMEptg8Z4BgB7U7hMlUCoo68eiOoLcce5Y+LS+ZZy52d4OI
RKHnTOtGH1mP1aNagisLnlzCMaD7XEM6BYSLVg0YZMZWYyAuzO5Ms1/Nw2B11ELL
vVWSaSTrtjC/0/fC/b+UfdLaXW0p8Qr/EHw1E3E3vah1f1YkSmDQSfmb8zVHVCca
7MyE2y7AFPdLpu2Fh3ayN562iHrBxyWrirBxNuQ0ss9xnZXVbqFbMckNjBm9Xh5k
/MLRDqkVvfbfSpIn/0vHBFQBkunAuNTHxhRkAwpIjNnN69O/2Oy+nu1sGmvMgWFL
7296LvY+5tpSfTGD1vQw+Z3Dk0ipZABax3lFzWHshmpECIizcUiblIIk4LXiXmsU
YqVqtiG/DBFm4kuT7RSbLn+x6JGxqV7a7YshI+btdm5aMcJ79wzqS2CBSkdaLHcV
RrAwwFNAB7alPiUtnZDbZPS45OIcSW6LOa8u8scybwsR+d/Mo8TaWvh5BVf/DMTe
c49anYdikc/Iq2a4WW5fQE4JQ5YtBLrQAZpS/QZOzlAE7bfT0TDeJDhRGiRyopdG
Xae4N6hylyJlApbAVbCc5sC3Vsaa9Mm3f9tAFIZoroLQ0jnlgUvmUHcWz6hhyM/X
InxpnXLCDrhXPg9o3r5SxHzVMPdIRQc+fFljS4iJ1WK4LaiaP7VZukYIVspSS6wN
SdfidMnGkcXpAFUJmU5jdZ60FOQrg/oAOS1tp0+vJDmv36RoMRg3PkMIyXjCZIoT
bQvWwWcyjjht2RCOpS6BJdSDEa0cytYNhoST5ftnKK2eJxpLw2NEBAi4ySG0merh
hV99TtAnL5Gzdy/2tiTIEc7z5HbtZC8q90NNXkL1SuoIGV/a3Vwu+tckoR9vWvEU
Yc6ZrhVt2BGB3UxsLfjDBzq6zR4J5DcMd1X/myVWPRZubf9Sfz+I3rl4mAgn+gtW
rqQDhfwWJOh9uWwDTfvdTgKYwis42ErLRhV5kJXUu6IDNDscuOqJ2lDvYJ4Akymd
BuxAhvRmZhl9oU8/gIFECACsL1SXrVNQoowXdMxx8mvjYoco+cRberFmQ4t0+bgy
JdZi+a7hSNeAyXUJLvq7mLJDR7a9vzuo0iVwfrv7Uw/SBxRMWQtUYUGQSaUWryym
HMhgQ3rBvkCzu+JgoKOgLqqoZd5pjaT6T+BPTRj8fkm8BYuXmPUh2e3TdvoDXuFs
lu8xmjhSdObXWPh/Jziaks85ohk9jtdWe0UkNqeIH++ro13OXyKd8hoSdKsjzOEg
F+Ezf9IchhCAH3IKIMuj/jnapZXtz6DAaBCBtJFBgLH0BWYAQjwlfIrSivqd5Cpz
AbqK0NiOn1fOuuxMXuVs2t3fdZX2m5SP+eheoBXucNGw3hps22zOwnp+3Uz3DDH9
xG3XfXnpT3hWY0WLDrgtVfrwRn0uuuWonUrAjoE+Nn4qr1J8/5iDR1+PJQc6ZqOu
smvDrKovTOzKFFGyt1WP8Z1ENHbpv9PTncgYGCCb7vcWhWeMnVSVoVm7QTPOXZDM
hENhQT5Ttt3WX/8pfh1ebOHWwAjqJVARR/MHUaQsZbaB8rAtHoOnf4AKVHNohkL/
Ed2/Ge9PEIxOIY5rkS2idhwAwfkjLX1STVb40+Z+fgRMCMGP3nLrwAiuHC8Wooj5
WD5wzDzVz31Yjx+3aze4i0BbfYfvh+EXyfQnRrZk+m1RP1pmVWrbKvRUJTQooQDV
YPhlS+hQpCu8iY8yrlUlv9rf84vT9/EIszflrnOFpj2GEugkWGC8b1WiyCPUqcNs
faGBnksKCnnLjMhR1worOmVeOWOlSiMBB7YFv2D9PTgq52d6Av0EErFUJYD+aiyX
V4uXEiZ+9Jr1FqmP0TLVQAiyb1Fr68dnfymwTVV0SEfNtY96jD4f1yKLK0Nz3dnb
Tya69vdPEhgXoyqBwn1Gfmqa5K/xhPaPGspjNpzerj2bVgCbNQhtCeXj4p+X13eF
ZnKU5q8ponTUaQqkTlxU/YDi0/u6a5c4Lw/IvN9tjJFaro0k8dmpsUXVw5tjvkJP
bXtGNoF5vYpYeljRx+QWo7UnU21uxGJgB9sVWYDitiKiKTcvaW+SSh8piqzeoStH
N989Wy3jFbH0Qy7pl5Ifd3zYc/tC92TkwgDyuKv7zU1eXFbJWTOw1BaBBjBk/xkh
4S84XECauuBTTFBEbexDPZb3Du6SVhqfo7kuZomcn0nJ/6cQ+WyNjMyHu3p8WoI7
QsokpWSxf7oO76AwRFF+59a+xLqn5a4SbGye9+gpoVdDJ1WMbDcIKNxT0+HtPteF
IsCkdOsFbZtK7ySI6CyiP5SiDA/2wmUo1q+bpIUCDXvjyCK4uStz7/cu27ixKQdp
DtPDfjkIcHo2GyxH1s2GVA185zEdHISDmsksyv4Q0XcNwnu+jq16w9tAol7dJuSq
mNFiG8/qKFeAFUMIBLjMv62jDOGOQEdAdf0PWLfawI4RYBtfuDZukiC2OdG8Pka2
9xK9+PvcR+kKwJPVMgZI+3sV18Wi81d4OhiVTfnhhd9uzAWohH2XPxJXowpOMsmx
gKmzlySTm76fH3FCSz5IH4nLmpLAUUwNduIFHBb4XB6fcP8DNVSGSh/dfXRkpa8B
TDnqqFxy5YE9b4Ovcj27y+nPaGexXlGXGhdhkotVpkDpeU7A2duHO8I+NQYfEaXr
Vjr4uj6b4JOgJDLitM6NYKcG2pZ5cd/lM2ajRgOcclJevVY47oNwtnxUfUuXVUeF
8vJVe1rvxjJ+DwB1YOBW6DWMcIBD2YdnpoyQ5MvdpalR7evwJRRRgAhBVovq/6co
BkiLR0kWjgPjuy+hdqn5imHaGGr8IbShrlvAIj9dOVbC8t9+96DWN8oUzR4ftkMH
oQjtLBybTw95+/bDEs7Ovk9AZwQlQMf1L2gQ6+505hvaikc4zW77E3R1df4BKxXq
6pR+ZbeqQuO4msk8OQ3UYaD5mI9hKwRjWGei/iEq+R8YG+YGrX2x2+6fRRbarbMf
bpdWBV2a29AcPCRWpFSCyoHXGBnDdbdFIGUn4LDfYhDwV0eU8+HAh+tC6fKujCUH
53XN+CtiLzOFdzLpmoSwP6KdZll2L7ysL1CjYC8R6VtPyU5MW/jYW4w8vDvm1Mn8
0rMOWwl8kBMn4yuz6hOzLEoGfK2PTuTqK49bzX8CRoK0P/EO9pivFLeguGR0KLbt
O5wCQWfQ4+ukiqei2sb7bBRgYjuDWKIS5s0ppHC/ZHFZVGcnTxEdxNEccQGHtXQY
BGF3RekMPHSHGudk5T4mKFLkPz0nfgpswV2FGPD+mj9BKDKEoLXpkQvDpOA60hPI
3ftr4YW2GZ3gzVd/eJ8+r6Ka34uJjFX/X2OMBA2m2W2ZxiJWjQJjtszSSvQL54Or
kk85019N53LWMcF4EpW3WFBtLD2qs4sSCgGToYlQoOrVLiPXvw9baD9kC/G39fxS
eq4wvqhiMhA2rWnfPdE2X/Wo1V/cKLg/t7JWmQ4v2Iv7V7ubYmuauQelYP/E1kIs
/HNw4EAQlUYPdPntKG+W/S8g75YweeyS11erGNpL555Sr28qTgwpl2sXb9YOVpsb
QgJhmCZr/t5+JlKeYxJIBSAwVLUdDx0bL7vwUjQUE/a029T1JJvUAmYqCCPyOqzl
XkCjUi0r9wpS2nHF3+LxELy7hcg8s0dr+oh9IXxtnBkp73euszFEJ4h8Cq1sgGPF
aBmIyBGK/55J4Ku/XCSiqQ4bEHD6O3qLsnCJWzP8UHK09jpjTEF9/JrGhG84ymJd
qnaz4q88F7Tb7I0IKb2A2tztHIiN/WByvT9U35FTLfPIGEdt3tg6U6eTwS/kKTOd
IUuPS0rVvz1I6rPaZJysbP2Ryhf/u1hUJy+jBIFsugKpWL2vAhC7sm3Dk1kID+Zc
5wjPuh0PK7dcOnmIUtifVnXfOgU9Av7lSSW2KYbX2nvCdYcoiZXVaQd2oXBZ7PLu
aspUM2Ri9oiS8kDVaz8kkYa0Rtdokk7EWNyFYELWRZLNpa2RP/r5CZlvLBDWkyPL
TOdWrITqfEAjlbmlsV7dDeY3Tpdi8j+cUqg/zfY0sjHU2Qsqt95Y2SBWqbmIawK0
0PiN/vpSAcCRC6LuO2R8yZG1qc5uGAXBZbMKlx/O1o0IbuD6tyb+wBT3LUu9bJZf
wChmB9cyaOfGZRqhmRzzQ03rXDsGZ17/zpioRBrUYc6jIkKuW/DF/s0Otf/q4DzN
xBsRWOKnXUy7JohejPt2ljTqgzkipnCF3KLMLmXVE0jmfNAJyvspfPMX1KvveBuk
bZLv6WfJQnCGQXLgQ8MGqIqGIwC8VqBJi+u5KWR+q4MYdcoxAMesZumFS7TV/LVU
Ip3MFYmebdrv2A5RBnFkwnUBWCiy5uyC+VU4Yp2XMdaWjOEF3ZW8qeiNF/Oyd2UF
RSqfzLZIvmRYGb6F8z1DxAPnZw6fRIPOpFvUZNS7C4xzPe68al0tVYDrzlhID9Q2
uvTHKZ07MOLivEWN0cda641KFYWDURcftgQ0xYejsdGjgQNPHTzKAsNFweCjzRJL
GWe3edyayKAEHuciiLF8V2e+7sDWolVr3z8qzlHIyIaLXwXz6c+Y8vt1T76gRnQq
BQEKXgQA7hXQiGtf5e+GZufGW78xNeqbbXX8ftjOKHn5PuXEleHQaf7jZf5rLSgQ
PY+GhM3xOZIYMIOSFuOanXWWv5u+uU4qE467VkOTOiv71HlCqHQoN2hi/RfBAW3V
5+C3Me3t49BvruSimbhpGQIqerrtGt6VLd+sRQCsyTLSWhns4CntXLQrfekNAHfB
5l6+HP+FmOLNQoMWlo4RixRzBZfjAXdqyRODCjeXoHwOUWy5DftA9lz1xtJnQafF
ohhEMcua5UE7r62MwfgUFnxtVKYQPpu+tMbQ221MSWYtsDUBG3AekzCenMxuJXXO
39WLia+oVTPsg/EinXSzBoVmrTLnLUkm9gUPbAacsAB2FitdTZYxpRe70H2J8Nx7
8F0X2+tTIkztU3OAZZLXlks1TJdeKhrzcrrNigBFLPsVBc03/qNrXZjY2q1RAMDZ
7Gi6xDyHjV1gfhQ0AwJ7MQYaJdMuuSG53pGay64T1eIG/1FDU6Ahmg+OYwoLEtMo
qqcnFkXkx7tup2XUfNybYRI3PpBrlOdQ1/7fF5MKbK9LFMJts028lOc0l41amLpF
50Xdqp8eQyOeTTt2KhWX+mNs4CO9g8GkyvJBQBFKxtv4wH2LNBmsdnADiyhuRGqI
Etg5Ar3MdPIfqC57OuHhCqakJ+WyipOiK/wHQcj5tFqwpzglsB+o0rtuhFJgTk3f
qLxR2lcbsYJGNS29s5vWvlNUD0+b14t4I+VmHU0ETdFwuSlZibEPLP+k2YPAWaF7
Y4R6OU77CkpWgiqf2WfJI3QCL0yLuMWzsUXgkQh6FqMkYkUkxqzC96gZJOTZIy4p
nwj2qoS4SHzpt88qcthn2WhwBd5G1cVd4Yw8sAEN3Ua9NmLdjbo2gLXq9BNKQ1p6
4g6DlO+ETQS9CPKnPBfG/3sj5B4qSCeLXv2X+Fw3icD2eUl2X0MPM4tSLsUvrwC3
Xeep7HM4TO0Q7Ei2QKvXD/Q8Qj95lfVdM8uLI1IIgK8Ue7cC/A0ix39inuxyMXrx
LPt/aLmvLkZ32MHzz/cmAqarA5M/zjK9dlGZQj6FOmTsipzrmbmHwT4/lertKxss
aJMBOSzcIlo4QbZFjTZZzNfTI5FQeSNIGQspBnsx71FqA3QnQr41VEZdF/qgqld8
rQolo/e75oMV6B5w0M+Ivi7okSC84MsNZ9msyVPh65fE5fipaVRewBKcjJ/0Hkrh
3WgPH8ALEBzEVD3VoqRVE9Utd1wWSzCAuF2kVIeIk8konT/G1Pl1sUREPzVbixv/
uZszqPpdHJtMdT36lqQTU9+Vca8ujmD7dxhUkwQps+tc/1aeX3WlNZ1gQ/kr3DFa
i8FfMGzUPBFGJn/YUJ8jbXeXwfvrQJrelj2bGdW4yqi8bw+MbZumCgyuyx+eUDD6
dXK+crDnzQahHzuEWRyt2Rqcu+mWv8URYPvofY8elxiB7yhYppOLGujzTZCFNhJ9
rkmuOpXPdB5xweAcqESujMOOgDFG4a4SvE5y1oJ/Rs/jySaAcu29i1aqwh/OP/Ad
rDsYI6FOFzhOwWL+CrbcoZBxz+jonJiLABJMMAGkbfgVzmzjbdzmaW4/Tdz/LeNb
+R/3qak0VyEzedlj7VrYDhovNWTgYE66u8yf+MYIQlt+zXZauSeqAZnSrEfToJ2v
U15xzYZesJ9rLinIylGXwupnfGj8w++ve892L5pQdX/Cw+hYTCxprOlRlEYWSXGH
EAKK4KXm4MiyBHXp/FnzVybTAnWlq1Ysj4Nbus/8duv5FGve6TXR5WQE9bU2jUZQ
YHe6vDebenAwnNksvFAF/2ltzQFs3OCNGKJ/Bamjn8KwynXpiG0MwCqtbD/3VNhg
dzaHFrFvw/9hYKZJxzyVErvxP5arok5xBOOpfOU4Oj6ca0jCPjI+SH4KqSir3YXo
UmuS/ea8DUnOmfOTZm67ONXKkqvkwf7w6MfmT5s7nFa5FhEPyrTZc7wIN+VrRR8h
/Cz5SSgSxcNgESNUGB8pjtRoE+MoXMJ+dOgZnKikYyceD+RsylQMuVGkehxmO0cT
4vrAxqgfb3EsQhhbCJAMO76jyxlx4am24fkQWcmj9Xj3kGWiVxleu4+5fvjMhZHc
qwJL7qBQmY4spwsKk3SXIFJ1j9uLYzBm0V7Y4Bo/vaGphratUqPPQG1rIIptDMrs
KqIF+2h+8Y+An0zJv2SpIfeHTX3R0V1BrjMfnGrXPJckkQRMyd4UJJZ8X9dhKcit
Az1YylbXUVFutkm7wRfDqragGTF4moDQgd1qJMpu8AmkvkK7gyP1Btl8zm4J5UwE
Mx0MJFkwm3EasSsk5J1iC/NI8vwg+inEoY7iioAZupJEz45WLLJrjTYl68aZgBMv
MC4O1K/Il3EBXv+/q3wYQGUTUhUUyIfbi5INAzZAHwG193UEuzyU7hUHdfqLBdNg
CWzfhTzXLPf8myJU/USmeOaXGVAEil92PWGeDzuNwqfbAYGVpXQyLy+eTXMbfn1J
dZ028povkYYWULQwMeKtyEifLswxyegdnEZxKv0BJ9VOXujcjC50GKcAOjuykfjf
3i9zCU9yYNfvmH5tuDtQ6OCxBZ00r3R4k6Qp1aEEE3gtHClCIpOvtLOcxUQN9+yP
tIvEOcCgSMMEQoIrUNglQY2oUfGIO8Ev66894PHzDvSf2Y1y+pykHv+oW2cIXlBD
wemgWRnz+f24tDOUstjj7Q0kNraZQ1P+Z6wwoUP0mkXZahZ2KPHkXkKKlE/k8CoC
KrmLBzUzW8jHTiMw6UCr2RM/mGeSPC0Uj0diRNMjzLuW+2W9b1gUfnI/TtHAbNMf
p2vNdFtBbv9JQtXA53mt+TpgXT8M4yYwZ5Z+I+wKr23B2V0YR3Gjn7o8kmocX2sW
K5dCkI/Mp1Y380+cG69NS7ab4XdLoYoKjG1MFahbhhBcIYVvlOFp5DOWNB6bRdUm
Ze8pLjIObDWDqLTne/qaGWXABGtULGnccT4jv7EC0YLtuNwp+RvgzA5gDLpclrkC
m3mt7DtNukW4Ek4CEJPRr/1HPE2lmAmE0Q4SKIdzwQymxpVZkN/MpvvnUB95d/Sy
qgo/1cFNqqbQ2S4C0zF0FWPk3G+FGb9XxhX3X1FoK206cC5nY5O+Xe9I3inuVOvm
3J68EkpnQK1AEhYxiCTRr2uMIqrYDa/X6M9PGeisJgsxOFLrMlxIeldoylcfYT5q
Q9VdkBtlpZqaLHY/SE5GGyEm1Hoztt1bI+2ceygB9+mCQsWxpuNyt22fKe7dVLvD
DImenpMZW0scM/YrJGlzrbC5aGAK/3DRWr5zywQ84ogU9Ioy4FqjnSDO21BAGVKx
NJZ2A/qMEsescWR9opCUhiKm+SCXdZWHuGSZ8D9cdbbRqmm49qQEELFgjwGhmwRq
DU3AbO24x3JqvE6eP2tmaL8u2PPKeOpO1IDzkDHTfL5D6GH/6uHh3voE9ZWD/0s1
78GjJiMcrXARC+vINXxlZaJvlqWMxgDZg1JN5TeVv2X68SfQDiecxTNnlgpim5Oq
3aaJkNTod0PwpSn2QISPmU7og//45GeolhutNNOEXIk+iZZ+HZ6+xANIz3AB39KH
V4ToRehrxyfBbKmsbcs7GP8VF+yckgQN0dJMs/fxgGb9bwSQ3kh0e+BsNuU7kc/w
QE2Fe+c+AAy+jX9pzh+HBMq/qz43EmLIQyanbZ5NYNChR5SYtXA0w1B3TbzeIvNu
Ov0RyScC6vxKJgROtK9HqSD8PLXV6VdWfF3jGZNeVhxTeF7+wKbWDiYdz/pDT2gZ
uRL33paNcez1agLF1m5sUBystn5BhHA+8jI/Az3d9ustgx5O1a/WO+uZBbcuX7gY
OzNxE5vNO4JJAqoMcom5xghnSiCr/+cv+TwQxx1ugo+DkcQmWBtuWz/YL7yJjGVA
iCpTX+Zl5CaRWz/YUDD30ttTPwFuA4hQry4YJne7yYJmVJZ5d2W4v4/PCkhgyfpC
agcu6hTLrqV1RK+jp9v8L7g7TwxaiCWfVWowRnetGNCnJKzFXHr7EaYcJwHZ98Al
u9MeKgDAq7K1QvMjywF0cU9bt4EcTfnc9TDx8luaad87VXSo18NIBtyi7v6MWUJX
yiqbWUE8OETPxsaQHabIlLSkFR3Et97iLAVBJ7WkiyXRrVgZN0fVkUZWjK83dfEN
BohtPecTPgcMfcw5wOp3rtRK0Aw0J2zIqK09xGPSgeRwyLR5/bnFIokEZ1AOCgBo
iurK8j6bYeZ3nYcRr80uyjC6LhMIw70RIWNYNgnkPCgZ+8GqU7Mtuumy9BMhEpK3
Ceerg7tXDY/75uxFdDyZaaZfsiDVHxNHMmwRVXwIVmBHNZmPycH4EnR2MicYzXaD
qX6oa84tIZ0xQnAchbVOT8UCiQMdytyxtWgoaKFqzKrKId813ve4t8j42IU8Qadj
JKkJ4I0/a6Gb4n+MMwCR0QG1io1+DItksYcyp6ocKlDFU0/BZJPYtBBdCDlWYnxH
6OOKPjO7u02g1J126q0HClfwn/SgX5KPHgq2OMyHJvH1AopsyMfywNT98Hhr+Mi7
NIdb6zbPEKKJ00gmHQHcCvbyzYDRslrR/nmXbTPHGiJ+uUaDUhFgYkrd9MLJNRz/
Fq+uQoESuzCUFr3fERStnefZxodiFyXMuXFMgzvBO3sxIoiOgp29KRsimMlM+diV
yM3iQ63gCyA+chnD2EM7DYJvVVepwyz+IJKsGJbCIz5vYCtRrYXL6hnQnJk4Enmx
2wjpZ8024FTLx3lnodzvH76R8mAemEaOJXGF/iuWWToNaqNERoARy3DZuygZLF57
kx1+HQaG7p7x8GTi0T3OudyWxj+LcgnCrmQJV3Ldr9T79IMdArHRqg5bbSfQeXuU
oWIuTQmghc6dPGQhyF2K3wt0DpO7Q+z4gW7CSGXh6avwh+hjZnDNTFNKbhcUiTSD
+dLvY+6khSzwU2m96SV8Nr/sjq0H/+RkNoOthFpuXlJmTJYjbOQEKAtHm1pG+Kna
t1rvuoTp3xUrNj8ZNVinkCQEAyUtx9yczrAcM2jybaIeXBfin4SwcRMn2LSXfPlW
nlonc3EjrDKIxGu91giP0giX6GHXSMVxWwmycycmwFTJ7w51avOewkn0DOdmmQ4P
EDD1HzTPWWYAmep8qyPLyoVGYGICuwsdwUTmf4zXxKu7DzAhGhlKyEwMsa8+FeaF
TggBC6WALvPdzHIz4RuhMy5ChSCXbiVLJMGA+QXYV7u8GIxMfLIAovLHJ6vYiOvV
fuVpv/703EZbPQV0L+RNHsfw6+bqbbGq/Z7SgxYz58/NvHpznKJ8hr3tGNHU6nsn
jW+yVa4H42VWT6hWZANWJVFYINtVslW3EWV2hhWEPfb8+YN9JosBMxQDLTnJyf3Z
e+kex1KflxoNFb08rsicK0rCuUSGKtedD5II5g2T2sxLwTPLKrXqF0xZQ6N6cjyj
V+8ns5MHeXPi9WfWJ4Gw5YVvyF8clRKY9TFLegkVoWIaZ+F5xHgHvyjcKth4r9/z
4h9Fw1PziJdJi1LkMp2jNSWkOkpcEv3aKowVcdC3nf36K7/F2S+BhSLrMDr3XV/Y
tZxWfAZq62Oe8e7Bgzp1kJuY+N1ItJnrvuXc9yKfaTp24bI+I7if5HWi3nAQm/GR
chxBuCZ9MAJ21SFmW4GUf4dqm2PA26uiwrWZYKb4Xrf6SXUQEJHIisTCDM/FrBsj
tql6Kj0N+JL8WinA0+bmZMg02IP1by4PexOsgiy9mCPh6pADK4aE/iW4HCgera91
+D5KWktqIu8GMdADMuHzNuPO+3h9kqH/fq0uPkyJxR4FJr4ww2uSH1Yg2apfx9zm
4iCdgEWuOaFVJ/G+rwDUCkXD3wYjEyt5OKinZfOdwW6XWNPJXPcizKIrhtfkGhln
sdcdWq6btAM0utBmLGZVduCjoKdQ/YKV3OCJsZvK3Ta9/62gSveQGxVnIfLfF4F7
dF95gNHF3+EzA7glSoOKWEoALyFwnYtqs2xh3/KquGWwYj6E+x+wIunylmW8y4wT
hogxq7Hyj+fEPeCF/FMpVMk1FViyDLssC2NsEKW0M/tOmNf8uDFdLV/whQM4pW97
IJh07dQVT+vmnuePvfB2s6cnQzOdIfyPdeGtnzwCwWND11GdC3lFUaL0r3GJn7Zq
kB0uz7nttfoWKhw7R4l1O64CHf267EHvDycEmkWIjG+E7opqRQ1OqdW93QhlAwv4
tEdMRKZFL+gHTyEPU44wbmgMDF3CIBIZQXR4w5/vmT1L4Pey/Ru2zNNfU+ntnwg7
HHDRlVlVQpBqZqWCpxeYfTrt1OknzbHOP1JlldAookZiFxKj+reptEOS4vYX5Duo
9eCPVtTZFuCihTZUBDOcEWVVD4DRxqych9XmbXy3Ll0SUe66NrFgsLQ0QKz7HVtZ
uEkozcD/eHBELnBnQbnlu1/ebRkkbt7yJU2oVGH6Zbk9jC6s3LKLKGt0Pj5MIeqH
6vgdtMd6hBOIYnTMg+Db3NYHHZ2nsf65z+4SA5/edm/73lkr3FclG35OL09yb755
ev/cO7qGzhGVHLi6LcXhhbxywGn40gu3QzqG9Pd2yWjjvmMm67c/adq04h0nnK1c
FuW3mZJlYpyUDg9RJYu80zzpsVm92zsXi8YV1dQ1BQyU3Cqzel+xP/BS5RNaDwip
2Bn9yqApz9Zgj91UIqM8uAyr5k/7C/auyVKWXYCbgFjABHVQf91tm7CMdI+ki0hb
yURh980bBW2U6g1CE8/GLf8/d8M1Y4GrK5Es0VdLK5u9u+8vKuivibWYklYOzL2N
CAnt1lr1zimIzB4XVtyIIHZHFbonf0Pa4Vu+AD5dLHVrbBYmXndIl7BCPNnq4vej
kX6xECax1JUKOHy+Mh8rAE8jt4iwMX/WbidiVP3002c0ik1lCt2NEOQRPjcjgB8V
R8/2M5ItTv+CDEVU9y42v92/OIYnrEuOIQNxu0OgTeeugx2zXKEVaj3Ig5UcPaqX
lFtU/7ZapZ7V49U3mo+WAvaYXOxsQiNdf0HM9AQM9/aiQ5+N/mBD6PD63fzOFqbq
uzHBUPIakAQfPbYT7pPnSfpY3oN5MOi7q/T5cbb7XqFZSB+oWyO/I3ziXm5/msl1
OrlTyRpD3TwZuPUq28ymXGLP0kOSVYas9dxWt8ZKqKePTEjRSvjSeSvoheRycaLZ
jw1dh7yWwC5Q+FUuzVOfJONk8E70ScXy5qlovLC8UvlY+GyMpSMqJRT3FF6Ew4dZ
03tsxd8kCrogj4U0wAVqi4YqN1s220xztIyKVCZuhh6qbi+cpRALcTbzs0ZZluEi
k2LrRDC1XPmE7MOazrlIhDYHgOEFzfnchptan0aFOyRUTEqC+0SFYAT1JDHmJ7jo
YgQb4HK/oAb5m0mhe0iOZCRE2Qq3MBkgGrGlrClygaIX20Xwr2TYrz/Qn7BRH2QR
tM9BNX+/8pYLLmGbVDw86nU0HNGIzqdqvshxuZurbXAVUptp47h0KXOuzQkSGM1w
AvWdDgMvgjTndC+TA6oXXhewCpAblhPRQ3u6XakEZdMnORmSWA3LOnK/xjTZF3Dt
GhyN80bX+h6GwZEP8cvlmPVKrXAXZ2YtyTgrw8YbgCf4IRMB31TTEu5yj//D1X8/
ICPrtsdXd5ynSSxR56DL75N5HI8Barc9ynQ6GS0weg8mX99k02h2w1yEM5dIY33j
1ripU30K1DBhXYYWyJYE+0pB2cueoZVEBvl+sxuos1nBFLQiMCCERHGb0RFXe/+4
QbObF2B690QrBVdzfDD/CphQCtjqLC4/gkUhQNrRHcy8PwUHYLUwFbEuPEvljX8x
kRLpEyryX6fgnnv9cM1AOGk5fF0ObV9DSjCwQPRRoSg+w9VyEoJgyFWDlDFgwvlB
M1mqC4zACgPrfgB1VUYP+TYmS61hK5QjaAJlF0TLTnHagIVHq2iglU9eebj+vLP8
AY74aYxO8XuQJ6xgUh4jVQvk8qW1pCWCwdcc5dFr3dOFBSwUZuOO4UMhO6xZ/OPB
Ec9RbPdbEbZYncNRrvU8TIi4Ws3IsdVomaPd/zCQI04RSWtGE/+biHxlsLLAnl12
/4+ma2z2FhcLGPGJrlL0B0/KKdBfTeHCYPPpfh6ByENHp3PPOhaBIfuxHoC6Q5YP
18wiAP4/SiiiFQAiQ8+e9zupcM3egkxaqfHDu50N7iEYLPJ0sAIabzkgMvEl0I8l
oSHiv4q87o4ZFLFg/LQWFHiZ8xGuvcmcZsM+MMYhglUr2TRULcLQzyjTXO8mTbfU
Q0ZuDyGk+w/1t0symvM3wTrx1fuiVhWfSgU7IkAGEZkuiCp3MRsUSSi8sq9aissF
Jqa4i87D7bsbPQ6pUz0uyes7nFEJ/ralXVdRydEvc94VEXyixXyepWdaWnhoKnjd
sCovWqgKq30He3ZkvOR8bNDMn51YufDcnvhRngAbMLPv6ATDBLcdCFN7ujMlx0ls
vNivZD8zSAroUKewprD310hYOXMkOuqMcL6GgD18iQs6HVro99tVkmfqNDDUwERS
sjGzgR994v/VxhfwxC4N3nzxMiS0+vEAHAhBiUjyPSUZuZ/SD+HsUytpqtZOt6fQ
2JWqlNpw7ONQFqDBvQ0KZIIy7OcJmyDo65/C1oeN7SL8m0+gFeX6FEhoh48DUwCg
SKWVqnQuF8Pv+DmProLVDvH8SgEGvCfnQ7KO56oPm9JJmmMJqPGYGJT/e4S5gDie
VyoZ6Jvo96qsouxyUh+I6zD2efcC6hIsowYDkHfCwfFCnKchEScFVckG592Istxv
vZbbP3D4aUSNOMFDvSofBtVymcAQSz3Mebmzr3oIRl0MRFJgJyxQffS2cpOZ0XSr
I8Ty8rUsCZbFlZUMT/RANzuqve7434GAG7DTzYUxHCvH8XGCvAodcvdWFdXoKN6O
5cibTWxbYY++GISCBoI/SqDxCJ8H2ujS4kKICLYpf3gzMGQsoFdhNgpGGnRGNcIf
Dyzw8L/sKAQKoFauW7apFusKs2GfMxqfXyN51XHOs/jYibmZr1C0Kn7NPzIseDjn
Uxml2pq2+a5/0+E548Pg5tQALAgU4DfMeiVwey+vPu8xuTPv89C+j+0Rd50oSBJB
QKr/nkl5yBHgGWoesCWEyhH3wF+Wbz8BYPk+X23Ah1oOhrhXgmRA7FdH4hoFOxVb
bTGUXgFXxLnBRb/f8Y5kRZmt+ag7oazJGnM72QMeEGWM8t/F3AjEEGARNSEo2aDI
BAPZB8I6MnfM3Cb51y2lgdGR/iUqSntZgYFPVoYnqeAf7A+LZIahqrUextet4C2t
Wxjgs1+GA9n+rJQ6tQqduU/mJ1D91aqJcNTN2ql8bqFHZtUwBfclJhTXUxIKlAt+
NfPCE49VGljjycaVGjU9rKDSFe225qUmCEvHmQV58BsR96Y28yM8n/XQwxRDA2A7
4XKZuYAXWMoz7VHejozOTwYFKR2GXmX/M1zyjQRcEaLuDvznrEPJshUadihhYoBz
xga9E0HkNp5GYpj7W/v7Urh01t8IhI5sf5CNIeIv59NFoekKNFUedg63/Bor6ATv
4tJax3mVWP+NBpnnjuJZwfOnL6Jtl2ts9VPvAvxxffzg8MIJcNhsfHAyMMG/6ELk
TPb6kjJ20zoB6Q0Qlb5eVdExTixZhMl5WXlGmQ7DVH5TMI+qnbzCNC8pahRjZ508
91vK+hrd7KRxL1u6v+TXQkRx4x32E0bghKPwu2dmo5L+Iwi2NWl6etBUCnSM9kCY
jEdn60dTCzDzLh8zuFlQ/wVa6EShzVkL0X8i2+c3KKeWgmDq4GQEQ7EfHExkUwpR
empcm9A2hGgsYqjeeMDmtLCzHKSGmWfZ8qvcwvHpSznadNgCbDPv9id4APK/aClF
/61WlcZRYwQU7krMaS4nuZgvauMbqz9UD5Fa3Qa7wQzP9JCqx140Jz/JRxAjVSwW
TGcQiIyI8wN+GAG2J0C7bLXbzLJEo6nVd4UiUv5Gv29+wegBfRMhvCPzVhu3J6Aj
JywY66baTklTGZ0xNFQIfxfE3BStd9xvJlv4fTVrzhAOMb/Obcww73VfvkIA8UwQ
7hp02O9yzWlXs6M3br0sFsDmlNBvq+yCFmToIBqDLOdG+FKQg6Wz0pXBq+e5+5Y6
fEX61bf/CM+h3GgntUVpjdAdpsT9xOmuY0mqAPpHUHh4rWMYedS6Et5Z1xDwaG7I
YJaPqsio6uuBsH6PeuxI/qNqhwtkh3h8IufX0/7Qa/SFXKtoPbTtfnR+FK4KOD7Z
WrkoM3zIOpl0anJQ+107thtwTPbx79ig7BoHAzcnCS9vtXyPh7j9UiTiTMR+jiUh
mlLrnVj0tg+5tgSNZSGhfQvSx2vza3TpLrwjkmKVOpDlObXRk//hhoCgz1VzcQHn
v21XoKwbBEC3ZmmVw9WnGz1PAi2rrvL55TDbIGwMSUenRqOYQn2HwQ+eYT1g6MKL
Dw1sYlPbnDWrWR13Qjk2BE4332RBpiSxEq3JAgXn9fH2mbtaDrjzo8fWaYc2PfzB
auI15DhmTHelbQ3mB1oXHU6xVNkY9yoDnN2DGM6XHGQctQPNLhryujF2nkOhVx9c
T7uAbC6wEUeSonyzBJlXelmMRFiV9+s9SV+s9+0FuJaAAsTZmtYrMdVxdgohddBC
qiodeXdZ2zhevVKlhgHYokGccQLz6ocRyvsEY4DKUFUQNkwzb46OpEN+OBLdnn/d
Q0vtw8Ur0zOU93KEOOW9HvvAKvo1hX4jl58ha/gcVH5jrm1nolp/NuG9VsXF+n0h
Nzg/1elCV7e983nR6SWu7hgGwXINvI2LMWTUqqoca//iJTaVpnYy4TphKIQNhcnR
cElrrr45V6TlGwRzaDm2nBxEyK2m7W4BITFprVJjLyaqL0pm+oMEX7ebNPGkShqL
Y+TIW3eiJrxZ6xyVos5Waer4YLHGS/FYRqMQ+HVQstZTntcy/RWPbDodCKKQ/zS1
t+I7kbYV8Ejw3UNxURW55ohaIehztL3DG5J+AwpsLGIdV9MLiNgdpGVa0yyr47ns
oQJufiYr5XV8+rtLziKhJ9gbwhbg8J9GL+HbBmhCZwzb70M0tiNops3t5ZPkGKe5
Y77Go2gCvIhVxGx/77aghWY3PCnWEsJm3wcCnV4J34weaxGBhyDU9cIJayxxs/J4
hVlUPGHhiTbr2YGJkYoT/n7EUIgP+UPgH6loJ9r/aiuC+RmeH+e7S7xuV0HViotO
NxCemy2gAFjIUn+LYpPHc1hdIwgeWXcA3RMMH/BJo4au3k/POiS/cPHvSPzaN3h9
jumKrp2OKe1FzbpS/l1H+umfOrRwR8SQYgChhr44jxbrFPdkI46UcziKsZuRwlbH
A4+/D7yWipFBWyk4nXDBmAMFHyV3jIIhAOeOZ/HGbC3Duh8UZh2audMXMz1bTzG2
houFIecklB9r4NBzmqa4NMTrrjjyjluH4s2wSy4nWBncLLimN0K+7C7DOB7PdGiv
K/v/z1SVvweRxSmda+3Bz5NbBfFthG3ogDyqo2oqiR0OrYuGZqfYW1M4nv911iSM
bzveGBxiCZyGg1vE/1tOiDtTzSbOArguL6ijZHIdwleQk+jpw041bJvvsCaHBjqe
t2qIT45i5N4lD0foFi8AAfS2w7jb7OC/LoN29eK0MBFwcKSnUhWjKMaqPAwS6fqF
Q0tSBYWS5zfeQ7m6atFBNRWJhpmjUObtTvkvOgiAtIZWbF0bWRsehHsYhwHEfN4l
OARvo7XPYUoIdlLQvXkVU0M0unbQQ/u1GBSOaJKBU3dPNC1nsWRSuuDjwKoGOTsm
llJxWejjup2/NlUsnpKm6etRdsVQLBPuhg4UcvWQs5c21LUU/pIcwUtbtVzNLEjs
gvAxOkVu0K35v4PAHV1IivJ6CfkIPn1mpY371ucvxu1GZjUMva3C1+SuSjczf7rQ
jX3I9859taR0pzKrDsOsGBaaUBXk3kp0Fw3u3iaVck5HLA6dc+1VTEsgEveK3t8+
wWBvf84s+kv83wpDU9/RoxFLcQCxXKyAh3uagOlUGX1yTLiqJEXo6YR4C5I2ky8X
mGDj+GmdCFfO0+snpT6YnBHCfGkBSee/2YEv1FWNtczhIA0p6IIKha9OUvt+VqhE
x+Wse3Uvy4D/3Aeeh6fBxUH8PfMRzTx3XMzsZG4xj+/Ia4gYdcIi8MXNraN0rQvF
BinyCeTF0MwnE1s2R8pz0NgyL0RlIancEQkWilI8KgycWlFNx2roOsjrtTjgNL8A
TE2PC4zMp9mIha5DSRsAyCmy9L01fTZpkMsZsrLZ7IN/8Saf+LHMOyo69YAJ9N6Q
8YR0IHN+hCIniK+03M7eNFXjktWtoUGb0esbENg16yw4EixjKcLygZ5x2iFlUOpp
yznlTbN+lvVMNDOd+7KSuABE2folBGpAFUNmYLLQrQEAcQ+E8pQ7/LrdPkXQtkrF
6gEvtlmSRJrWAsPhLLI/CdDaVDupsRCrr6Bi2F4Q7kvIFXY1doQPckmQG51Gi8Ng
Vj1D8Z0y1/alsLeu3A9k+HoYzbbFuFfE8MVwXQPH5RUfRPxA98O1fB9SNwYhdKvk
fo7TRtJayXSwIJjJNC2i0B4XO2lPB/yOIpKXjWzPYxf/ALwpRKxya4SnlGmzIwrj
rKXfHUo7S/ZktZdsdfZV91E19KReOWWx5XdQtlRU8V3c4i/rx2fsZlmlbA3aJOE+
e7AyAAbn0PpuN56m7XtsV+TkTnT5m7jpehYMbQpxQAzmzCNymC+rIMS7fmhCWVyL
WtyHvH2iS6Uj/C2nNp46k9PY/6d/kpk2dUJXlmoqJQG0694zmVMo84q45o+P3+qA
9hs84Lw4oLBbG8jmOlzuqMRb2PsEsm23eVkE8QUvvKaeHivjMfj5ShCu7e3MRe4g
BdZId2iAMyCSQURpEEBO3CLH9ffMNjxNR15qrRZ5r6oKajUes/x/FH7PX0zioSr1
XEGMTPxzJBmVPF2X4KInO+26UvKd9c1nTuSC4UaQTBcwnfysj/J2aKAZq/W7UO2B
Ae4IEGyk9pWAn6SARGdk7LU7qMyWLV9MY7VWAArF6zq+aS7/vEJ07mN31KmS1JX1
aDxxoemJzsLtUch0NF2X9nLAF2mcrLHCcKqxpRuWHK3Y/9pQrgg4iA6+KSXISRZZ
QRLfjDIO22o7Z7lOoIPMHdcJqg8XCzzY6Is2mTgDqh01O+1t4MMXJc8eScX6sJ0G
r2Ya7w1ymndZyHAi/QaynKefV0brG8mGHiWccWoobZEvZmBfdyUxDFRA6a4autTQ
F+bsFr7dwOHI9Xli/mE2Q0hxSBHf2IBfQOeeHNIQvCM8mMPhkpAX3v/JAk4Azlih
ZLLpzskyzHPEYalguZRAjPnL6Wf4C0z+JOoHvc2ucrRLRD5xPV2GXpdj5nX3Z7Fz
SnODWZTGBmb6Jc89GrfFbo4UaNqsNLdXVezUA0ifoeRu8l/Y6oZQWTwujH1d+y3+
LvhrmyBr4P3Fcn9KjjksiSjgrSh+exvfQ3bm0rcZln+5wubbS4tr8MOhrUwXg1Ny
jDyQdOHzZLt62wt+V2IukaNohFVxoYfWaGgGZLUA/flMskiheu3+m+m82FMlxfqa
zYu1MFoSSG7xgRhQ+h0xSLJYD57zj0d18TOSKwa90Yojx9k34sqLFJ+iRhBRyoWY
GYQ+O84QlZ4vqVkLWNFczK17FuhGQ9AzUN02rkX9JtLD2QYCYzrrK0xqlGx62v/5
WIkTa/vnR1TS1lqeC1zGUkhY4labLigD5B+rKZxWHYbNJY97iOppVsFbfKvk0hoE
Q/60vnYpdk7rm4TCuhpmOUSC+uInA9hTCBeBT984w3xOMwj+7jGXLdugx4Ei8CVN
+iomeL2L2edauKQb7LK0LkQZPIPIMHuh4oLauct/emkT12q0ZUlMZFuHDDDfQqP1
UbHA6l669ULVOLwr71vTd3HPm3pjXDQU38H952xIcBL6f6TKAgjWZJBawQ4edvTY
fAHuuNxS7c95qDozlFn/dHX8EpVdgwQjlCzja7YQAsXeyK4pAVxnYigNvvJviSFD
UVY42wENhqwSCi6VxxqnYludLogBHSdBUX8A8zyE+lyPnyfoyO2u0A9QxwkMnWwv
SiHfrN3tFCO0PwduFbCUitmqHL/YC7n6v/ZWFj6L+/CqWs94fmQ4QgZHYF/GBecB
GdkBn2TNjaZUpWkr4YdZMypiJKwwONheS7dtro9wSXo7YZ2KZYEfbbICMXhP1RWU
s5xBsda7KWhYFMUddy3DJlV8GHPZiv3XRuqgOhCSs4lC7jG0vajEm6YsLoJUOG6W
EfDKZTSMPRrxYwuEHnuEy8aUOIpoVOvKB2S1jQE5f6xy1/iSYmeAyMiW+1IJ/hsI
F11keXJQ1sTox5pbiH7321R1IHsjK1gEgmcaVvraYaGuxDTk3jS7qnm8rzwspKwg
n1PBbNlp5WoGtMbcpACTmLscfC4lTmvRyBCYb7bd54E9jEPhQ5erUHTckI1l0eb1
m35K843ji7vJ+nCvFQjYotH0Oa9r+G4KdzUK83YTg0PkbwuQz7PF+1y+51qcJiJ1
PufAjYMDe5nFpexLwQXoPFWtHt4ZoSQmm+hN3DEW5mLhDpCG8E7N4fMdsQNCbPTZ
MwheJiDUI/uM/YNud5jMoYUEmHSb8nlssAlfGICRHN2w5b//4lm71kTFP81pfgaa
gHvrlWRDn46atRKuVuk02ZbdCG7ANaYOUbl0RLb1oeYKeXBRvML+6IEE7D/FpEt9
Lo+ZpNM/jrfilDCp5IijwYRtjgyrUen39o5VAJ2S6MjcGRKXw1a2Irszaxjg+0Dt
IbUBBZboEQ2D084bV6bkn4tgxizcGzbJqaIQKBGkXh1JD4avOadIK/puUriPxBog
vMFcpRb7IctVLW9tYwgcCwg3vUQBcgMKfymJ943uCC+7fP3NaF5KQcCtEu5vZYeW
S6zLfd918dxSjtdc+w16X6kQNhi8BjaVLn7t4kBrD0jhJzYE/gNW88OrU/lfVTMY
CwHNHcNs4C0gil+1OXGPypOV9uviab/oAKINmMLFOtQdcCvDM/WRezuuHRt56SBk
4UPqie8TEbFmMOJP3rqhd1RLrYrGJChhfT7Cuh6Si18EhJBz6j7FXLG4n+gpi4I1
ZdGQtAinl9xpoYF/p89FvrzFJwOjCpYTvcn9Hpo611tiew/7Lfn108maS8HiSeQe
raoxqjw9rdG394FcE2gzkulOjYxqU2mNr0OSJ9qRIQpN1VbI4QyY/AZIpDww3QK3
V5ZHrRzJzowYqPvWVDto+Ie++ToPS/DMGxdfeC7JYXVDNvWNP3ClGhHcd0esuqOQ
Rl/k41xOaOUww0D5T1/Wy57LFOHEeHnNyNenAlKtYdeleaZaSCQECFpJIl+ffxlO
bFeZtHMLOudAaj9BKw9+KZMK/ldSp3+7AwNqhZwC760XqUwkn/+PwvIf4qoRxMtP
z7EdWHT6TJrRcB3Lj5lLc015JNm5S3WRiVoXY1kLajgzHG6tucMqO/XhepBqOKzC
yYMX5gIwjaXIpBR8iI2iK7SoUcn6rIEy5UO6gH61oJsR1pHI4eBVOgPoBJBRtRZV
disshAXmAGAZ/hBVnjxYXXrCMWXltNQvgFOXiE30biKguJKOEk7UjuUtlp/ZqhHr
ezUCeS0BbVjr/740OuDrcf1KFi/dQZ8VSj1yUwYUN0+s9IH/0dwcK6YFVQ4JrU0Y
uBsd58P65pxCD7R3iGGg0YpDy1Ez+wI25wKc7NBwjKgDpPgZ/FYAVkshRpQPnTK2
kj0LzBnPNtJC6KLygfhZ5OohXOB3HEGFszDSL6xNndslOwo1t8/Jlb2FktDZ1HiF
38AtnkaYtBzyK4z+fwOZVYYsMpKEvDILrWkBrj9wNHjA8/aTKO4NtVdtZLJfaHPU
rVZOv9FMKTOqXXImp7hOzFDqiPY3Mu4UUuW1ILgxyod5g1ZYhvB/4ghFZJIzGT9F
tu6krzgP2Ui6bM96b+mdylSagUdgXlnv4FLkRFm8XTz3KDUYNzd8XSx96DysdN7e
LKWG1uJvl8ZGwIj9ezDuGTXBHjUiyTtx7QT+8PAy/nxCzkGN2pP1DsQJAZvLUrvd
o9jMKrDcpOBuEerIPpmMP7Mq87/5sD06EWXhMTHWaS9CZk93EF2Opaqxlz5AmPcR
DEjole/JdLP5qn65B/KkeHY7R3RkMn72zGlN2khrbcJnvspRKiOdzXplYzenmeNP
vnmP8pZzImDxjlaDT530x5xabqRha5dQR7Rrm6WoAEpBMd+9fKWwHWpthE16TzI1
JLgK12eakNOU+V5PTmeFjFlhm7iCz2YlmHv4iB5R9I7OvuN5KCIEp/uhN/NNgELf
NphHq5zU94PaLxTZB6pb+zMJY77c7ihUDcMapKqB6NbyU+V8g8iY5/B2OiUU5Yiv
mlfKLggiuznzFsYDFKhBr02QAH8NUFaR5y64deDnnHQYO5zU4oNr6Y6AeSvgU3E+
ToFGl7Dp4MjRpa15QydYkMDzsYHDQkEnkFHLZqUuuN+q4i0kXzRq6dGP2YsmRVCo
JHQL+ZBTMo7CB1siu8+0WgRlssauU+Xt2pAUWfjgHJnXN0+jYQmGfFLNYHsdxwng
aLE8/cyPx0S/7As5lnVDqc1BjqIrmPSkp+nr2dLN0EPqkkrlbpNq9wJFeZGGQ/WR
H7jtwNTGlFZyxZ1MDq5x7CdX8xRVsT+++aB3E/ZmlPNOeTCI9FsMSBtsO1WXJm7o
N2o2/u+fRw0oSwcYYxd80I9pBS0nxVb5dDNLLn7qa4gWlei5pwX/gc+UPJwI4mZ0
WFfjHKADt6Nl6i+SPFvg88AeyBw73IdycEYUQBLQ1DVqR9sa/v9axnpgAcmHMhY9
8MZj1r2dgrl1AD7WjCZRrhqwmZ7ujwZg5+A3qT/5YMamudxgTlOalq0WvO3MIVI7
t+zh3MOHAdZdxhWyFVKml6R+r4vGGTZLPmBDRUzUTlfLqOCqfm/u5y9AnzwQChK8
lCGjCuHW6AMNpU7cjcYeqykh1dYo4kZ9XsTxVqbTVKzmiImQktNN1C/cwtvLo/BZ
9SlVfVbeEo0wlVjStwnUsaUJQOOemBN31KqyNbZtNdQewEBbnxTIWJONSmRo4D5G
qquJF+4KTwEmS4Mq+6dhzzJNOG9Rd5jw6itMrj0riaG7E1V7TD4kNVBOP5Y0PvBC
9g6LJw1o1AmfqEyYj/vshhoxtkUjRaXwJTXfHc+8HGzvnuFRmjwaBQyPbR1crExD
nmPCdW0gvY+hAOliM0PGePESfkeSUL63RyzMusWc8CZ+8/KWjJkxVT5fpPOy4YJu
Ac4Liw7wPdQBy/jzH874dViA4LVwOxPSNXaiQzCfOOcAj3gMmumzW5sSoPM5rW1e
fhxKXJOnD12GUF6gJfI6fBKdXE8wXHbT+lBIuekax5e2mstKP3wsdKtu1w6cloLe
jPTWSmWUrFFJMfmIaknQ6e7KMoz57T8A2EnQHc6FHqzpl8iZkFxNGWRIB5crGQrk
BP/o3r0asx7pX9rwckWeUBBu2PBbA7nI+lnexKxVxnCHK4bGYQTNhJS8VDk1bHDK
FXQTIMkbycfVFoZAKbPG7PcHYlBE+Ucuzv30y+m5IlhE0E2C8B6aDGPPvuQGXmRX
DTmOG4sui3fzH/4EYsIJGRYkCtM9TO4A8kR4+RDWnQ75AxVXUvLximeK05XFLkyr
zSrOKbIQnAlgY9J+mq3tBtznwUfEWBmpOZMc9/i+rZ5smoFD1L6YLlP/dKjATvHB
iTa2cK617qfPyFnvr8cwvWtJtooPxCQvKadGSKjPrpLIo1tRryI+pQ+GX1FDf9dq
JSytV2p3rcYyBF2qTwfv7KzFA6I5EGVgOD8K5vYVlLAqYr174/D+03T0zc7cuTl8
DaalOTiLtzfGG51vMRAECSXCj8xlUa/XY3A8FmGDwAw+HRJ28ciFxgI+NisHPxLl
NCdT+K0dLEEguLOku3zqcsMK9zJ34BUhZecfE5ejH99vYTwOViSjSNzTaP4v1BPe
bycJAiHPJLRYUTf/g3CXMWILEga4ei8x/RgC0sbsiep0O1g/Oyiq7in/hQw/V5Vk
IoKJyx5AXGsi1hyECOl/ZVAv7z+OhY9KGpCjAHNI/GSdHIZV8rq10k7qcOgyafxU
zyYRBEVPyE0lsBmNz4UqAHJp1u9M8fcceYVDwwvvcBsrxrbFI/wAjkaVOpeXtTD/
S7CRE0+AzD4Y/RpdPJpVuVpVmIL9g0/O6YMF8uigIC34LrDk3N859zrwvmLnwvM2
/wcuxnxmI3hLuxR9A4MdbRZtsIqN4etdfJDAl4QnQfystVIygS4ouczZt+4uPctS
DbjR82yW2uDE7GtmrNs9icmR9uy0CQxNEMiwEWauAwiq4qyKEY++vjj7ebNFeQg/
JgvW5kttoprMtvSLeuZI22roMBR9xkJmoJfjhtNzOwopVL/BScDJi9UWjc7bxHDF
8ebaE+N1ef9Z1izRFRkpOZ9LnM1SDQaEus7pC5IqA1P1lRdFVsoUnvH0yJ02mAPH
NPlW95onTFJvsc/YwhPOtVA1NoRawZGwzDRo0RBznNxGl75oW4+tZ9MpyvIs+weV
DnQHWXoX9Bdy/+jbqyUR1ZAF6IM7ZmUSL2QP5LAwlhZkJPyktOs9Ee2z6DcIVga0
p/4MnJ1gmVhhblD+x4CtjfrVuE3e8IdY9YMhIv0c8P7hgxeXLM8u6gmjSz2vAkZC
8r/I1vs2GvL5BrhDg52apCL6oNLE5hW+3hPqVnJpTUCvZMdTXhzuzIVCj4uqhize
F6FENCu4xDkgcPxw45vvgqmmtU9EzbLP0e++ylZ8d2joHvbzGvL8wbgPi06g0RN+
6nRuPFx8CLHewCptO5rShjTYulIFGfHjBrTgeHpQN8AQh0qHrLgzMpaq/cod0HHs
5HTGmS5BR+hC2Cr0IGCFXG6HAhIOmsHaTr4i/Xo7XpAFxc/KFAp+7/vHjH65/4jZ
ToJxABmjmxUCHWTMy7qEx7Kk0/U4TCHh5EuX3dN7fz6RBdSkdoyYyPHkmkzvymTS
asMNWWK7RYoRU5WElZuYupgkfcWM4zvrGEEblsnXY9byehXFXIdyjjhr2NcvRMKk
h9GJyusV4sZc3srEM+76hjIW2HpjoMsVACvyouNI0Z0bPQ+AD+/XFmEd4VnTgZ7j
ulFXQ8Ca2vXr2cchQDTGbCGMxt4iVILRlIgqFWK1vubfiRLvH9Ju87ZjPPxusXeR
+MlwCs5DjLnbeCg+aZqpnqsQkHvtEBJYIEJg7i0bNrNNypDopo55sYn75+0Oa1h3
4Uh2ragS+Oun+7+kjqy4M3sLkY8qjzoK1RSkIw6tOsa+7iZrL2nrgw+Mbt6maPD1
aH0DCctMr6IGVMW9yv6kQFrmlz3P7JVth9ZxfgrI6wKLY+uQ8A80hFSqpEUeyLKk
wibzPlPEQvzqXXN6NH9GHgxO/iVVq2lI6oMDwDhpO+DhM8+2KHG2JyJ4fa9qLda7
SvXqQrCUQjaP6XxUhdD1s+eSYbdx1XFPdPUkt8YPFEuPMPJOWxpKLkDOuKX/mpQQ
eGGOfPUOmB/gSRM53Kad8gWDZrbDvCfQKG9qJp0OFKSZaC2+M11k7uo3hr+ox+YB
Jblg/T6ARhRrxHYE0N+pa8oMHQeUG/DCYZKFlpHlSELw6rGzufJP2TEMKroj8ulL
IEtg0TUCWpRyT9C7ovj1eyfYpKrNewEW0/FMgfDB/7C4L9Ob5FcMLbu8jECnCwg9
We0v0rPgjC/XUfyW6PDX+gmZS0Pyq6/l/UeW68ptrEYK9NZQChLsoLnp33CRXdBa
z6n82jvoP9wD6p9TG7axMS1FsxNwdv95CublzaGXb6HyYo34TJtUFWzsXhkGBw89
OC4S92aLSN0ebpeheziCrlsg8hdKmIm/QbuzFSRkxc04EFuCxV1P3xe6uk0HPI3V
ro31dbnrVhGFvrEVl+7/vG/L9lYy16o9tvHPDuTeco9sV54xtQmPUFUHUoDyUFe7
uYfhnQq+0Mh4ohdww3VcXE49hR2X0cd7AGdcT72Q8kpxmeqs7iww0kROy7VY7Eli
42UhMA4/1JO/QT4b9rIRJkYHW6YJ9JRKjUsgXvFfZATv2wpQi+p7RHOtzbh+IPw3
6c1mqCMCS7S95sDz3HgnIdP2MXe6KaIzH7aaoPa+5RVvWPo6q7HXnVUaPTg2Ouy5
FoTKtIgsn1TMRBPaLRkq6lKvM5fZQR7HUvYmJp7pXf+YTOQa6ppv/nD0hO4ors+e
ddeOKsPTfvTsdx/SLSQdM6EoPnoIN4/b6hP2x/GuJAIBFYZsl6WCZgTite48SDDk
5xV4doVx2XQGD6sFBXZ9YvbjMRUcF02jtInxk8xAPsvDO+m8tZ7Bw2Q5RWpxc1r+
tv+5OwB3Rls1/V8k6AJ357vMxjrDp+zEPktwBr8KUv1Z8tkIdrEPOhcIASf058N6
uJgYjPYu528upA4tj8iAektu29cYRvJqprvBp8KGp1lFTqEUm0PmavnzRscvB1OZ
6p6WTdnuB9LRDfD6ZJy/60Fe3zqQybjg+DvcChwEMKM5hMIjGGQi96s7ClT0T3mv
+tRW72hHfJcyHNA9dZiTSDy+o+wFFBQsQBsLHBuvLkDlIVlXvmynHTd3Z72eG1Eh
XYt6rKOeX+fMllhEGPj5ndAibTsXxaAddFYMHqC74JGU67a0PcFjQSrbf+CPwOcd
5ZCizjcF3Xi/p0fwcYcFLIPh4wq1UnQMmj4ejBdJpMO8G9MA9iseYNmDtUh2it1u
JWzyFOAR3wwzPkK5eZOsA8X5eWFGSZdTlpgQTdz/CNzKUAEb37W8H7daoEPbnfH3
WtGJE+IeeyH5zS0hqCZ17m7mW8Ue0bSe7p8SZEHXQqgevXV9XbiVGsVgRzk5Mi7I
T1+6zB1FwevOBn3XlbpZfDrJvllGzOtFqLsEIgNn5RDWyYpS2xZ94HFH+KL/z4ki
y3lRMjI45j9hQEnWF6nquOvYGhA1H7+OFAwdBuGccojMP/obQzcYjLrX0WLBy9bp
3l36V0gPbz2e+KMgyYP5Rqrc4Bhc1gM6YziBr7H4/5Av95r2LLbaHOuRafMcmyoF
2s9y8IVE1BXab6xBY9gHzkxSk4uHCPqaILPWtapT6KfKD4AZlRtY1NV6S2x3SKqc
+RsGDn0qUd3MJo57hhXEXqKYJKZka2Cu688FSDwlxarejR7sADC5QPd85dMSCVxw
B0f65KiqVjGxyKdHG51iDbhW4Hm5KIRtFYphAEtnrFaRes7259G/axrWHnERKVYa
o4t//hxgCa+2u+7gGCa1II4b6k1Yzj9tk9CGsMXx2+v0Pwp78AElXNU6BmZFfofI
UVtMYlIKVbMsYZFsLmsi5topN0tfUoUu0AwkCcIzxG7C4qcDWOeKYb/Lz5+GSCuN
DgOIl0zoTJvPMQL8+WEhFxqoQUZpG/B8/Pn1fRaTclonMwO092g0YZ19Fj3/H1s/
ELL4S1xP8Ru+Dbvd9TcJiFhJhA0jf5jXNk9gePV0h0rHBQ7WpQzGVyaTh9SU7vfv
QtqA/7i+apwGk5NJj+40FaC0ItVoZnMMhCBUZTFF7Q9jOnHTJVzsp9Zg9AafIK44
MskAI+eCdNqt2D8PRbJ6EKPUGOvm8/+qDFu8DgqD2jFGis53CrLmrR/3hDyg6Wfq
PVAKlceZyBKrjmZGLbc0/G9D80jN5FjMvgi5uiKl89OZKJxAum+P2makNh7tj5Bk
Q04ZHmrRw0CpiAF3OjIAnJ542TPm1MCGYynWquu1Xbay0qzCAWCcl4RyQu4gmCjA
o2Pv/f2zyYkCalcS2F4y2qj+qxrCEqi4TsYHJRqd5PtFP/C7chdt+bI33h5yKRGS
jalxnuZdI9kp/nxp2crfQiUIpsSZn1wJ9YnK+N85dvbvH5nJrWUDL8vnTYsVJEGT
A+FHBoVP23nVAVUPy2LFaRUFkjTjYJgHOC0WuyL8k5b9q5WtMQDVq9mIwaxIGqk3
rCs7NN5aI78QNjo33+fptpHOVbHon++211QhqVeguGL/w9CZ9SODMAoa6RFBz6fc
tVleZSlFryBddfuPCVl19ehHUuuFNumStYUZOYEutVcyQDPV6JxfbAJRXea/njPM
YiJL6elELY1s1OP5HlZoyiLVSmwK39a3J318oaFkMcUYZCdNxES/TFGyKAvdNeMB
+uImrduM/su0exYwsaZh+gQYawocNW5YCui8nLyGqc3Y3rTGl+1TlhFJzIvHnzQy
uy+Cp3CAB8ztSivXJNupU7PTVF47hy0ccHynQQ+tU9/CZjDpqdL+TYn2y8Fr08Lx
RivzfXuGaqk6WGw6GGEI2t/xFhhU1zOStQ8c4I7uLfjHKjULFHoIBYSwpoxzwBtb
BaPh38NZV1z4OryStkUQJRxxOADADoHEmQ4HfJIbmqvzFnG1bEPBswBZ99l1xpSm
+t9SIt+6Ig+Gba97jXZl0wN0xFkUow7h5O+Yg6z43aFA5QsYq7Jtvl+tL4/a/2gu
S+ffAhJ2Abjgu2uqpO+EcjAmbUWQUwRSKNmoSA3huxBW/Maj2K0hfrJ1Abv9bagK
+eehHV9oVpJYY532RKRj0viM14jgkGCffi5aA8YqrFIvygxIofvVvlWONDXwAXY8
Vr4f5Xw3U+DSTJSgALfUxCRGwYPlzjKWfsoJ86sBBhXvSuGJnXW3PCIC+LqyZEyr
69gY/dxX6y7ePDsduexPgCQZbNRFVmSIzJaAiy3ZXEAn+4+YT0ew21AZjB/VkZgJ
mGBrGDhvbTZlmFAa2CEksKkLY8AOpwowaq+5W8EUhi199wClFE/XazWgXLbJ40/Q
ExeVRUDUD3w/wTDs8q9we8sxBUjsGREpJEdhIlz+k5GFfTYwmg5aGbt7q+6KyPhE
XmT9AcJWeSSjwEGza3xaMwParWBXRfSbipre9jtYMz2zKglwx+cb3lejyc8i6UI1
SOi7da09XYfcKUAI5LAd6I5KV/D7p3DWrLJ6l9IJjxZtXZ7PUxO7I0ztCoDbzktT
zsGyzBP6qW9aiS6HePUv30PKdZRIPy95pxqrYMxYbQltXgv++qoDTPfa6QGzplEo
ih7M3cvy5KyWJXvdmXE5anFmLvCaX1pQL637+bXPH7rkRD7M9UIcAqZ/uC+9liuo
mkhg6rKYk3SbgMOABV46+tKmCdq1QGbv75gdQQ3lCw/OlwM8Q2xmlg/SM3KzQ7rT
E0UvrDiY4JrbUVkCA5I4FH4OgZ76vYv9AZNawDDGyRQ07KcpawrbrLNe6KGBE+Mh
vdhMHvbtBx+A26ndBo0hkhysVhcm1l9+iEFYAdkeLmExnl+WY7tnubjI7CFqRDfN
FWbQYr/FIn6T4dxkcRwYyTZjrUw+jMCOhX2wzT2WGfTee2SXXaqMqDcDWh4kW9ec
Ozvbiu9he6ufFnmNpObciUKP600zQqOEM2R4LwgAQcFegCeLBnwA3RpgeNxjLvTL
082T/Cpv+8KHZ/7VeiFhmAE9KiJLXYTVPRegvN0dKs6z0ZtALgCugRO0/b9t+IjI
SoYKGxuHLdATzd42hpxgS4tnm11iWPPHEw5BaWw8KjnZXX6KDkjIVzh8d2YtCfvY
SZ+l9VB9H8yC0vdhx2zOchJ0N7ZDtwDkWge296VohjwhxvaoOo2JmTU+ZrO+WRKs
6eBvTV15nQ/55xPLyE9EQpK3bOfsl2/GekNeV4C7gnIQsSw04OripcFST69tLZXP
yKl2Zv2QB6JKGO5wVPbSawnlGt0UWDszMFLuCN569zwTnvMtTU2PWqxBToJhb9V1
+vFTm2tDzZbYnKDj9vxMc6d+UMe93GDUJnO6S9J5Xw91dHjLovagblUVJsGaovlq
n+PCQ5xdQ/jhP6xSR9jz8S6G7aAwLT70LU7tHzwAkf0yYaDZDr5v+lacga8bve0S
UWzoy/Ipfm4DcemqW5823b4DaTagrixfMfHDDaDxB94hq/QxeMImaqfwC9RNbnbJ
dXMlrbaGB4fyCV16iEQh1BN8XT5LbEfYBkFpRdBsOlN7VKXoah4NtICPF43jkOFM
E0IcZkxCztmF80smkUtBfDLSx2KL+xDQMwy5ZlYD0qN79HN5vNCUzhkQMxs6KlAg
Q9Ieu87V0qf+JpfCjccSeuoI6SsfWGozG/GWmf/i2vCB8kWu9FYO7SN3z9oGAs5j
q+W0KJqiz+Vrupw55Hxkkq/gLdVyY67hIHTcCFpx+vXhb0LEIONR2o8p4NwEBnxN
TI5kdyMG65jfjbrCrSuGXGae5pdEVOojrBybvsxpNTYZoJYsHYSE2guXGkSIh6xo
Mzv+8Lcm/EKF5difMyl0mg+ViYzltH2qZsAwoY9iD3DITd1wMxrXerww/VTfjfCt
pFjitP1gmiBs4fGedphW+KewvR3wU5lWVFAD1UOSWB1mVLuU03Pr+BdJjASspHfM
Y3IGRrJ1p4kwheXvZErrxU7kcnjLG5e1f2ek55UtwjvR8u45fIbtrA7SNXRfgvkP
9bFaUp747hTKjt4uIS44z55j5XeaqaH1vKk4Sfat8cQJg6WWhRJjddDpoI2sS1Qq
zGawdrGDUJVHrgBsZi/pqBwuDoMg0kLpS95/vLINk6DE53AQTxBTVYpXlgixGE4B
MZ5HvvPS0A3mHVRcil1HzV7h/sd8StaM2XiDodl9FyLnwIaF4rC4MfOBOAQczEz6
q++Sa6IPjXN5XM/8x9GybHDIC9gW7ThJSOoM1W/g2M1TqC/G9S7sOcvUr9JURFLM
M7Id1d/XEES3klmFPz8v2lcUaJaeTyUgQ6XbiLbASLqWO4t/avyuQgMT27XtxGxK
w0KAIIr3w8LOfhuV3vxXRXjE6EZHOFskweM+ATQWM/jMp1y1NxyP34nFi8ucEHAd
1v063CU9KwuwmmEpUrMwR+h+/4DgCHbfuKi3Nkp4SnNGRZUOkOYmLXBaCE8p3jdo
SCB4aXeLauOmY0xPwqUssRIe9iEG2ovB6vvztwn6pbI0OqLCokEeSh5mowz00wFa
I9aX3maabqkqHASP9ujRLFjtbQ00k1G5zxug0JCBb5Dr624Lux/OOewd+nE+e6KE
pkSj5Soi+vuX+05S8Y61S+Ta0QkoZvUVF28oDRfGuKtrLHk4Ha8QlH/xVe03ZoqY
GQlgle+wGCF28lg0C1ExPCouv+cm2EZ4VKotvzXOulhDrWbc6Giaw+9YouVTRqI+
ou8vJHxoNLIDQs+WkcWuS70xuPPVIEcg1iEtqo0oXte7EHqEM0oOTDws0yOj6V6O
nXscWehRVNTsrsP2as0PwocTasNFXXtHAkjDUa844oQKE6pOcf7E8Ie6M2hrl9Jf
vgk8QM1RnuhvibtQHYo6dipHYSBJlGpHGCNWDPuOWngQ5LNUiHLKGZ9qGe7qdLUp
OGUAVv4/tduM539Ex8gIUE9KEc/7Zh+mgTauBjKwikJqP0pq0XLflpGEVRnPZGwe
4Tw0P7SxQQPmcypDj4EzsQS/cof/ETYMJCWoODrLMr0MCKcB2BuiEYZeguXVy34r
NtaWNLnSoVpRc5qF4dAh3v8LbVyijZCUXW/AVuXVb3B505/H3RaBu5nXRo1TV5mz
5RxwkMunhJyvwdtGJ7jCvQdKwMNWWMPFshSpjtaRlX/Swwhnff0IR40snQnv6mQX
YhB03lZAF8PsQfN0lrN5ZQHZREoxmXaN0dljcvkxop1OtwL2nHZcQJXE/wAPPka9
/N1DkPKbtGo2ODK+B41tlIHDXvkusGaSAl95mEoHxn84yv4IelSOeAaBYQ6iqbWw
BoYQyJtV4aXKYgeC2RyKX/ctP2ycz3j3b8FNAdQN7BXXYzJM9Twuqzw2kNFqKNtp
2AofAxQKcLi1CoYMGYRvMsNZmeT01GkhZPh+bKTYNscDXMAWA6VeVU1uTl6unqRo
tn0FzlMma+gzjNvBB7gGVtN7TegjycqdwxyUt/Ou47YPMx4GH9iDI5qFtcdsYG4Z
QJvkcHQjpRtpXzomk/CKI4CATm5ZUH9wsbLXqaBRyZZknnAKhDobQWDz5wxun3LV
gbr2OXdM7GeAQ8HfRWYUKO8W6zV/yzJfqtMP1IuT/jEzhFcROUyxvw13gvJxlRRz
z8TY3vKGs1CJW3U2BgKIyCu+S2cksTmJ4kVFvO9azHQnAFUXgM+jL4dxyziIrFG+
oiLR497USrZdCo0cp5NQmaVq9MynpAwjudoWMY9Ze8UvRj3vx8vomrFW0vJ0fZba
hisFt6QrbmB6YVSs3gG1GcCmkd2zAPDb8xrmjgeN8jQmURomu3AKIi9fkBkK2DbX
bcEc4nZ9pP2rkAM0EjAw90GJFCeWN7ufFMx/QYKFOymyQrZPaboaqpTttZm2VWXh
rlFRwJrBGZk0lcyf2MLvTPZHYmvmzO3+M9DC6ZPgEc6ZxcdbSsNZQ7Nqb7oOtFWG
fj2QPLIfHmVffJeJfTRZNmsCoFfyLuqW91+rHoyQFZtJ/0QxRheO+Q4+iY1otm8q
irbeH3B+/pIQcu58Th0ieRcssUAWl1nRs/HdswAj9HESWyUmVeT1VRjcL4j0Ub++
Fxf66sEDuHDfYT1V+M8fL/+1j3iTGOp8qkHBnuz2WLN+05wfbkssRVEVu0692Im7
YJXR/LQd7/KKOf9Qxc4Rid/iRbo3LnFGfiFDnvUiPz3Xb2+bpsDcqX1q0KL53qAm
KC5YU7pBYe7RqAas4Zdbg7OxWXbhqjHd7jsy8HsiXMZfeFtYhXqvaeEQ9bacuVnA
UHz4p5xQ2Av4sxShnt4xiEkNdTi8gryYg+mkvhD1wAbRrIfbBJAj5TJg9kyUBk7u
cyCzVFJ7ewRoe81QLsNJNVqG552hzLz8UZMud3ENr9MXLQqy8kU93PJ/qgxT4D5p
nRimb7FMmNVSqWcikYM3qJ76GjmTV5cNKoyIfZyE+uMdASn3+bM7jctL1+ErOj08
JgKeNUt4A63fnI33gefYKDgrwzRY3MLBKJy8Db3NAPKVA5o1rskN+T8GRkxzgnU2
4+PWwcgKYiw16ZcOfZvtLaNFe/G8Quq8ATOctv/QIedWTvtqhJ5jDVbBuKimby8o
ykzlWsuDoKPrmTMHcM4Jc+XE7o9zT9Dhp9H0DRZmJSNklckXAocxMgDjcmKTBVnk
DVGLrz7gtUb/nlTV5r6+VVMLz3vtT32IU2GxzFHpRBEWUCwhd9aLRr8FgBPFW5/g
ragzO0AoufKWTT2ClXGvBx6fqxl1gMoWCxyu8/KquKjdpfUeBQ8z5EEAz/t6zkZm
WKmCTC0cReXhwZPDKgLF7FkWtDESKCgwKHJbWLHVglOKFXODJt9hKv6JYLwAMgET
EsuboV3veKKpjcR1Y0G0fukCogPUYYJc1XTFrM85PDApgIpj5qmVyD5f16tpat6W
FCh/xXsLmQqzT3l8NaeLjlFYy4+UU1IxIBlMk49R4hqXM6vd/OSBHYSADgjw1kny
Xh3bjCKjhc/EmjJfBA5shd43iZ2O9nw+wHUvYme5YUFtEsMX45vrdhyOdt8wudiF
0jgaj+DLdiKj88UHDrIo9aNSrTFyW16bVLXwJ2LY09LbrfrxRrRo3YPgUhxioDHI
+iKs1iN6afwOb9oGSpClZ29akzIrXHx88wB0o/tmjDuhqk/x38u2FRB5RtMhF6/y
LWxdNScMRQvBvlTH1dYmfTNAkeI5FS99AgdWsnnsEp9nE0wAZMP8MVMMxqUy/+6f
Gxk05AUGocVLlOsS9w5bvruL5PIu2xH0IA84+7MSDVxaQs0/UwQ7dVtvv7Ati1WP
mnaQyGpGDhN9tGEQgRMrZdx+Bv+xoG6T2d99dxA5Fr2jqtlW/AZvWGW0+6Sm0man
0XMwkRCGe4LPAIxi0YiurRSKkitJR9zgZ2qpM4+wA0UnUDXEqvrO+kHl+s9j1m+W
Cq8ECjm5V8atJeA09i5NVteJAJdkEyKpsNsyYHKY6skVvctjUqU0Pqh1HoGtEuXV
B5TZY20nii0BsUfe/4eC1rO7iq+nU3AiZGay6+exZVlXkGidhuMyWLuprvc0FOyy
Q2x10abgZ9fzkDRlTpa0CZs6X6QNoF7J2P8HgOhxtkKe4YvQJ+C3gLJP2b2mJqfT
x4Us8amJWCAsHb5SAIALCBHsyRPWLwsRoJKEr5y6yX8f81W6L9DUyoHzq2AfP1mT
U0wQcIEQYKMZ7yWKdFJOg34HHy5CDC+Z8Bvx5doJpmMXaI/TtgZ6NnpFIg8gWybh
MroWEMMqjIq/oPZ3NBDp9CYN8azViI79tSeFiSgCpS7yyEPzptqoxdUp4ItC4uay
ANItZwyAx7yFUZStwxfXaJLQ2+quQsea2oukAybB3LxgjOA4nUPaqUVSq+ALj0Kf
bYRGuP7aQn1ziRBJz/HWu7sckyqQXkcD+2RPmvwzcAnC29kNi+kGEEL22bG4n182
zh4DHFBoH4j5C04c9oBEjHq48LLT55ZLJK7hsmji8mX9INZz09VAi+0o5tNWiNHl
sP5/nF+yB4THclWLvuj9o1cpdsf1sN4rr0pRwOb+8i2/nMENZLus3i6sMSEQ1czu
0dM7E7g+bxIHPAjp0Q24fqcJTms4pMTRROzAlNZkSiPUB4U/NsP1yfvd0XIAqduS
WEjVoJ/fU4+EKtNL0+sVg9MDawVYWUYtcRxcDTpkUVhTWaDaFauiCLyh+TAIIMiE
MZCFsn+htB+P5yrF2vAWRWHXaVx9mcS/Yy8I4sxDa6Tr44SPiceDU40cRBkkgt3G
uxlfg3S4dv0QUu/QzQprzoO4GOcoFgmYx0pXaqDDHFt7x9v7V1roQXhb1TFBASdF
mnvdqjrsYjoPIjf+JQmOZWPf8OJaz5YLJRDoPNzrgnf8q8cm2ZzSrQ0GQgk9bjDd
w3Z/PHYQ7cu3odZL+EBpyppe1e2NEFMACy6g5cd/LHEcLnP9avX4V/ZDtSk2bc8z
+G5SEawP93pjXsyNYUHyFuMhG96J3a5YoAV45vkTArIz2hgdunB9K1zutwTat4V1
SxfqYxF6oYGqe5sBtqO5xEwT2RqjLa+sbPKZrDCf/yg5GoxE7/dlE4pCSR+aRnbH
i2wVVwI8MsRF+kTOd/lQQoKQ8Z+6pRlzBsVtAbc88jkR+9v4QinoJSUM42CoQf39
mzTt4mAIvTiF/GVnn4j0+KJp7M6dmiyqLsMTJCrIjUZlD+rw5zfRR+n2YOL8liO0
lQWEB6LVk9+ff9EvSlf2mZ1VmyC5xTBHVP4/qT9LlLIR8aDeeJKLEtjfNQsl8E69
dEYabZkpdlMzkFV61MCQGQeRr604XLyaOIaRL4p2C1UT3PummOdkp8i0l7hW6BCy
VE6kGtwBSsV7YmtrhiLLs20+/bQ99hK2qGM2o3RHedJqdWVOJYPG1aa7Ef+wPSUJ
5QTqllpN+hyFkkQx7nc05sTWFXyXH+blXGSyLfY1811R19nxG6DKBJ/uSvAYW4Hm
DTBfh8pTLQhEOOiybQNa7n6NffqBXdmGrdPiCDoW18RVrShl7i6jlNOsqDdIzzg+
4QwQKq6+qRSbX4MgJZ3gN8VM+Z5Ex48BRvLnZxDcc/SprjLjCgoRSo2/soAoj+bt
HYTj0ChhuGDU6TCF6pKfr27yO5QrK+bDROuQjxelAY+iPtbkdsoGhN8Xx7+go8wq
Bxv6QXhhh4uf3K5F6L1HVg6jDEcH3h/EFjTYk85/C1SIay1m5LoKn8n+EE/QLQb/
QfXI0BQqGb9klIGX+tmF8Kth9YeDSVp2qRoBxO4p9sYXBI3LeE/stVe913Efkk0a
JhrZcaJUzq8IqNpwrlung/aV42U3ExfG/GwfHC+bYpH8rTbazdFt3lfBlDnlE4Nj
KhcrZjcFZVjBtJx8RmXXtUfgXV6UO01zNadjt5kRfVhwwSKXK8cWnAZzqhqqsj/A
xEb8ycV+P/f3D8hq40KDuuaP1/wTsneTz/1dH8sH7PfIfybao74f9daYqU5W2dO1
5i8vLEntpAFbG6IZtb/qXM4Z+ImkAWSjcVFGxGEnPAGhNz1//kM7tS0aVy8s0+AY
ydTqkjfMBuGe+HCZSPRY9L+2emnqOqo5Mo8kfY3GP2ZWJrRHpCzRhf/33O3fZEei
rqzdfz9oNVnQ3nxreNtoBgYZNvW59ecsNpPpe1ji/xw5rlHGU90km7U7diLVX7n8
wmTDzBb0YoIpLOH9DFL2oY6O39T3o5nQWNR2Qev5tmrsMzXQdDAGIdG6ZWgJF6B2
5zo1yqJaFgp8OpUu1FqceW4CdzCwQunkmtoLkd1dayjVK4IR28WJozzt8gjx4ldz
3Tsxq2b80bL7oNWraLWbFqjruGH7xK4FASGEm3zRtJadzFOC6K2wzUz9Lwk1QmF0
Zvy91TreeAo1t4voNrTuowyNLUA4P0uBeFRSxdRb4Lzef+IWXXUqKfmtljAw6Cuv
8JiHSA0Awcb1BgizlLQwzLkzYz9I5ntscOgaMo/EoEpe/YmhF3lRFk2Wpo08CDuA
6yvKDwjDJm/aZJ8a2FC1hqkiNEq9YG8L0t2ICnwWVsKjpY4Qr49gJ+QzWrrO6xIY
lzJRlnr5PhvgTMbiZw5ymkdEs3JUNQ7a5Rg5mUgKx1KhgmPBDUnQotmYRTl1ScW1
oTkzV+XVXU7aIE7VeeLpWh3Sa+RvvE9lClZ+rNiQwd/EWhMdvHEd3KCuIjZA7laG
YdxUvxUV490Hl4OcVEuxABrXiGBtCg/Q/mOC7ri8XnB4d3ikyXzUOyhhOjA74qgM
gkNXIYPpiohfHmS97Gju+chmgpiAM5ZMSOKoDQO4wQz5HDq+MnvZSWr9xqkoUie2
hO0JqZaXlm8HeLjSn/FI0+qInDB3/Ni14L6q6cDiu1F+oBlcun6dz+OX1yZ1aVlG
xRdErOdtHRVMaJkbq0+U0X14v53lQhUYQeNWQaxrhzZaNevwdDzgrh6ZVIF/g5kd
ncfllVJn5EAkCw+imZz0bDKzb06wHwsnVkYDTWCGFcy0xlYyv19JhACgmMxlQAy9
t5UWonXVSBegSTaGyDJ2UqEgMvpVvzVJSesV1ko3FDisPAlUz9KtmmsLTCC/qGw9
BtKb2jjWBh0+1GlU4h/AqVUTISMkXMEXkfnyqGE1mMk8Vww8z0/7uqHrEeQC/9Gs
rgSNrDmmhRE608l5KlzVOuENB1RWSN71FbJQT9D1SAn+D3IioIWOCyDN2RZJ7/X8
RDp19f0tLYg4r3StqXl9z/gm1wNEIwm6fKmdZ2soOS/oOy8CPKlBMYK5hB7/hIEl
eso7B5izg7cu4pUw4tKodmGxD+KlYTwVw/nM5xW6r2Hw/nuH4lAN0K4z5HZJAKK1
qNSS1CY0bliz7BWnWxMjGesYGMlk9xWEjHJIH5JOmQqndf3NfKr8DD8ySg2tEVIy
gDTf0YRUWtkwHfegqQqqHGR1yUh1JlbeDqRX77xEvnvghCzUFoKzS2CCV+3T6aTr
bZ4L0VC8nRe7LmTsefm/nU8Dxrg/caYE29Qhf0m3Tx/T0TbmumaqQXMuf4EAD9e+
man+kF4JZlKRr96kHE1e6jSn+0UCT85dE4ptZCmYQL+TpcEThrp1rojRamqpwwvh
R5BsfQqV8hAvOwbo5GQEoO9pa0jTjMkCCP/82lvlGD6c8bcqc0IchGtBkaTtyZo1
a7dTsfD0g+ioYYHm/kdnYkoQ4LCN9unjT5WwR/a7oNAMTyo23U6lG3/UCFrH1mYL
hgCF8kZym8a6lMm5Z2aADUHsDoS4qVul+InOJgI+KqF5n+UM/Fn69u2Kx4lZlyTE
FiT0ErH2ZCA/sjYBF4gba9jyxHL6pOt+4dhzK+ls8il0tI9ehFEa+egtTIBYZQLO
lx9mpCnn8IXLdR9rznTxJBhDrOu4V29VXukL1IIzv4w2ulvrZWuPuxEPoKnO7QEz
WCdlMQzcZq8fOhpVZX5zPXzPjUUQoMkJ5CRco42n96RQR+XQwoBdVQZ6rd3EWDaw
v9Du6DovQlzERnJ6Uese+vAcZg5OE+6/Ro6qQK+0QbSogMKubqxAuEqx5NO2y4Mm
2mpJR3293VlghaoOFWsGMfXMaF7I+G2viiZsPR98oRpHjRZuvypvrysZpDJcJiNd
XWSVEuxHeuB3RLEicCWM/lSAgN2j1v4sHblYf0ZqZTfMBLkYph79KI+dLynRhqre
HtAJbPZPpmDLt/yq3m2u42UGIlyFSCgHGHkeoqszuEw+CvQQVIyx3u8Swwt+cksU
HU2C7+Ksi9totF+ayaqPCKhnKMjI1lYESjj/Bv5WbHq5cSXwF6oKoi3ze5Zr/qBZ
aikZjeR+0KWq86bXEsAuiyEjxCz9t0xhv5ZKdg98ESrQUzsakjAubPlA8+aRhPj9
6dmhCKvUAgDG1v1Fs1y6sGePFcQaFs6aH2T+wxJV06SrIuMVsjVyo2k3LG7aDPYm
aQYbNftNi8oJTMVzHS/DjaHZHT4PgU7/2idGTA+kpt8zbU6Mah9BZn+0OqOSvbAO
0ihBIS6HoacGI/MhjRxJTSeFYUOYQCJpckfHTpQZ7LAkTrN4aOegXnewzUPoSRcD
EvB2EW9nmJ+KoQ9oTrQqwF7B1Kl6KnQmP8j0RhzQfl4l6ZIGmcIxVVvgrE2WL6v+
b/l1NjUOqblNQjFBoOF4cvLGQr0ak9VK40w+jRIEq3WedveGmn8wkjZEKPjTbAJ7
CSBVX+P3LWzOXJv7jSR5HaccyQM9Fp5jj7lsg5A3KhYjhxt6vdqThoY+SOrb5LmF
0Bv2LBFgh4Zv7b3BaoqrkI+QJaOB4Sp+eqmCbL+6zFICzmT5tmNp/mjAeHJlmDM5
BFnYXFmD6Xjy3JzRLV68Hmn7jRNKNGtmE4RZz13THLf02ZMcPa1lXZ7oZA11GQlv
/5X40rXbHqYAEZcFYl5Kw7MqQoGBnvBJBIIDAqZSNUdutX5BQHiXQMQVgAtRMr6Z
W9P3mYZk6HLL93ydWGkKjPFGhteX0bvkOPu0wmuBOov2CZBzoSCfaTh9hJK9z/Wq
SFWm8BSXwD6dKOlCetLZnh8ZiUvf4lUR6t8rbOT+auWNzPeYBG7OEQ8Dv+ReENQ8
liT6vPM5LpGc8UhH82FHw8jyFFXBeA+PHDoxpXnESAGhRpPcMHqK5/E+Am8Ivm99
S4+TL3wPdN702l410M5E2TzmYVJcd6gwUNk275WuXBMlGS1193k/1vypNNuBupeH
ahbDEg3dQ3Ys/l/wTUH5tHggvlmNeKoS3zuZLeF0v4iO3gnLNJmkEXa4aAdS1t4o
JqYHHVP8Qfte9JXQC0WlZ5aPukFs/KEpRVxheohzdVmIkHv9JdWCB45qFWeAy5tG
6b4b4idzUFuF5XgqLBtk7+cKqaxIa/FXwbkSZAuw4aQm1733nKy9ke7AxiPpF21V
k32uNl19kaTxDKiQOBiDvOFoTxrUEUDaM7GIhMb5k3o6ns7+wtPtYnN7z0EDQvbd
pRE2flIwl1WwhmWjTcDH5PgJQYWa2IaQGmlsOsGtWDK8mh53NPpYWxnwliaPoHIm
eIHxf34vZaCl0Wu/t3Hn3NEXrTi0GboP02ZyhbU86hZlOWGw5iRK0lGJ/7M9L53i
yQarvV5gfZ9vx6I1h3zTO2Ixd4elqZIo1WKzyTYB5gXNoh5/tUrwf0F9L9T7aAhk
PbZVIa0qFomZlkO1CmE7zJEKfjMlCA+jhC2Sl70IH/2i/vi7cnpE9pFTNySwaSaG
PsuHbX5r8mDY4xaNSSZ23hKrcO/6XAMCQAPIY7CcT9S3oAmjqclG9QcQGucxzjaW
eyFO4nB62q5qgjrIQdVDuWJx/Atea9jRzMP1HalvHAJr6QE0qI4kBaVqoXk1SgtJ
tkq++6NHnRFr8cW3QoXz9t2eMKWBGem8sc4Yy7TN76yGWjq9ghHSMgZ/w82FR24a
1VyorKaAMlPMyPxLYdZvwQ8kKWyUemJPJyBylYmcklDf1c/DCaGUxqUCcL2P8gGN
BToq1pcr5ouJOvEUqaHZdaQNzpG32y/sDDP8fbiv+x32hvTS6/9rqtTmbHfcm3G2
ccmpP6RKmN9Kjk4/aktv6eQ562jZGf4JZSMA5x8xJE9yh5kme0Y29mCE4oBvW2D7
PSYDAQXlV1c4tEFpi/1w/k2cMNh/DEAN6gMsH0sS+xtz9iu+nZITHM+AWDzB7Go1
/0eDaUT1lAXAu/1+l8etjFyycnZqm6KwLEhEABGph42Al3kJKeD+9ABmmvlT1bLb
ci1tZuiDD3Y2Uvl0cEct9QJmk5pFjkEMKnQnr+fgLauW4XnVMuXsaw8qTxCAUIG/
Kh4CQpNR45FIwO+BySPAO7zpxtWbQASd9CezmCYSeMu1onZ1z3tXp+VKPQNUXodW
ig3sVqX2+VYFgEAnxoFlADOQzRxj7P9ehI1m50h699jUGd0/FgKNn5yvHieyvI/m
yMH6w40BQSWCbT6nMHknudYzHHzI/c55QnvLtGL/Uzu2s5jAZZfiyI2vQpb91ZLl
XAxF2xIY+FpP610JmsKuOrKxhvYqRJgR24vD7n4UxmehTEucJv6OwVaNqPjZg365
pnXmmy/PPv+PDKQcppn2m8zwjBnhlTvnT6LA9PsZAEqlv+lmB58mW2CPfxLsnP9i
F98aFEisTcEsTRhcfqWlTjXVFzGtZqkTIpAVdIvm5Osl3zFaBraqPkD971iqpZTA
N+xYMV+X7hkShhYHM6Z2qJAp9CxaJlns/L+UKtSPo3DFfKr/52aM/+RZPaU8FzYc
O49P4fVRXJi1C2ZkDZZcqx3eO4uQ18wMRmwR395x0lwjYN9TJE7EG0JlXAJ2nRPv
i5xHRE8aWmY60dsMfAjTaMtMWBuC2sRdeUur3u05SYQuiyt86q5KbPxUj8QsnWi+
DqW+K9Py/y41Cuam8zmuM7kMjbyNa/Q4MxRqshL67aLodZGPiKb2EjcI9k9ooDTz
yTOyQyElnlDo6AOrjYhMTSd9UvniF5cYX5D5VqJkS14nnbzZsQTJn6Okwkz4+b5W
3ac5S/aupv0akZz2u5VvrMGsUzyEE6adkorAjMDU09XmqKHyQRWZo87KfH6YG+Fq
+hvam3zUGvM001Ttem/a6D6B+JGmCni8kSMjh9798yTvaBgVLRugudAS4kwNNKNf
lbTwXsolGsUx4Q9eQ3X8BXdHLk8O70tV0lqAVmxleIVmO5WdoGq9pAo/n9zSrs1q
Ro4+UjaBqSyxTJwArVEaeRe0x6/Y5h49OJbNOhYCfIU9E8+q/bBfc12lueCLcgOh
cI8gL1FkrTWxSPHXAg5vnjtw3akrSj0cynJOLn1E9FTOKFkhsbxW0EAkiEsyw6lp
wblgVS7PgZQMkVYd4V3+spN8HbfhQ1l/MRX6NL32qsJ581KEy8YzWMDzuRImy1ph
0dEI3tz8stNtvPBD5KvAkvPVpfytNsfQzslhMMKli3GwxdIc02uQxjzXMQa+ufjj
W5RPMlgpbgwqqAhFkMihxr6I6ryIOP9ln6eIuzz3Pr9L3WpsHUoRY/tkwmQQ1ND5
9OHMV8erXNpD7w0YQBXg2qsmwmb+5dmn6iaHc4r90/0fXZIhP6kmUEbXaR6Z0wyu
XMwH83oxpQwU5Nh0+2iPBkpRnQra5fcfPsv+/AocsDVGJYtmTj/SUSLBFKEmhmL/
UlGsvSKTKwviEqBfLanelQ2Ggg7nxrNtnHqynNpW0pta29HPXkIG0hz6+meCE0PV
luEjB1VyKGAoX5TOTzWiVzCdjLeohkuzZywzzp8vbF4cb+572RQt+I4pB/KcCuV4
6EhoW0pE+boKm9/nZzkXxclcKntQnhjjbEU1YzT54wRXqWBzF4TTOohJiFz5srfH
kYjbdkORl4MT3oX+rgIsrMmQWIa6g8oiRBP3fdh4WUloYBN9ylKz8A2W6Bc3SqPy
1B+7xz8XA6ea8Oc/uVxuJ+fKW9xhmrCgU3zpOUixLVnTwkwoWv4iAhy0DJ2srmaO
nF5+uM/FbRzPYSUWh/Zl/dYfLSCSX06YdgTOgTXQzuBGv4mu2yPC/1aDr9L9eJ/l
pJeRmslSr9xEJJU5+lhU8pGORkMhwFY4dkBhWcEZa5miAJgsF6BV9q70hAfuMTq0
/JBC0fmVCAEsQS74KR9t6UtBowCPT5s5Tr6Z+PXAlhawhvY0QPq9ur+66v/1Bv0s
j1ILDzgj8A3PTFNx8mde/8jlFwagklD0Sc9iLDjDkVN2BiSpkWXkcRlSTNocpoSo
ze/k9wh4+biIrhZfgT/eiOdb9tY7PHLDR6O4gThaB0RcolSPSCp0PIVqS55Klvto
ilIzkZPBD8eQaMgzosz/ZZmLIGZFhWAK/0kk6UGYOOgUlZ0DfIAxpWbh4Qz0LlPU
/ZA8BKaCR1Oz1tiD3GUGGbhode4q9KMJZdjNp0b0fFBEMY3TRvtFF/XV7sOGTVwL
+Fc3m/94ysx6rPgDC9aJ+U9jbHGPptggbSGALmWONQhmXjNSkvSkjL5ExrEKeN0b
1lNtg9+7mHojjx6bVxm4QXAsbj1wiQjfukJy1daaQP9KJE5KyfK3XlP9ooZgEKeZ
gMxXLPbYcK0CgKn6rToE2sbWrUMPO6E2TOhczU3ffhTvEesQJefcscr83c9dTI1m
1KZ4oqkeC6u/fUiXTH/Q8AOuf+b8/GNXl6CwseoIqKSph3xDXgnWqvl+ralaI7Ac
Y+APSfZmlvMeL4OPSuio4mkT6bnbfK9pNwH2PD9IdX2ZyBsXAWWqJjl5Irw57UOq
MjrwduicNs0aSseX9clVTWrpNQTRI51AgNTxcBwwwzif9Jmm82O28pSBESScV8/L
g5VDZpxJQdoZg/bh9ZF5527wR83/fElcaccBw0casUgX09ThzLLMSU/v+Nng7ysS
CJGoVtorsAyEvhZIwQbKtGETA6sQbHjU1lUbYw7L2cIIvB8ZCWIzMR/hn+OjNxgs
rm9t064lqzARCqYiNzZRNN0xsj4+KhlnRVTUxNmsa3pFfGiuSbEV7UqNumftCnoZ
i7uujVsjS/Y7Ux7f/6ji2N51mSgI/FCFdyyFoYb6yV+rdWa6kSBuhyo5uH5sE6+5
RDLKQz6kRy2GBKBllRPkEPTlUGrg57o8XDDHEMhp1pLM1NlLBW6oHbBLsD2KXIRh
iitPJpvrN0Wcn5f7+WwrtQqpPca3l1d6N52PNMylE4RAvdEtixO46fF5sTnSpvZi
ZwQ1SAr1idJ7EhtedkYaNIlAHF6ha/OseGaqOieBvhd1udAnKJcAkUOUSwUHBO28
6VLxGpt5JQZeRPyTzlsStQltvcVDhuBmGE2vrl3NyanR2Nmy4ZaX4jiATs/T1aKp
EqvTpjWV6rgT3Pldd9V1uCX7FEqkygjN0l7v5PFNKj9EIibw0PpoZ1Sixlxm2zBo
IugN1niqqB3brwY7k0LPVbG6ZC5TxpOFRUJuEpErr9bYLFsx/whq6MVAbzhPIhJW
gwUXObbI6fenyKF29sVRxEg6+2KN9612D4EWBDDR3mtk1rKN6vPmzK6FXeCwkMtx
4rdcS11LyPryH25wZOGVjeJw+xBWAku4mjh/Q3lDKuUAHF9QEknuA7oXcM0oj791
ZTx13t5OEjPacnRAsPaDsXTIyaZuDWoLfO5gaLnAlHd8Hg2nzp4Tk1fyykt4eU48
C+lto7jahjORuDzY7sTKtafhvGOxG9CypVoYPiTBy5LxkV/AUEGSibT4Z9SInbn1
jMNxiyix5CSy9QCOXek52zV8vPvGtK/bvMQFjupBM8ZBq0tRg5xL3lJc9o+/eXWB
HMbTIe4eIpoO9sCm76uI75LQS7FMWXvUdiQVapchxw2EbVb3ZFdg1whZwJBs4H/F
51tWAxhl3ZhhGg4YUSo6EEalQXJUrOAtOz7K2XMRcmYddnrKvW5x2qy5zishdX8s
SZ0aP5siKMo8/9o9FSr7DcLznffs3PkSW8mqYFh1fZrhOGERh+lJsvHlF3GM52R/
0lUy9z6DyZG1KJRCQZea1qxWCdCUtLqG7VmdOXGmHWpnEnM2PMrHvgIOeGnClyvw
fjjvyg0MNVG+mJ1OeCiLoRaijGN47JQn1Fn9Xi3PBmClA1QLLSHa0TPHInSvLPfd
XKz7mDD+iuSyNNbuNfclwV0OJ8quQ91SgWfvtMpst20J70bUChJYldjTFBwUsSTL
TAo3rVJkjUvQFR31TdIJtGVy9Hk4nUr9BbG1tXcq7dIu+qdqavTsX5J7c0Um9lDy
rXZF35bQWpKoSw4x92say9JSEEy3cR0k6u75Uu9wQFvULyDu83TKQjtWR2ERLD9j
78qa1dnOW44oFTKGgHG++hcelmKcnCKXN304sm0fBtPUGsGWTA/L7noB32V0TxgX
fqeGX4JibGr95VIPiuQYujSNY8W5LZwCIuWR4yBhwhSvPv7HGNOMYTYUuQrH2S0L
53cn8DZvC6fPF/7eTbBHdmIOWsHhgBeIAvqFNTBjopFEqEETfgYjSgeCRjN4RNO8
YVnu/yx0+9hzCLq5c9m5dVfvkrW+ulyNWmYAtxdQXTgevRHEiTme8Wsn901BB2ne
4gTz4EWe8JbX3orqfIfhyLXrCaMV+Wf3mfU3DYYfrP7bnnDs8Z3XbJlpBIH9nzYj
zkRpslU3gWtK6/qAk1rtYqer2E/+sQWtQzHXOMIsBM9GN/BiHTYS1yEeln6gO9Ew
1KIFRgZ0YfeIQhKQVvVfYxxLjyPyEcU1t1Ge61WXmAejccVlNaqcNBQKzXvKXtfO
UEMKgFwwRnfuiLJtqROGpqnXAhelJiV9xM6HYQ6maJVlZeAmYCJwETm53uhKvVLa
56R+eEdB4oQ91sHzm21mkFXjfRu91Du46KVR9FHRt0/pYZYo6ams+HTBEFS4IaKP
4voA4nsiC/N+9sQBIQADVSyFOG/va/+7RQKbGiOXXt3IPmts0iAiPSC45Q/rEugL
CqJmNRLKkaaDxCEj12vnjvlrLyVqt/rw35jYF6kf6AWnRaeNP+UrZpQdEvDnQite
Y2769AMphsm53lhOFWWCgLmKAm+UslvZcxcq1SHLDqzohGfKOHeeX6DPjU4ASLsq
05AJA26Hr+8IqLPWHI5CURIVqYdrk7dRixnkBGudmdaL1jywSEq5tX5IH2jIesF6
PWfysAYBF+2R15xB38n2gQ6gXzbze8nw9mIDGMrzy+CGgOJn7kSkCvJbSIkexzbH
UTJ8zPOz5c55ErLtDGZVmvMrzLyxmMY+tbEkCcs9lVqOBQ7WevlbCcjNkDmVfq9Y
559GVe71eg+r9hi3BZUGSmRr0xDkyuOr6ETH7FwE26fQhqmdFbMgU4Sh4vjJec9k
WfjlKNVAzFobmX0/kkMDyNnIpfyrbpPOQecvtotirWoPGDivhTdiP5IxOL0cKyOd
veAf/6waoA1ZcNLzV8it9uKTjslGII6ii4HcZLpeBgOG5C99MTqppnZnjsGNpD9/
KmiecMx4pAAc0+71SAGLE819Wfoz3ydWnjN76dAUM3X8R4hC/fJb4ekzmwZPDqDA
ajizNr4Ta+dj1HWpOsue6TdGpMGUTs5Sg5kY2dnqpXM/b4UxXU3+mw+7wEWw7mcY
NfbUOawn0ssfpjMH1SKXfs1ijb9f162+QckL04XA5GBKNlXW1VFIL4EKnvWOEugc
0FSdf5P0JRd2tIwA0AAyD/NBjTN2odPC96b4I9Rq7A/IopobdgMmnMnz09GkCt9R
6L0lKj1p82ilVubLyrHf+5Tcl5kh82IbQQS7Oc7/VEZrtwU3QBYW6ypIv5jpvzKN
smn/cLDtlKO0lrzu7BwI3zJBYGqwJ+EYzkEOtlAiyv+MUP0S8EgCXaPo/uUGnJ3l
+E4yh8ytnYZVqdMy8Cd8xeUYCcGWO/1kN3KLhlFHmNIUqvwhOvlDVgOPwoX2Uqn9
mt80fVep0Aa6l/Gkgg+ZNY1gImVj5LHZU1s44mf1wrFHp2AdKU1jN1aW5imSuuZY
1fWj1IMsuDIJRh/gCFLf4Ivx6AAm6x8trmPu5baukzcQ62+j6CkVwM11tRUQIqVK
FWuUYW5NXrt3edX1s+AND/VrtR7TLis64fTP38UZFMeYabpOgh/NV3NkpyqXTz+Q
dxu2jlQR7i7z1OvHA8wnCQX6zfOh9L/pEzWttEvXL59f8RXrjb+K4f7t4/mnGh08
qvVg5vHLruv1pO43CHJLiOTp9GNwQovg30PZp4K5n1UUJg7PhRennN+6noHcWcRa
r1lYnxLr/8ZiEGLidQtzh/Yan1wAuGNFiTEvEd/PaBsIkRehLrY3kZz+pxYCOZoh
kyAGQQvow7RoOn9ATpDSGSflGmQdPhzHZT+0XRBQuJyhLUniPAkdfneoa/qMFZau
7XmRL42e7VQjPNuqKM7j1goqqQuvgR03A8eWCBysP3ZYOIe3NK4zJAOtzNtMZ8eO
a0hyUbHQ2r80atnoNgeycrhLHg2nWa+cICA///4TAIZ7FUTau7YJDqUpyOyLA5KA
gv/ncUuHes6IIabXkrA9ggiMGByefK7+fqSnL9PhX2llNhYOrQSyZnSCSaB/u4J3
KgtWX7WgrCdRrOgNsarWpIZlCxz/LGT+gOY/bf3ZnTmid2QhiWo+rIWDCgEsu4bA
iImvFsIwCeMfR5pZMpjL7WH6G2HxQwYV6tg+DJ4aA7FjmYpoVHNOzbOEoIxfrtqS
ibfrxkx5MpneukdqcFLKIN8htsV6N1PthHAdMNBI08I3Od26dZYR2fEQ1sYz4PDc
x1H7NIieZbeVaOaYqprpKg64JonhiudBHOw5M5gO9EuLNIgFKrNnZWaFmBWQNSHW
5Mg336W34ESY84Uy1SuKAWsbAjoflOaEUP96sT2A7lqVdIBe2uw+AqxeIgEPVYFB
7/LGHbLLkMpbiZyOd6EfjdQQsbHaOyigc/s+Hyqjg9MUvEvrs0rqBlHimI1Utttf
gCydVwTHUJyrKxkS/ueY3SUo9CXG6r417W5R7hEOLUpLLRLOtwsjc635z3cz1EBl
vxMToudIbC+uhVsONfdQ4+Bi6cYD+lDixh1f3BjAN1bQEzm4IBXkPq3/tZfqkqjQ
IO9ka4jXzmup1okbzEl2s6rbYFu5y7SB9rI1xGZUcIKQsfTD2N+Rv6bZtwcK5U3i
wWTm637N+U1zv2DSRw2mr3aaF8fJzAYHOMR1dHw46suju5pb7bL1v8I/PqPhE3BW
rHzPMolA7ZztohEJsQ6syGG9TyOqo1MOzJPdmqSAK0s1HPtSbSbJAjFmVgZbqVc1
0Y4h2UUtKqabNqsleMpBHvpzCEVRv0m0DhMdeMKOawBdULhRDwxxs/aXHI8qMSbK
sreRaaY6+l5mc8L+DJNGoW9LbN4O621dIQXlrjBhAI3rHlYdxxorf0p4p95NN15n
T3cNxRYa4WHVh5qmMsXdltadKgyX4QapGwDuccyCY2a6mXCSC8a9f8SHhC7mfokK
bnCMnb/CYYnX3rzUR1LyY/Y0Kur0KVJ0F1U6q7ST46T9ZCqRoKzas2PYjuYoaIOB
DCtHFA0EhwkWKimavRxH0cLJRRAf7KrilVKCtacNeIJYbQcGfsQ3D9X93K6ZWHbh
2VIgwBl8tBkkH4aiVayZzuhbQOBG4ry2KEnTgEAYOTBjzWv0VN6koZsDIYyZyALz
MYXxuXTkd66RwM0100cqEcGTysjfKMQ70t6LIMGDCbGy71Z4+i6zx/Yjx19654gk
2w5BYSZb14cnY9upGI9jccCLeaMdHyg/v+zxr44jCexnmY2pyHLS+abdbgCJxsKu
Aiqm8FBsJHkRRTlBBi2MXU6DkuQmMFj3FmAEhCkPUKnhAMdd2fJRJaXxlRu6kRpX
dYtewlPilAxcvgO469EAE5PahcHQKoxmfiIX7vbMzSyw162SoudAdH2PU2xxJWL+
FEMAKWA+6+kdShuVTiWQTy5vfcPBp8rTQ3LCB4rKQSC0h398h/rWl0EWDRHUCRlA
7uniQXMJNpoFDoq2iO8WCbm9zfJmfGtg3hKdsxiRz9Th9NxN0CZ1ClLveSJK3IZC
FVqMqQXCzaCSE2p+4ybtOd32YtFAFneGIi24Tbo3N+qGJrEb8CVqaZIpDWzVo0Uh
5b2JGaaMsNzB1FLUuK16Spxymw6N3xdO5cfx+eys0iNkkR/B5xpAM7wYXjrNMPOp
ESDdIxSr4j6ghL4A2h6I4Ys5JZnYuxJLALAMYbxeHUUNWG7srCUwnsWR/puLNRzr
si/QvCHPVFeTe0pAUZsFYy1DdM96QUMfJBist1kj8qENksW6AuLZ0P+gNh199Aa4
XBtfvou05HnZaHTo6W+en/eSjQmqDQNZGj+F+UCzoBsNXhLCMpnoZaFpvyXL2hVB
PMzrYpgq51912x/tG+cs2HGEzLx2o9RDEOMfPHEG+KLm4rXw8wExo/pFW0t+xUdS
VC5gHJKEYBMrx3RPW2yPp65plJKscqqMvlBpYwEzwgGpiRMetJfhtW0uXImlxYU3
0BpJNUKo24UrY+wgp4vr0k0XF07+amgKyLpmcNUDWLXJa6X5fHtKLiU03dcELMvH
Zqf+rak4qmxvsbesYge4PHkFs/ISQWJ9cWImToVL0QU+ltJO0Xs39y8ggt5N/wYA
zUxvBsaYB6EGBLLPobmyb9i8Y3WsXKZL3oq9Jo1HGS1/w3YIyVGOSBSvPWrliW+5
5UiQpHzZWsVsm+dmm9zz21xRLXbPzk/LmIC8senFskAwJ66+ZB119qZ2QCcwaPvg
FdtxeeRWW3FrlxR81+IysQcTW9dpltQHGaiQP/oz4QbjIWseBWDcpWnw+jaxyEOV
NpA0NGHziqttc2UIcGyCs49f+xA8AbsJ5yiRIziiwIAW3UNaky7AgiTREMW6zI+M
If4Gx1m5Y+4jBe1SPMsemv0n/gpnVW+6i42yuRcmXihc/0Q4bWz7kipz6qi1scUG
zU3CJCT5XYySkeUjwBTnDqLXqyRDqBfDRLJCdxSUs7n69ZZ3TchHdnHN4zXEVwO2
jTWoXvw76TsTj0XN3AIAkogwfMO5ZiUxPc3UlMd+3kDMOgS6GklPrU2+dEDb6yiJ
KQze3257+SLz0iv01d4vwKrz4XuAB5d53/Lpncb3XeAfoOECJPDMjHAZDIwad0IZ
jv2UxVphKoXROrD/UgwwQSqy2YNNtpJYnJMdXaiUMJUlibDG82iYUZyAWGWE+zqv
zoTank7EfhqzyEIkC+vByHSG5cP3xJHu0LFs9RYlX5HEZlmEp+imOmaza6UoA4WC
f5dz9oHMmSc3n21Pq+Emwyej0lsvXyK2363YJ/2Qv6alWMQtu//qb9OlrIkqm6tM
yMb131op2LrMoFsZol3IlzI/oM3cwRNo31xfYCgOMheX6ILPZCWsGlFDshNWah74
wdquw0OfH9EqAwdggS8pVTDMz+d61NTp7jAnfhZDW3e1KnanNIC5Moq8A0yBWCGh
kEgHI93t7Ks8FMLFKZWnGvryu4E57MmA0/K9rX8EbX8lStoeTNMSIFGFq/xDP7cv
Gw445u1oy61YcicFAnietPMJLQPZvbL9Rsy7t0vmKnqcJLzwVSdqe5J+8gBUCDVK
l7JvYBUa6r5HNQTsRR4yhUju0xIan3jFZNyC9YFeWMD3qa3DZw1awlsMbsX2sW0+
lzzfXKOkCxO9ACoyJsSWlsFpMrA+rqGD/M1DdUU0q2vG8QDdeQgDDSK4YIENRR9f
P2mOB4Nnslf//boKpaWxejbjH5MvXt9OjmNjis/y42q3hXF9Yow6eVlgUJS8D6xV
mfCL/pr8nUKoppo2htODo4YUnpHAfX4hZ6g9mIyvRG/2o3PUpMKqRmiWddY/rJcU
hWgvGRLJEEmi+SyfVfWBz9b9o7ms1xIs/QeCchI5Pdyl5ztjR630oAUYK5/LlvCM
whpLmS0HrYCBl81n6JktFkQJ1dSLb7EZYuWPqatkqzoXrxt7nfx7os95Zwb5PB7G
bb7Ld8h3NgS61iLs1GL1mKffqg1F0r/UPbOBY2AVLS9/arfbx9nmHnrTw7vW+jVh
vg6DwWpAtFAvLEWK/Tt9tw8hSQSanS4esDXNcczUAP3AfMnnXvOjitkO3mJMV5qT
7lubnga6ej7JYu+bmZIjGkvpbhChCQj9FMFeIfeeSXRCm0PyGJ9EcEp+KSH2ljbO
FTx083HBePYor/cmYxS/YQKyiALVrBR3hEOc1IIZEv+Ps9FO9aOWhgrAUJKjFueC
TCkamHNlJwgAGEWoGRQs1+cybQhCuKiZg4gXNwCQZ5rw9vyxkB4vDW1jFpY+xMq2
IYTACUG/z2v3p9ep2fpRvJ1JTkJ2IUVff5kFRxl6K7te69L8XN/frN2kSXuOaBaV
1CmPyWZkRpSHMXbSGnB8paIHezTDjPsDuNmUQVkfFExt42TK2Zr2z2hO/HPMHhTY
aloW4QbI9teIkS1tbiBLeBGVneUou8SaijyuvoKJ4SgnDPmVV7NtFTrBIDLFmWky
JjCZNF3KRFKw7DHkNtmohDvNQGo7jB+bmBS2dipLsmPRYQL8a8ohp+OJgrpOfoiC
aWNft+WhiVUtJa2Ku7uYsOOpLwE/m2rGK4GKTkIk6ccM8/UmhXZf0P4S9j53jPV4
GkGS3IhErs1x5Q5EGCy9EHA4osD7FcTuYqbCzwV6WFr0yBOxneMiOYGTlOQjw+I1
6Q6dl0Gd/g82tSMmRYKccWWv/2HRBlK0s4mcvZxYqOYWSDfM0CkHUvul6tZ7gxD2
e5mzluXuojPU2KrmO+vAJXpOOCpAHb3N9uTUCY4ViHTnNP1c1ZGEsJZsvkJ72wg1
2JrcxjOt6/nundZTbaSbQopaqHPLXGytpM/oFaKVM+HiTxmtahwxnJHc5XHmOmuL
irPONN7fz+5/p4OY953RShLqy3H7aSr19sEgBFkH1FyOhge+1xf3Wuv72UXcG1ja
oCeVATZWkdu5seBKH1AxyKX2SUd5Qg6AgiM5+Zc+H5yRVGV/8nkv+bzvOocEiNde
FOTEP+DatfTykTmAdEImY8XJBr9Md1+YD30h2YF7SicWkrmLuhHZCsT8hkMdLVcM
dnAe/yXJE/MMAvNclABPsrDjKRHR5aipZMEXfAlmmE0OLqHGgvcGhRHeL7AWuuCG
Fwbtc9Tk7p7IwUvoMEC/s5Tt8A6iDVAjKIV9k2mLLq6hcgZ8hS8PrP4QR26l62Gk
7eL14W5fEvfrRFNxTAmULx7OiKEaKopeJBDuma6GEVKy/jvz+nv+m7JHoNNDpXDL
MwGizzeShdMg2ALbEPWKFzg9cCrzOenIjDnDHzwEmLJiksi5hcXmEWZprkoBCe/m
RmPMAhHNxRxiF+uUxLfBg1mm8EspKJYVrWDC4yDF8MUN4NyKd3nxTjVYp1zD0j36
QP66bv8YFNpBUNiZ9Op+iEtVGHUfyQ+aXj8xr/WYU5Jhr3TV2EIcVQrnDsxpsNFn
O/FlDhRWZdkec3otsq3XCpt6yoMnwvoadibPNue+vysCKORW/oUja1pHf5FL0Q+v
oGdQ1m7LWLB21cadb6VmuYpoW3iIrdtNeScVfVwxX4s1ao8TBZja47MJYzNMdtYa
6TMhla3ia3C2qAVvpBNRWqxHFqOLuvsFrp4k6Sv2Bng3fjel6UTyzV/0BwaEDXew
HUlMslaY/J0G8V/xAm42l+MwR2/q3DDnIp6cxxlKYlVM2deYT5L48DQhQ964QlH2
p5ZtIM+htKis+nPQAM7LEaZ2ZeWAw9FH03lAZLuM+Mg2eobEum0/xD+mtDbegwar
sdXDadD7g7LaO+xsMCpQbS9qvbXcudlqHTd94OHV854waztatFh2DXfBM6N7Ij0a
i2HOjtBHbhU+ccdSiA7q4sjvKcWt3WcsvgEuKOr5cEMP9xzK6jtwqF5Fdxgc2ATw
cqrw1op7ztOx5SxXXnp9Op0Bv7g0q0kfTZGaVmmc6upMk89Z1pPnfKW2Kra4Oio0
ee2/roLk6RZKy7AO7jQcZzA2RI1FCNxGWNEQ389aup1wMIlTFkHIlWHh5Xl3o41l
BkQRHHgWLDj87b04fDYAlcErnfDvBvABlXrOhIvuCm2TeedKuqKvenSJB+MtrqJa
6rDRthmX7VQmlbrMUiWksJQCzJIqS13i3rqDovRKuyI6Wf0JyDA1q5nXIe3ZgRxL
Ya6GdVRlVbdyP/O1+ABLFNwGJ85Nh/0dXVNNZ5Q36upslnm+K+vHDLyI242ZlFss
ezNlT0WxpkjMCcnTl92juIyU+DiPON+ENL7SBVAFenirflyihyZgyebmW47aFSam
kdRFqm9KsOQX4Nji4RL8Xv6iyCBpy0ZTx5OM55jjLfm4ul7Dldoxkhi3zkggifAR
OOp6UwZ1wpbnSsCgxJTu17kB11dxSLI9AWlmeDgjk1F2S1xiwgYG+Q37hVsHv7Y3
yT1sf1ikwWdfCD3lZD/lNHLL8Is0tMKc/MgeJE0nHc7w338GTnAFZu6VDNjGiwj7
z2CDatrt9//kZ5UT7mkLk0H9naN7fit/gfqoK1EuZ+P+U5+zdXFMOHKm5t9Ulx7T
2iavGfw5IVbKZMECdTCMJZxYXmJFANEa71/ojMsV9X6mTHsGTBZ+qrfYDQCL6FSO
nHb+NVIMS1X5Ze2Pm2GVGsePyUOp1XcJndF7KxGRuJbAs+QpT5CvZgSAmeEwruXw
pJ178nK8vIzNm/CiJLvw8K7wTFpXdQM4+0NaxdhgueLVl/TqMkwbZ/LWu4Vby5aY
XDwUD/3BcLp/sgo8AJsj6Vkmw+ucCKQ4Uj4f0K7VkPLg/xPTovIHi83gimlNCX3e
TvP76kTJVAxaU4WqeaMZktL/GYCqEJwcXXslqWQrHZjoQR045YhKffUOPTZdqTVw
UDf0O59efEv06P0mgBWx9tUd9Kei7sV6bOiwviAAEF87EolvwWvnb2/QdZxTO+d0
eE7tLIN1nOI25ymKXeDzpqIcY9iH4Wrk6UW6orC/wo+uV2yzhKolYsr1zhnz0x7F
Xc0vaQufY6oNFQSp9bS0+nH1nLu9RQT5BVfIxfirN1MN6jHuFplA2zWJD4YkhN7t
aJbL+0ZbNoVQCOHlxVZ5Am+fy1+jZccaZwtjVeil/SRbfV/rLjuqNg3ydCG0e22Q
8ziJ2oEFQVxoygX24gBGiYMHjwaUHWWmO18MbeX81KS1E4r2OxWamZKNl3QoxkrA
EIDf6FaZiIaF6V0ly1QJu0eHdg9X351m1FRONFpCWTBImYf1q+Ju5pDEJWk/Kexl
JQQ94uMbKawV8tjEqVWzKhqwls7I6lmEf9gBV8UFAT+n6mj2js8p3RSqHZNJflAp
lwPEgR9qZZNPWecpNOTncb+89n9ul52LM+JhSDVvs+0kZoqGF6VqGdr+A6RLzMUE
yDoeNClFLhVcvjwBOTHObkh8dlyJfr3EGZZ6i5ROgbwYc8J4vlPsv5rnTrhI6xku
iWp6zIwVbtzqElXIBSIt3nCjF5aIZmnewG3Nk6MkTbUp3l2NyAOmDwFmfcAX6URO
2XFVW3nQDmof6oqo7VlgTqYgNJUabWGPZSwJIMDVyVVAPa9TuMJYBMOIiQujHLXp
JfwYagfl3ElOFse0bQBZ6jAso/sHH2uJx/jdFLR26hElBCTtab2tHr0V8NGSmvLi
GoEfMfzvIDnPKnzp8TmtHZsBZi7yJSkpcydDMDg636HkKdjdqgStpnf7hPpcYlt8
90wCxljfOis8cGslijVHZWHmKiUXb7wKckWudGXs+8MVJ2yK+JOBtMixnxiclcew
vY580mLBNMz1I8U1lI2bFXcshGOlBopgfCCnFAmXnDxrXY7hrS8XaFnRRKe4PAPO
DttLmAZ10yVze6bSe/NW8N+9c6PLw8XkibcU4cUsCBWGQ1t9SRsuZ+T7UTtLZg3F
tBRqQWPgoaU7pqNinhvR7q4ff2aPKrfxIdmsIPYq69eAnp1KvlTPYN/TbM8vauPe
y0NJGTRbARKVqT8kYE40OuexsOCqdyXAArQiX77ydLtwpLuqYu70ac4QTrMgxO2U
8F0WxhhEJHrrDIyQuxlfbmGFwQShOzUtEXstxeHkhTjHN0IBwTpGm5hpvhN+b6VB
hqDktB/4yJwF1bfD5U8yr7ALCzajP15dMf9AolviwyZQvauMhsp8OleEKEM8VZNQ
MekEi2Vsw0hWWHZ0Fh177iEwfCOel/DGKsSOeszap/tCOMu6JZs9hMi/sjX/Sd7i
eXQttZ14hMJnEVJj1bizl5L2vrSbmjT1ESz2rxslhPc5aA0/BsU3Ge00bdQ8dvJZ
pkBLGAB/kTviuo32oUsiPZCq782x+hXDkgokY6RomS74C8GjCBSyVm0WZeMNSX7g
6+GbZdoWie8JXiQKXFSl6qzMU4qQbzT7cYVgfBY8BHvTADmu00z5Px1TRydjWYY2
9aMaA+K0qz/5tzmk06QffbCvRjlACoNOjrKQyEd6nrW45H9WB4bSdwxQqvCPq+QK
6/FLr5TWWj1nzet+9XU2rmMSjaTlci8I1liM9XZ5ggUcsp+NTVnmfOKWiIOU0RQg
aLOXoSKd5OkVqtt/j82HsRsqjnWa/+pvwyv61zLS/QgklwXyTU/r0DkhcCzPxHHm
I5ZTDT3X2o/1rx4NWH4SAkYPS88VzmfaG0gjD5oTpGENnIxHQ+Rkv5MNmnO0V7Rg
ut1g5GW/G7ptO2WxzZXmwY/ASc/DsdJDQszQhd9DwiNXoNIQ7VzD/w+w9qZCJSXX
TOwAFV03j+aFlxklrC5uvBDfjFXZTM3l9CWHjf6H9LPmELUJ6MSY7AIyZHIUCtSC
mSPdq248mVHvMFys8ilmtzEbZwQ8M3PWHWoizmWmigdjOsp0ccssiEN9umcJlnBk
GAbXZB8iMAgBhwW5ivD3BUiEcRv8dUGss7YiIgrEfBo3F4V0uHWjmzmLUuEG/Fpz
L2wEPcG1v0gz6fTS7fVI6JUKl8a8WK1oNFdYmTtL8b0UfUQziNbigXZEOHFU7Is1
PJE6/OZ8jtSloXziDUiXI2aT6FHgMjXfCMKvCPFMFsysMuJc/WcwiA1jmqTs4KT8
ZcsK4NlZ1unNprsW+BcVUHbv7VOc5Z7EVVMTy9Sw8BL5jyVMUwZl/tpYpyuTEzDy
hPM1KLlKB3/3qXfaHtZi80Uk/atEqzBoX2FfmxE13XTekPy+ZlfXbbUKYRn34Wfs
s7hHbpaSAn8JaJzFO6+XodKj9BXRuVAYXEtkhjoSkw1bZQbXQNHV0YhAwedI7VK2
5M6cYTJ7M3nitR/896E07XW/usnasUt5sATr6FCP3Q4D7QFSJ1WQVhss9ymBmEew
+R0x/Bl1FFBZlyK/O/870Ewjr6ECGeTIylFd/t8ojy1phNlSPHcFXWqtQxgeGdBO
tpV1nTnF8wNRY9A5F7SXEaCW6eHF9TAOJV/sa7FwYynAKqmpnqmeaKNO9Mrlm8zX
GcWLlXFP1JjCfGX9OkLDtrwSWrCKHPGY+KPho872kdJ+FDBj7dhhLrFYpXBAe6OJ
J6OXtliX4JnemauD7zh+w0LeJhxIbsNTrmZkswjNyirDfTpjX/1G9Ty07dbE4+uf
+5JT62TDELm/ACtT6kjP4A9ZTT6X7EN7zlZLyggX6AAxWMt+HsFbz6WQJ8qYmns6
rf2tHENmV4ZWSZKA2Uv6aJ4fUz1MERKVAXXhcBLUcw5lmhJk78OHsixLTyJy+F9u
prisdqsYyV7yJmvnFYPDXIMxAF9XESY1Nofgbm1nBusVKjYb3d2YReIuI1xu+4R0
k9JxcEE8KiULjd6nRL1OrFs1Y7AvdCDYrs/MZtDx4YaB4z499AJoMx7T1zS4BQ6O
RNDaK0XktfBnG4tQAPXDIL2s2CPVNRt8Mr6b3rPkigTETjgbkgI9W6SFOnP1yZNi
23mJZQkGq3DFDzdDcTT2IC+2qMYUnOwwwFCOO6cjXAq3bcmI4za2f9zX3UGidMIc
TYPrnuBfmgndBeTSsMaiheFgF9v6OqhW3bcB2l/r2U5eumOYUNbDYhwqhQUlG5+r
cdBjt5RYoONq7OpTo0OqqvbSLY6v+aLz5QRp4Zd8qzhvKHPMy/Zki77kQHMXeV7U
SHZZhjKzsJqNJ/BV1Zg9piRisJYbU7yA6Y1oeMsqLjSz7+U/rDatJ8IlKEXZE1Fv
d7rlt0UWNULfmBCruWTZMBUFxOxPMn954xjyqM62SH4qe9HoFBr1ofzonLlLEmWf
9DjGQ8wZU67qyxNot65WiOUwd6ktziBGbxGXWgXrSPXXXeMRaZUGFOdbFsBfnfNh
vBr07wxo5VwK4ViuVjE2At4SYMTRRPdPyGiMySqhDJj8ON2BPZcstoo+NHMQIosK
ChTCkj4qa/m2qy83ZvQ3zzxqm0IFX5DVinEKswEOPCM4nixzOt6tSX2Dts8xgA2Z
c5IFmIziDQsq07CS9H3RJHQUArioE6uRf369vUg1+4Z9vUS38ItbfhWLCF1Gdm2U
wbEw75E+/WuSle6v4zPZ+KUTdr9Pcm2b+mFQDsNoqgPu+duxIrAJfkGeYN0OQHYx
mpNMTpIK8+ynkiy9iKJiWJI+ECitQwiYpO+oOttPvFLeA/zPNwhsjlAWw7DBL6DK
Ea5owP4IznsutgflCcz9Dbx19wupNNLXGFJY/AobWN9SD82OvnbGsifNZtrJtQyn
Xx87aqmGu0BX2qFjG/4jactQelOQSmxRq4RoLkBU3KcE/k18nwxtKwEwdsmnjPEQ
awArEmGuM/0l01boy2rHIbtjnuA3xTd9rZjKuuGkQHVrsVsCrvYCY8Fx+7CJ+10V
HedEIEAXkVi2IDxbN8bQTkdDu+0MrkhDBXDD6CcIzWySdq3DFOTLmpUlVpi6uXIP
3c4IBCPVCQ8YDp/W3DHHuLWNNcGUZopBHlfVS47pndL0D25azkml9LWk+dakQXME
+4mHgxd+nlNgwTvSShpjgdL4MQTPdRfxlKGtX0zQ1RDq0RJsePUjXrrXkT7UeS2N
SMNPL5iBucbXBbbP5tv/O2jF2rt/3wvVXs65kijo33YSQH0/cd3T9WE7FPzPUnnO
KiMktnj1hsRbXDyIZ0noUtMCrDPJBhbgjfZAkkCnTg9krvWkfvl/s8o6Xmd0ucnS
o/JDHH3dfGawUye4/IaBVCo1glDdj7IbcaJNH4xhCbRti4/ICgm1SZscB4KW15E/
7OiNcCWEd0QqLpiSA5blwb966tHdmHhEc2PmeRV/KcEzcmNr2y4sRAcog0UTdzUp
XCqhutIJzmtwyW2vcIZ+kiLNFLUh9VtLhtdGoRvNOhTaPjxAJoLDL6ni7ZOLsR0b
jYaL+FodgRMO1stSOzROQafrL9E65Ws1CxGfgaF0wDDR4pPXqqwAzsIqQQywWjxH
EymK2fBKhIavZKRzTGjr30MXrOTt0FtZIKadZApacQJDFyLWcE16Z7Us1CAlObAc
HIDAvGvJIjwLLiwEPFUFEncKjw0PK2syXI89KR+B2XBN211e7JRCbY78T0MBTwEd
GH+7I+1nhgQ/K9fwX0XKxADW/++EyI+3EbpZWS9f7zIdqFX1y6A+G20R2ajFrBVJ
c2mcBYKG/hy84MnOsTxMdCSDoQNeCWel76DZIZWLjUwXndOFLyDtZHDo4b35SmNI
99sUj+tDo+ECvXvPwPOGpzWLtantKjaPj/xUPy5ayZgD21vENz7uWSwUgSBfjLAD
gzAhsMSY7fCtQElICtRLsGDEpc9DcEO66tP2lKtncKB3kRMprH7rPwBG7PLqEoJg
wStMUEH/y+WNJu+/vmVH27G2MvNNqbO83ehmt63/m2ZjZcB1SlMPC9yEL8CisqvF
2CkbGL2PdH2bsWjNFButD5OHonMsCjJ5eCSYE/qBue9HHJD+ga8k1bStByz9DowF
pTMPLvRsVOs116AYIUQsvoRXkKBWxD5mVLwRvRQPaUekxbCAuGd9IrEs3Pvhjnik
zvAg7r5yWGpwa4hq6/Qo2/Pb42uFJjuBS0jvbqqQ8SbdMI/hM7I35/l8m2e8Xsjd
9ly/y6y+mqmdE9v39eo1DzuVjZ9r0WLXByAGWdWjlZku6HUJK+hF3JiWCUPSn7E4
uiynl86GxGwWJlUunUFIwjPpZ1Erw4eEjzHqyhDdZOqA+R7kee+/PJGKrII8kRZc
/4nDijdX0psymR9loi6XBnU5osh0KGhcz5xdhok//fSzWTBhxDSeIl+RzBr84vrX
1v+4L5yIvnPDaVssnklIittpmjOCYZc5MV3oJAAWGyultZsTvgVc3proLxvil3sY
xU/NgkZAebeazAUOxL/L6Tlt6pbFyglTjYfNmzEfPfhy8A03GixgA2RHgw4Ggx9W
m8wM2K02Qxpnvy5CH8vSMdDixwR87sXvepmQPj/rPo7qQxY+dO3SLAnKfQDVr/At
Odqu4amGuk4kbeqOkVX4gUcnP6YccuxJR0jZAe0F9guWV8NUaCy8/SAi96W1rMCj
pqaTXKB9HUa9hxSgScfnKMTqVQOYacJ0uJ35O7jDPYQOhWteFMLqtnrB5WwMFvOe
dvpvl9vXrppET2dnbzStY1hdLK0lgqzvayUF1eZUfqdYblDiF7fEnr9UaXnzY1+x
W8uRyp5vfVN0a0o3roTQT+bnq9fuRO0bROh5Jk/KCMmX5PDDpE+IP3gHTydc7LXP
vzlEOfvq6mReqzrprUActv5qvuaAFmx4l0sNPbUwyRvPjBont0Y7tbB75wzidv++
jMFd4b76GdhEkGZYdqK+q1+tDrWhDVo6TGUN4rLHr4ZaZS9aJL2TFggzWFe0gnVm
97QLFrbi2UJmPSDKE2V0JiqwnBJ7cOqxAE83GGNxz9Kp60RT6sgP78Dmv9jqIscS
YHRyGu3+noUf+Vzx4S5VlFi+wOmddgfR8qk+LL8NTTbRSqfekRaKXRYmE3Qe6c2T
jcCNjaGYxcopAdWLYBkpL64fh1TLC0sIzMSr3F673ndIAZnymm7EHbiF202d5sNQ
VgRuxjSly2MRCHvIofdwt3cJ4Z1nZApfoqyCH/GpmRHHm0U9Kw85ldAEVEe5Xz5C
63ndl8JMOsayrRLFr+K2kvunPv/PEXHmQSAM47QX4k8iO7uFbKTQb22onua2vrkP
vlm+58PDeGXkaMiyu2TmZJjDC1GUZnvt6FFFe0JBGBLrARGlTd0lMd/jMViyCMlM
1xKZFleZRnoj9xY94Lv2ohV5mE8F4KAO6/TYcBAEXdd+Kt6Z//yudqDLdR1nqRyH
b93EVoGQ5btc94hpWaPuBmNt8o/EJ8mOKqC7/SYjX7MmP809Wm8ouZ9/kinXYcus
c7ITo26Yc2g+I4z4WVJGkqQVR7adRwSemmWdmRMYmCxGKnk/rurbe/xvJQ9hjSII
LRD+p58QWEQPOdVTc5kV+CcwKdwvHXeloENTFiFdwatPuqcpqXK67u6N1HgSvmXl
8q6FSSAywGULpxxKQJRIx67WyBHC83k+AGgH6Qk/MDPJLhfj6LcFiDZLauZCmP9B
CAT3zjfCexWDTQtfAIZSBfDOKN/14QODF30Sxv23Q5qpVehj6PMAZCsRDn4vnPnB
Ic0ZgXbrdAGLinSon/FGUXNDeMI7njyI6uvQd2w7nUmTvIgKMZKBJ8hlhFlxQePf
CpiZMlv6WLlWDAXsUC3Qd6MmGd684qcUiLwRVvQWf22MuG2voMNrqnCh9emxcmwN
X1yRKI/z6PhxwkxUh8TByFvHKxVxH5DO4WPInEv8uplM1BvwhLq77Y8PAlwPZ/nS
agmTcBhzI7M7Mo/MX/STCRshHKXrwCgMQ5FAXeiqzjpMZuFBLYMCu1Tl0kPOVd1n
LDASBXmRpJADZybCvWdxj62wjp/fxEQUURI6nxxTZ5GBNKhwwvv18EW0cGQbac1E
wkZp3oxneCsizEsGVU/FIzR3962WJmXBS9n3b+dy7nKNO3nMgHgMMHS2HyKwS5DY
b8NUjufsRMhW2SxEluMgCTyygNQ0TIfLPdMilMCQyqQmnPJmMnt14zQ2OuQuQKt/
WmetqYB7fpQaaN/v4I8PyI/BtZMvorsd+SKKyc3ohGIaXTJ9Yxd4AvUOzAep9Jmf
kY8FB0rh9g1y4PW59Fv7Faa8YnPaz5hDec+vi5OG5N0u4oZdIeEUBBeOxehRyK2q
VGmsCdddUmAQ02ZOqrchj2vh37xxATRDosIVd4ltBX25wClEl+tbPvF0RASq2cAB
PIq7iC5SHLP54/Gjo7OC0aCpcAYYSGVHjh8CsMC6/Bg+6Z3R3cGroGapc3rDWtsd
QuPHPV28JKPhp5e3K/ZVza45AGzxSVtY9iwHarusupV18194ECmLQwrN0kf+K8lQ
WusU48duJTaNx5wUH0imBqPk/rhxMgs5996VOugwCutWJ7kkSTPlRD1NUwtt4/Nd
/Ax0JhxK0JYlLyT/NsHxfUaReukFnFE0MGI7fs5Wh4fg4BfUq4MnMT+HTUPGm/ek
LjBeSJEI12AIp7sMQp3tMz7wQOqeJEOHxp1xgnFy9hjU3pN+t96I06Mpkwc+yztM
HNum4Vl+u1vXf8BK/z6znaHgLakPyhB/0111p/dWGk8cy8z4kiKMDRlk8LEG8zYV
CtMqgJE/N3uQ2vpCokIjDScwWsmSfYhBjTbP/Duv9ALua3XQa26F0ksKs3MEFki7
704C5EMpWnzZmTzwfhwE6RLUYegjitBfS98ldSkGh85pPdWCj2Lv62ZbZD1mcENP
LFoq6A0y/hMnPrO9BY9i9IPAipJNf5GBIuFiId3PxzfldJEu6g1VgfslXX3aWYyz
LaKnojyRphxlD2c7WrPWlKUZlrewLgkRwhiI/oEqGa2KFvbruACmQjZf07DYhrvK
mzPVT+PVJ+QaLXzv/kIODQwna14qYzIbC5K5fP9y18xEmGDsqJ0+BvzWfCtr28oB
9xJs+RVvVcturEU1eTw63LeFrwIa/872ziu4C++dY9kY0Pr/+F8emvYw35SBREoZ
QivKItNfOWcIVbbqzFcpfZ089zqOapzt/+h4VV4xMsv72XgmUekPNE1pSOsd5bRn
niGKeK/cFTQH17S0m5i7XzWsMIAUKfMK6MJCfjromHf/4Bji4mx7ST+/7TgbeO7M
bvx7dk4kR6C4itWOzujjsfx9ude7wh5xPGBAkaxKgCGq58jSah2G0TxzImAdnO4g
LWqymUdU4b2FY8zXMfLQrmTxwyGfcPrnEuNXo2DjpnRq7g8r1tUnh0hrFcQHeqGc
aBQ/fAglTiwARSECv5Dunstq2GkWCDs+zzSotUiW6HNJGjXvtO5K0RMJRqsZ3FDp
Mdf17oNioVFb4aRWoi61vFQrmWFVA+IleM9zwtgLnZ2atBGiPkbozNwjwvSZ7f7c
iEzWUm6u6HXNNzIayX3TTq/LF1UQSmjD1zbQl4dlccULz/RBWTfp5feP9N2Mw4eo
pxBAylT/TZs7L5AmgEZqMouSp6wiQsL+AnAUo4VbzFabs8oZhiKnHxxk+nn0crGq
u005dyGCqBas53L4ZvO81y86RATkM0KfZ47jKvra1kuTm502vaWOWvlPigcnyjAS
pqR3LAbGONAE06eXwBMtgBtlYWeoFafzJBBL+yG+SSsOhA6cnu9Bcg9KhPZa+ZEk
0mvYMgZqltHYP13mMFAgNXcZV7L82Bn2WqECuRr0VFCrKOGFzYRj6fpuDjjnUh1b
cRnwRMxug2ZMurhYL1KIj43z9h2PDgkIjm99jlosLs/EhznSZcr4PLql/MRjLycV
4Ft85drsLHNlH7ASs/gzhJ+baYrg3O5I4k65uYAiymAlGMpIxy7+l0stcv9/LJzA
k6bSHF9f3QL7ZN5P/hWniQFqm0SonFrnzRF70x4ljPpHD2krdCIOg4vPCMwVS89X
+92vb56l99cDnwDBMWTgPkpCObjklJieruQWnuxtvLmjL/6J7ceivoJoKd5jBlYj
5CsF5x0hEmZz2ZE+siVKIlqZm8toA35JlwoIt7iWjXuACmR4iEHntjmWxObQ0v4n
oVeLOAj1+/sQs80zC2VebFZMvXsJ8uxxoy1hIVxpmOG/F6O+wtt/WMwWF0Dj+trq
xtjy7TfLTtWtiE4UI+5G/9Pq6257VmdbdxF7+H7R8rfdpwp6HqpBBC3qwM28Ow64
ejjsAkcHcjVdhxbnR6T71c1jZ/tZNo+vN1KL2AHnPac4K+q+BYYdK215gMCbR3D+
LzPjCG8aXYclCJ5HXeV4z8UuD0W8RX5FhT/rRki7SuNBpw7fDo6868OOx2SPwkj1
ryJacUoNTjBYMbvLA/qynZGrhm8aSSt2AfEkNOtqwxBso4V0Nl7oYLSwWu1xTZuD
giDz2k3WmoDF+qUl8nmaeFm+mU+TZT/sljYcKf5REluDcENTBnvhH7s5O5oIdxV2
IZkKYXtYur7pJkOSmyXOT5FBVrQqSeIvUPrXp1aEEAw9mrHGXqrrnMzsnIj7S5VV
fIYM4oUte/+5sc3v7mMe4EsNBWA5SD+YCw98dIdg4jrXxdZvir0ohAurDbrwaOM5
5s9aPSezr4zj++PZyeWT4kEWohb1K/dGqYth3EQUshhheIUyB8cDnY1Eq37q3mi7
LBp+ocMHHWJTigFtssypcD5se2Fda0NeXm8EZz204XGJFen/ILGKgsx2EBm+Jyxt
I6wd2TCtuO/VrlVUvc3jb05s9aCUyfrMPuaqE/g16JvRohFkoMZH5KJn5hpfySd5
lEuFadLtGuDN7//GzP9ao5LK2qYcWePSJhv/9+HVKFki62p2D9c472Tj9Yy62zJV
faxXfYKmp9i7bHIn6FXkcgSN7L6H9TAb5TmSEe04etPlJKTWkUh0pb5hnK/QIC8g
WwlNE7sS2PuhAl8F+04ErPtW478TWRmk1dbcvLxnvhZj4kliSZvV9VfjghGr89fR
Rp//EP6rW6OP2cKS12oaC+y54EpvuDLkN7XYXf7rOxZ7JdDezewzkfi77o61iO8L
5247qal8CGln00FXrdtp9BDtiQUaDU6xFaUO1g9kLkHnf9Bv1MxsabQrWNklpLap
CcoEogDjlyVh0D3iOLQTnt3qvnE6iAuVf92SI391RyAq54273kz5UJwwVBXhPPGI
M8dMHWynm9KJEVxBOScEUMsWNWX+e2y3ohMLrDPSdHj1ICWxb6p1mwP4axr45X+l
lZlQmAIo4WYnRpp+Aw6ts73Neulb97THzcaTHE7fUeUxqP1XntXElR2FxxG0SY3i
3hN6z0CUf9ILjvrfWw4S9jvBLv4L9CE6Qtbg0kCG2aStCHnxsYXQzQgrcTfxH3zE
tJX6mvE4bfxPFM3wF3+oJsy/2c9x2CuGd4zGA75vpVtg3phAPKTrfyumA87fyK3A
V8JwAPYWYkXuqOj+OHzhuSMuZrtZC5vPsgTYA2t4o5lVE0CtlOej33xS3rg9fe7O
ijUJyLbDW5FB7/qSG1gv91N5PakHG9VOYUVkqck4MPDJEnxRnxz6+/3HHs3/+ntb
bGg6OFjaFuT1yNEyPepM0A4j3aP7toaLIYhUXGASEpr3LkshukpZ8G3xooRAun9F
1QTm49OR5egI+LgbYQ4Av5vDiuPmoxReKzV39+Gx+YvtbH2a/3xJ8OoUOFkN1UMI
RNIW0YGcC0x5Fx4WxOHfqIELebe5yr0OTMv5hSUk759kDFZdUy4JE3/gRPBU2Eb4
Fysf67NkNjCmI9hEGO8VvWxpf6I+7ShmDyo4fv2uQeQlHyFtAvhpUXtkQZaKSntn
Zxd6D3dd8Pmu96sniklNKttw81m1AFjB9eSJbb31HXoQo1lm3Wqm5csb99QzDMUo
q3DCJEoc4xH8TFqhc8+60HK6DFgThlMAZBbZRdCy/7Ih5I2smC+sAYDcsZqOTWgy
W4PPmw/nevgD5+JqYKKI1M4DrAhE8P6KaheRjJajKQ1gabmueelwPDExtDHNXc4O
M+JUCZ51iaIiCGF5whX9Lq0HM52rFyvwvENA9am+ED6U6WsinTpv77NX1PBgYEDv
6bJXvWunYAjSjIeqxiESWKDzaJ436h8aedoaQsST4QNCqr9LbJ8wAoX4BDku6YFI
pqT80R4BOUt9zpjumSPR9pnsCZ3miuayARH1f7By4Wef/GMkVu+MtDdBhXViyk/d
phsqfZA7AYFIWEF2r5M9adQXLyrHuaqJZ4gcjz40RHe1I/1cwkcmCLua8A2qyxi4
VQHRF4C3yUsOVwnNF6dehAZP06AF8kkIXDnp1DgleiBqKDPQsVENpEQQSM3gBC3t
HrvHiWsgJxE2/UYellVnATPZYphyyQs2G8P/7ZVxlXlZg4ea7mDYD0qIYPJxT1GS
Q1yypXjfPn63hnzjK7Q68/4wPU6isdehi8VC7KgRkhgBGLNGBO2SyZyQDwujihv3
VkN0yPfGUO0KxkenSGS+ftg+JAQNrpD9M/8sxy37Wfv+Ow3awsCzDhsIAQVpUV4i
fyfr6IdntPOzy++ftEWbq6IRE5n4OV2t+Mnt5oaNBBHisD6/uk2BZ/835Cix0K22
9PqpefJg1gWpuYqm5TxnIfhw5yaSR17M9iWCVnH29her+tKj0zyLonguCCBDu/QO
G46J+jjfGGzdRT2POP7NbMYEyM077lY4FQUGE3YX6EOMHIVUq1lb6VYjE6Wvn/sd
Jb9Ms9Y5WL1uE9/DGWwA6xw64S8zvYuVPM3BIpCNC+im5hcRxDuCQMx+ct55sliM
9p16uZDwkae6qv741Zm7lKQHHmHIIMxSOBTWZQw6k/zDV4sntqbvtzbtkAazs3px
l0dztgBSI0E4eOej79S0GbZoBVEqDX0rVLuBwisJRQrLH0ApPYbcKyJf4kQIl/1l
FVtp1zsG0efyvaZH44Ma0toSdlziCKS9RHbYMHUnzrR1+GAxKVVnoGMZNqpFq2CH
e78Kppdp63duBSsu3sAm2P7ECgkabLBZI2w246n1T/YC/yRqvmft8elJPyU7R/EJ
NdgMxBlKF5Z6UL413S3Kv+Kcjsv185g9kxuka/pDKBtvw9o6GzCcK29R9s4ExkbX
Zd3PH19HGQfhmpbKQeEm6uMCUUq4cLyxZHvDdtnCf1dK9UXohask4BzkLcN9fQuI
5Lpasvbql5p3SS1tjNn5Cw9sxrX8nz24sf6H3TgVOHwZ0wAM0QlVY/vJLIjBJaZt
c45NLRFpuukHdxMXAl4d8/rV/5uZYVZX7w5Xi5/Qk1AeIyJ2+f3mbiODr83t/VCv
TSmXxPt46s3/Nzb3ZAb4E8bOOMlTvr8nEobiCWInYANOU5lE0NGkW4+v0kLcj36a
WF6yQqZ5YHSB7pItpm1xWkHjjMykOBeZbqh2Z/p3PJkZUfxb87qXdmF6XpSz98lW
zG76eBWR8nHY4ocEn8O+yBKAdtgiiaWk4eItozqdv2ADO+A+g9Axql02RHpPUjo0
69sajWwt/HroxsjGT/anzNKHNc3QVh6iM0Qm7dhxceieB3pBkg9l2woLwm9VcQH/
qieZ2SXAXYJErzXcsYIDn/xSrMILEuwJf4URvI85znS/VbXkzUx3yd9F58i9P0yH
k1pmbz61LeILxps23d0pFmjbXDn2Bcyx/VAEp07DHaBMgMCEm12Fpy/Yy7BWF2cy
XPn8agaTYc/AhRAS48uLehxaIKtwQof2MuoQIGDtFiyH3ZHI6pzrUr2GVfI2w7ev
SzsFT52JIrjaGYCVAH4CwdZlNhtIJFE3XgTOZM/GdgVAwtrbzeE/RHd4ob4kT37+
gELVdm/jUC3E+Y6C+DYTcnSJ/BpEfcDtbl5DpEQsOTsLo2BmFTbdlzb/fbmKvpvu
SkgGz1ZEBGBavA7lqYl8rrOVPJ1FA/bi59YpQcoYPqwqehfTa01ilX/BqwcCR74X
PkiGal+vaChvPgN8N4/9dOnx4AFQaCWD32a5bMWTo9OvDhXhjIDXgrxJj1Rz0Ql/
E/v7ZXjYEyVx0RoNBS7xvGC60sRhXklRspxvLX6S73W6ibetGSyO47BA2cN/Qti5
iv/yYCeM5MIPygDe3K0hS229PSm4IbwACJk4wDxeOaPGuaKE3d0HCfnlkdGqKXVY
o1yH0xPyYOFLIriPiA6t13/zpNz1/wVc5IWhbMQU/g44XoZktQ+EV2A+AzMQkl1d
E+nL0eDb25LWlxgytOMsh/K6Fj3N/TD4Vqeo92NSS8fpZZLG3j/u526WdNClqx/V
rbcK5jKUkyRibF5O4jYbFpskwMXUhnxlp/WoZIae2tKw7PidrYzvwFMnaCYFitdj
V4kADVlwLutZjjoBq73XO27zlzJM4wkMoyr48J2fC+LTbnKhIlsy50MM2P8GZmDg
7hpHX0mKD6vtvwF1Cl1eaEdepMiQLkGLTiKPz/ifcq+FPBiEZBDQ9P/mmDiPSe8+
W/9nkr6P8v7frCH9TLIAcUGS3iQt643BEz7OGD86SGOFH7krN8rz9W3tv1vEWcqT
F+QQY7ZT4PUOW5rTzPVq94YWudBQHbzahfEHwy/XQfOGzLjH2wb588c+NXSWjJeD
/Zv1QqIaX5Sq+WbMsOUzJKNbjvEj7E/yUo1CHaEl8XfC8ff1rmyfGqlOkYtqCqUW
9HcovMKmATbjohOJG3ap+LMhV5iK1NfKJY5Or7REPoB0hsv5hgs6cNqrLLfg5PG2
NFo7qdgXD+iuztzWCJrku3WjSipNhcPiusgnzzYVR7jBjHeOkKtFflg+vvSu8rZA
rF9vrdDKcUheIp8Jyod87tETMikRBmkUF4C8KJbQSdcbkjehjWTNqQU6wLMopv4T
4pOXEwksEoYDcoI0J1T9UJ6Kzs49w5pksBZHf16olNIK4tUlNzhRvD+lMTcn5Mfy
dH7taZ9wK3YyNh0FJGGIRCndJYik13lJcMo2Jjm/CsSavCdOOD/iyvJjOKHBOTDQ
77aYWeahxfOg54J3vZkKdGQYKcHcOxER4QRcActbkR80fEO+/t2u4qUticocMBEp
OVon/8N0JlGt3QTNby0qb7f1N1lyHrsNoK5rKDOOUTGEbRB7YJE38gB+TjbuEbVc
OT6F4x+5N2IUJg2llISKrLblPtPxRJVLHAiuZ9NZUL7FOuYDFXjKxomnoB3zHnsr
tvJrgjQR+PVM+PJi1AgkUKHkkmB3molFc+4AaNLC8V+t6ARDOoSrqvCsm/TLq0rA
yBcVFz96xwx9JZaUbVMZ1RoMIJmXrEO0ojmveffCZrzQhRluJdeAHCeS7opWOZru
np6zR+0SlfXXBT16m7ax2dNxCsrBIlj8eITx4weYWk0ZtRSBU7XaHmQbEyYfmsuC
8n4rouVkGiY9cGpHe6Ui9y+mQIYxLLIt+d2VYsVWfQfKN7jt/AJewfTUwIoDurfU
iRXOzceuWvi02wV3CY2pX+54l6uPYbqyjSm6EhbkN2cOojkb3JFcOcwW6Wr18/b0
aJynhWoWc1lt+tQBGXd94E2OjBRw0e12inYCsBg7xf0UccI9a7Th+OB7MLwmE7f2
bvHhGlbp288YhvPjNpUaNnZbBrdZi3t76ezGMoD5E/ZDuQEn32+2+dZhWiZ4wR01
JtJCVNm2D1lQ9wqM7vv3klsU1Vw9PW82rg9pI54NMbVzDerY+pTz1N1YfToBZsWi
JuGu79+kOIt49ZjjBxa2VUnv2Ko2UE8nqwpJl4Uy8eL6NuaGSns5X5Rz2BAjiaEK
VDw1bwbvSgqRp5rEdzb6mAh7d//sQzTPqMsmmz4HdTm3+tTT1nV1JeREqgTjrIJU
JcWMMcb+ALZb8oP5uAqdW08mpXTkJpyP/TONY0Sz37FqscHQA6NmyfNZsY8RNn+2
ijmaA3wyGfTPaCLFiTy9HksM0gT9+dX0DAedW9DyPXuWRnoXhBxKEE2qWZPx2ApT
4DPNPBMvRFzRYf8kkHiYxtsgHFk25PF+eHDunvnawu5Sj/ip2mjXUAFBDxVN7Mij
BTDzXRYF75PssPX/9L0FJbJm3cKvotlOlrPICUQLxh81ZVKlGASpSds39CGVEhP6
Oc3UCxvAeY4h5HFfTorPPX414GF83ehHw3zAWfLt9luYjXd1ozlL2+FDPGoFez+M
HWzLyYIqFObyAe7ghN/4UBZTlIWjU3Gh49VRcwtS13YyueonjawDM9qgeapd2Tpy
ZCasrpVSXQfSbEmxN6HwMun7CKvMOZfMb8LSq12kE0keekjiDLS9PhEy8RQ1oOl8
fBWLaaJBAzz5MkDOf/MkJaCv8hL3WKI4BRYdRLmyEmkTCT4ryz11m+xqrTJNIlX1
Q6eJPgGxYR553VhiVihn1/xmYOn2qPoBR2DvwBq5ohyo6u7IU8SNQKc3VyDZeImw
/JpfXO7Y3oZJcfSas0Sw31npeRdFbv1b8diUdEp3ZRva44yUae8B2TsVfiWCKojV
MdRsXj8CxnBXjmjOlvhyv/IiQMgX/zl1mT5PMjWf09CvdgAo1y3fWwMA05Ee7HSk
Spn4UkEZp+AEWACnKYTimFypZg85bTV7rJnSQyxg45LgqRptXJM9mZIZLZM6gMWu
d9CL39IeUowZg4bYCtyn1lKmWzihhUUDADn15gGfkQiOMn+hVg9BSnU6jq6d+KNQ
GawTaX2BITG1LPYrGOJnYp1kGzDkOcQ5CoTDWaQHPMlGLoJu32rvX/LLfN2JozC8
3DfDcBN/lvsIRHv+TzYZpa4YwjZ17LpCsbwABt+1VN1OzZiqNEF/NLmk0sU4is+0
EsDoHaiWPwlbaQTRWMtG4AMJXiMGb+nTO2eH9NHhiV2PskYkIh4m2/rWGMjzPKVM
MD4xyrBHa/8GIh5Iq4z2cY909U7HZlrnxDJluIg30/jmLIL1duFgDSSFjJQvNFXE
4flt/5R2z4OuUIvQYKpwwttpzUM018j6jyLhePM35hW0nwdQqQtELnlTXRklj9s9
RwPYoIssB5nX7tDxT+XcWupyheSczyGJmfhAdg8Cect3HJr9L+NgE30+LXUk0C1Y
muO6pUwcwI3bFQ52yUdGUv/sOxQ6aoNMBVHz3ePoNydw++/P1lNv5OtnTaLMDh09
zo4Y1jwAz22YSEL6Bs/VC7J2LyP/QT00bp7Z0j3LgQFuS4yF/B6ttwP/At3BKLJ4
fQFouunCwVnziQvDx37RkStkjuhPdVEAnFQb20NLJP6+e48gALb78vdRTThsZXjO
zURqzFx0f2E023Ld46KtdJCJIu2oFOqIVXHp6vjAmyolXTD1+/B4hqd64hoYgtZy
q95Bf5hlkwzIeIwiBzK4AssvLwMY6mIZjHWY2z+/WFTiBmYvS9MbAlBjYVdw/Ok5
V/k7dS8q5q0iA5xPXNABEus57kzLyg8vxAwD9nAWgU25aDfVhXXYBhYv3PCgSTY6
Ba7sDg8wWK5n3wOUgZopEx0jAjrUVg6oQMO3UvB8Wr2rX/ZTRII/mVuKEaKY05pk
bF2smkIUr29xPKCwrn6EEjhUTERIiL7Tjwg931qQBgKTuioffjVjCQkXk3SlwxYC
4NSvXlWxv2IIrrVOnMUaJ3nUD1osrjKheHPb0rsq04hB/7mhLq5X6WIeE7i4v/ry
BQcbRpjgDIKLwWqFFRqv8H8rcmoerVyy4f2B4lHXEAMPWZbDHm92JGFXdQBIsUna
gkfC6Dj5OcJaikjaNbTl5WfeZgZvH4Z7LRvzc4+NHoCzUcsnReSmE1SwIx3rvL0L
JKe6G8X2+bOqdmo1HuNtfWMBGn0yEu9/uankjM0O7p6qVTZdrXBMCWcNie4fuv9L
xUtoSw++GaAuFa6aRhWFR7XGuV/QqRjTYQKLfjgvm2wD7fWX2TUwX4sqPAdRhBjE
tN+PCMBpjmAkwo1Pew35QXTfttEQTSFp+m+d6nud0Y3+1zAGMsbY6YmvorF3Xa/V
IiNckDbZt2QJeO8Jpuk4CwkC6zC6fgqsG93NSkMu12usGikGcG0gHEaN4ouTwWpk
8sVs1z/nju6HUY28FJMfB7sBGAFuoksb7h0Cgoeuv9CLY06ckBafK/XipGb5Xp+n
dvnDYIHAN3PQhTwSTxpJqvNmPbx4BI/YSggGHdqESoDozkspcCb4NtGxfm23aPbb
EBkmQRj2DiqHae3SfYz8yStiO8F/FQeOyrtyxTW/xeq/QjKxW1fnA4uIBu2bnWTS
Ztvzn6pjudIv6cb8TScaFjkeLhyL9bgfMVE45coACIp//AvzaU/BvFKebxKu00RA
CmSLprd4TTxRZo7W/6yv/Maky4e+xYk1Pk8LbFKGWj+t0mkXH75g1goI34JEFvwB
73053JzzCzDaSPt2Zl3SVBONqxu0NaPQZapVV9cgCARGOBX3g/zw8DKycdBDzx/s
o+EpU1WD56Tmb/HZURD+qC3qeTuhxbq78NWxdEzy4CloOfzxzeyWAfN6xiI2iMSf
XUtPOXK/6LUirG3fzqNnWj2Awp/MUylTYbG0mFPzFxR2m4klxKRkiFQQhm4KHytx
lknD6v8rdGU2z0ae9m1voKq+j3YeFTCFLfFMiIBI669HJAgNtW3S0p3EPY7W3Fs8
NpjfXqghkKZMOtQbnWJu11qrvNu+eLqlQ75QNcl3x9mYEB1NrTFk3zQutSkDOAab
fegrtCSuN5PJm82fHp5X4lFWm4hKLFzgEZfLY+5Jp9IWZZswwLrlzCPsToyykwyI
6gM1n7qyCJ/KusD5DJEBKk7j5HfgdKT5tOm7fnyBz7B3vR1u4kff5apnS4ffXztQ
RtqNutqY+m6dr9zWscoIuOERjW9MSFdzC9JDEBa09mo89Zf7lGGT2g2lrHcvqE94
n+BcRxwz8d3FXGxuQFOWL8lL2GSCgjJJlk8Kie8KSL4rMoOiy1UrrV0FkU4POXBD
64DwCJVBbzYVuyBYJ9LpQ+xmmzs0vsjKbZS0yH08kAwrSKsBSlXgVycTWvEHgCF0
F/Ym7W+ibvVrcMZgQniMpq5kSYsvU3kT/23heFgGKMCfEEbaUnxYYSWsjtXnxts0
vuEy6XlUUnz87GNisXOm0Q69yT/8J/VgcmEPnXLYqZ1+qUZ8jvL6LHDJ5vj/PYP7
D23ogHK68xNm4fOzIZ6eyZDbGkTWX/qa8EQGgqkbXo4nIFiQm0LzYqNpBfRbneZ/
YPFCxgjWoZVlLKQKmjFN/rGvTPcj1DM+6ejK1pIDlJtEOjIZgKZzHcQWlldEmLzi
CB7aVDmhbyMN2nR03ckDiA1+XHxEaXjzjlcZofEYQIP1oI5OjFnuw0FxeW0lV4co
ZgX4BkUXGM/wZgcicoynr8/ndotSKUOC8ak9s5ruodBYKBGtiJsouGT/tu0cfkQP
05ijdC0LJvqB4UGqhrFierLDPWIJwi8lUPttu3BWACHXRHHd5PFOsg5pSnckFkZP
VQtynQ9/R+P472JDqUsR5cs3p+QMG9s7fWh4hFFjNgNFcqmMBJopVJ5+ZHfvNbpU
Xd211Eddb06GvNKK9OuaUhBpSA8S9w9j2D4GXyWjhBhDHhZneqYDNbbFf0wpfiy3
NkF3PMuc9JFWxlPi3Ds8Aqn+TCgL+gubS3p+E6pcQasDDjfKoYV8nb5iWLzpu443
vrXnUnRhIcBoha6YcqdLkz6qXTPdgAfJ92pmnVxNthic3XAvvGEWqDgOycW61P7O
dHPaFKc4XggJG1PLkjQ7d7zgvk4JN+AMQ3Orm48PR2JqQIZdgSZqBYMtLJjbG2eS
KkkiGK23382aiYwbjZaRFthQGYFl6c+LZSKLQ8ROzi8KMLzL89wfbYrtuoOVy9KK
OEmEucrj+kfRhC37ykO6lYePU9GffSM/lVnhYcMJtbQ9t/BgXU4hgeEQfxnPJj5r
B1yc/5HT5LVpuKEEYHIvPl6/5c8IBQmodhcYeNlHx2ZpP9AiGnISxU86VHyAtRJl
GjadhxfHp4h4Q74sNkrV0vBpq5/GS9lu/97jr2AVo7Jftf4wXNGUPjU9uK3v2G7T
cxJu1gqgRU0AL0W1IlK+EVdzr3npP7Cw0RLyUFSJcmvRqkq6DjxxckzfwOk9RgAu
Q7OKZRYgyx4oyZAEtqE3flkgED9PBILvJ/IOEjLBXF2Lz93uqaAlvT/WE5fRXrgH
dtxw8yswkcTCfkMUdM0NeSodIeZo35P0a7649vCtAtm2so6PATZV0O4uvtfuyf7g
ExZ8q65cNX8S0tUdY6XeZGqTKwhWtqP1gmWtSOce4KJsvschVVB7YSGzoyctLf78
qxL88FgMx41fDemWyf2ydqrZMYTmKuPy//Qa1P9jPUbUjvrcX8YRLgldCzVnMAoq
KFzB9EeWX2NaEkxJfu6Cw2yVOjfUYLu8FdWyt6kyUepAMkmqjSRzJvPFalZz6VOz
gICBUkS2722gA+Aq2iz9ZEW9yYNXt+FqeoCoWxtHrw5TOV8aMFUbmWc5+f/MUIVl
LmX/PYnxxUKRcCpgXhUaX4qk1JJDSd/y2Emm1EiimB6T+aaRlk2aOnuM5pAVTTnp
opxh/6xUMEhKloCR23L5FVp3iQrSkdTSabZb9BfA+7S5r0cudgvHKWTs1LajlVUX
jPJOCnlYhWQHVE3BzJovlMQSpzPzbFTabtpyr9lxoJ65zDYT7/tW6QkQfXWlbu0N
OlVF2VtjZLUHJhLfPfoRqhrknJD7FCv3u46KOUv4eNatH/XyKRkjxxFVBslVWsW2
q/uHBRTVnjw3aWiapxRJEX+CkcfkjCx2buNCJRo+ON1/uSBVTwPEaa+XQrpSSMJ0
ZcTJl1BW1pCXN5fTQfZbk1p0d/QXMRuMfFNPs5IE3A7ODDvVa3DrxwvEb5OrzOOp
MXzMnc9chHo5YJ5FC0EYESG3DvZyBzoHzB1N1lsmCSt10Sy611TuQXbTGIjG0q3n
vvWjhiAA7lkbXcHfI3EpZnYf40+ljxMq5cTrntBByt/FLSqdbvd47NCrAlxesQlQ
LuFA4pCS+AL7o1gCuVpCmPZvZvq5nz82gOBngLQrAdAeMV+onCfM+GG3hxsy9B8W
YavE6Bb2oQjK8o8u6gVm/UHADudgq/t/KHAXa2mZU73sjqWAyIkaCuA9i4AFAskF
UbXKT1ClE9vL4Pzf7oyjdODN6xp1ZuSWHmCsvGlQqQkE0b+lLJCizUkEzJqs3S8U
8SV3kfNe9AtZ/J74/UVxHN/2sEclK05M1lDHZ0N2+Oz8UtXDk1lRXE95ytSBG492
+DlKTkWshiLAlK+GKuw2TxlhNUKKNZeV7A8GGwxVHBQgI1r+VtZONj3yVMA4ihTk
3ywmLfr+7ISha0DK+enYfMHQC1rMmO+xgSAI/2S1HcCTcjw9aIuYGXPYJ4qEEnet
pJPDSH1IpxtQXsrnVoaBAQNxW+sHWw9P4CnwVEHF2bvjRY8RZqI57qyPpl9XITub
S2PSJZzxPg2WxwQq2aK2UZsyOiSF40YpUKeomqju8KfFnX/7pns1RravyT1yNFNN
1HCt7NsWprx01QCnMhtjhaY4FHX6dotPMw+SNFagUc2h3T3RM3Fi18RMSax62u4x
ZARUMLBruCV3nsZbyg7bG6CMfIqyYGant4rbSiILb4aXAuFvCrasv5GTufYTEXyF
9WWEmmrhiiYuljH+9DJdX4h7MCX8ni16Smvn2dD+Vx9phOP+CibkF5CrRH4nYpmQ
gFtq4AdHq57yIRVlFVS81Khtnyh2aJnaNn+Ue/v9zTcCONwHF/KXHXDrJm0jLkfz
e2Z78BpDrzMpCLj0tBUoMbybjHXxgyakqf4Bm+DUlSluHy0MwyVowL/finud96JP
ybKYVC1yUU1mrKCijBtvA2ewzLT8vPyKvacVcpdobc/syTXkVmf8jALRT8W+FMA5
H/BUGT/HYQwixXZHXdy/BVTIORiZUQuf7B8Hi2H2qIGInvZH/reU0i3HK8v4Ss0+
5Vf8LFfQfB7tvqYqw34BgJ2CDw58p6PMOAajAQfx9dxBi59Mlhsz3ykuHW5nPwBO
qCjXhMS+8nTfSboQ4h0VcmMZdEMUg7FxEdEbxIp002Hpkky3MDol+LFGbWuAoTKe
NdWMgdZSHJ4+Q+aOpXi3DqDe/DV/40kQP7XXqnTCRh7XAtblxH1B8EnzQWsY21fH
sWoYWXzRUpWvzkRXY/0nqTwb9zGBu/mKzK4+u+mkkx2T3EEZm8kU9dd0FPZooiOI
xxWqijISKnVzbpss/DEwRF/yw4XSvucorH3YlCt1l/+4sd4QPcT1BNaF6I9K0yKl
k3bn6osD0n22sEn5yCBri5VcqoJfu1VNly/fcs9NtzQoNMltD2Xe179+t1CZvkzE
vYDu4qdD5VLinByznTVzM2fpciiqSthUUBfw8PaeJDZEK95wNZMiW+nAECmawtp8
ECm5yyQyHhA5rafF6lVZddmrjlhCqCn1Ol0L9NKnXll4slvtDH0M+zthJiwez1w8
wxLq1PwuKK1FuOX2jPKnh1H+52BHsE83Vfb0ucpQF4KbmQv5Cfi7opv5w7VSvsZE
ZWSBOQtQB5DuhZDScsOS97e6LtdgRDUFQSZL60WNE3pydp5yeG5rn1/vX329qOYz
tzAK3ViXtqUmWA6ZXkEsqzgUSSHGrxZDdx82EjcQFr7Y3nCYn6tcCqEXDRiRcH00
ccv8NNuKZFu1i3CugsEZoAKzsXyS8If5aqXwX7EjndvKSDBU0yJPRqg1V9rWp6o4
mPOGP92vUSgCN/xCJIxxnLUqBZtYFyVXr6JmE1orjaJX+1JSAoDIgDvXHfmF34/m
HIMNrCXtUfjVSvlNLnpZEF9FrF2Q5xZ5+gz94GzoJk3k05PJflu7MMl2UlalHeLs
j9+1S/MWBzPtomawWCCJv7WFmaiqpdPa679R7wtQlBE3pD00CQ8JXzXULbj6KkoP
wbLUsxRXJmKPJshErf9VEO8VPxJ1FLYigNUUBqUaTKeLkKgQOiRhyslcWTq8xmsE
UcIQEpn4U6Aiw0bRfE7jeGvCYTG3Kpzjw+NvsARwufxqCtTHrtjyqfSH8AFHjDEg
YRfTIl0i5VwO+gETaCIT5VR0IrZrJ/HCmwRN3ONkp9taZqqdUo4nmjsiKwpfzisO
6YA+3O/1kjgf+3gd9SUJxSTWsTbqurbI0Qvs5Olql2/8EgdpKQKfm3lxl1eTo/Yu
AajZClSO9aoWC5sWMr3TkV/CvSqdcJNzfKbmHZIzigAtsi6b3ezomHqOuWMBgBXk
OWQGBAdxx99JaRdfAUZzfXnZQDFHZNZjJFlA9jRcISCfDsPsJpsjzJD8nz1li22X
PSYGBNDpsWDQMNMTGDWMcvnDO6I08RlKEi0B0eop8KjXqUskzgSXfMZWInMBUVu2
i8R55pnZX+3yuxudVHhJB+vCibIRB37bpvXcXu6UjTJsA3/yA/2d+CvezWkte0gU
FnOhSH1lLuCGCopeH7wQ6UPFpaO+6at+yzq3WUGNFsrdBC9zCuQw9g2mAan2aNg5
fY+/D7cN0IlfArnnuGrtRBlrIsPBzJf82RqRkFJQkCg55ASp5n3j7sGQo0erDhyj
nAtPbkpQT2W1Dzq5nIoykUZ/rmnGKO36+/EFbrjlVRYFwA4eS0cy0U81JdGJ32EH
PETTw/f40S/O+uf7AolnjplAUxNuskduVNrnvBki01CrWutUnKAF7cnTvZTfpnD1
oFgsLLZq/DuJ/QtNxMij1g7SEuPyK3VhgboJSwofnYxQ8HGhPaj5ItO3vQD1n7NU
5Wve7ETnDUNUd1ZsAVgpYD79ajrjZijny4nIR4VwrXqhHHqNe2LITAfDKe8yZSAb
mST/a6NqtfzwQnNNeEut4/ZyrcrOuVd5Ejatlcg1ZpqS8uNaixhuc0bRK2u7NdbJ
LwBnIInBnGCt9F74lBoHhXaVAOe74elVf9BKMDI44Gfhf06KM/Re+QEWH4hYwpvX
KMjCagztnq0M7ZY8V7PhcXBfVBnCw+Rf1V5VbhjVeXuW8tJUECQujVoH5TcUqV7v
v/sKpfCIKtK8IQVyq9NqvQzVr2czH/o7HTwzKQ/mzqXwixuyNjLU2KkvJvwIOfD1
DGr/lMGGqMp3zwb+x+UIn7cGYaAsO6+CKlQmEFgC34/R4sYoCqhF2Vi8WRZ6JCjX
ssHshSc8+JX8aizMfwA5d+fvFVGKbXT7Kp7hdmib6LjYfPz2I+XD2EEATegIw+7Z
/a9pbY6qEszZgIND1F68/grRlzs34HT44iIawBy6T7tAL5FbdHa1GSFD55Sa7hIO
/bYlcumzsDqc9tRXdnxG4eFoq3+63fTo1YqiHmF1+ARRk6KMxzEkhE6xf839RrHw
L4S9tVGDSTAJs5iC3kH8gXVylnsdFFhypAVCLASXDi86w3JMAY6e9C+jWB7M/pVe
Vuy9cyNNYfiRgjcbvmf+C09BN3OEuhd5NjKGDNKLG/zPesq5ThluYoZbxqc2Evuh
nM4J5pyadnSTNnNKOtu9Egw/dXJSVLKfwR8fKCxCvziBWa2QAQRYGDRna0mv0cl6
Nkk4W6t3GEJNNYTBoY2EgSXwlC3i0g6gTOq9kwBjC850rnUsO69c/fD9r1CFc6zS
H39Bp7SPNPDImdr9aW9cyfzXzwir8ClVBa22eVbj2aWR4M5KmiPVadJSjOy/YIbL
hrDJCLFK/9N94kY2vkdIZKR+ryZsG1CXUsLBPef/XlmZhSvk4YWNkeeJfJNBD1lk
7XcCaJIzYl6l+Z1ywSNVXh1xSCy4fsNP6592KCfMVsYlJgicF/GKGCsE4rLJbqxb
WR2yRQTqS2gj1/nqifj7458UzFOGKOSdlH27p6k2JI1AgmXtgMGvOJ13fCUlxKvG
KVvI4VYjas1BNu4jSPknSH2OlDB9Se5BSBpSVYw3Q9xSSA8yku7/TBG+F++9onOK
gCE7kx0Siq1bHHmnSj0tWRep+O87/Q5TrDoDd1gLu5iUDoqKuJ+H9krvJ9FjPU8S
4Fv8mTS4zxpzpiKtvJFQW5iJb/BS7GI1eydlJvk+4+s6YSP3WipIYleTPWwbWPRg
I0dmJkYQkVaUL2A+t5ouQcbyss85ktDqLxWrPsP8xJmVToZL1UxKXruJbpKAbkKS
y8d575NYmmM8pDgO3GsdjxEPyD7FN3hwRlhupEKhQyczagWJQnOOmaAW88sCRfa+
Z5RWBMXnMh2Tuh6pspAy1XgnqmdL6LLPmS1lfACe4q9R5a2Z69qp/0qKfM3eOxIl
P16eduqLA9VqUGBaLNJsmsGpnRX686fRIkFzRJN4CwukG1mjkC/IJtAYPCu9jmD4
RS4VFp8jVYrUCr76hbSeKxJAYg5bl/tsSwUFJtEfO1SuMW3OeyifrrCjRzzqGh2f
oQ1ckIYO+TK9iEpo51PCpYYXZg55HHrfPDCA5yCpRmwu/p+lhEe20O+LA9ehVJgj
V5ZxgVSEM9sUa9H4EWans0kJhSby1GPRO4Oa+KJjyrJGLXISK9OSnguYB2rH9XOR
R9iiJJ/CULrSfbiZ9+TM1WvFQijER1hCRn/N61U7as3I01UMDYWEuwYWPLZt8cSs
iN5tsQReEoDFMMvkig37gBqruuqimNL74Gq3bmLRX1oJXrgiztXN+BOfrbqkvW76
egoY+j9KpYBwbFmuqf5l9Z34JhA0L/vadi42oE7CvY0jz3wI0kEpFAU2p4GhwuiL
Qm9vCVlQqwed7x/AhQaUCuSKshE6G1icjTshd6AvhVY9T37UIxna1mT86z9YzxH0
qx4HDOiCsPf3UHX5noNM8wv008CYimVzECnLdMpCV7z/I5E2Yse6H17gM+lYvosb
gNElxX9nKCS+hOGdsGqGWNQVpivkPUTDvkATkTazzLQaL77fsuFZXCm2pcC461v9
sO5czgT9mCDTfv/ZCbFKiyVo67to5Mu/0gGjFZEV6hhLiOzTbkWWHCDPjTN4TuX2
QjzmHSgLZlx3DYq2baBBfdyi4Q3xncBop3/qjN3xnpAj8Ex1sslIR0ax1HUzVM94
rz3UxRZI0PpGRyTCyDDmMBJ8X8l+z5KoPEteGf+EL1L9FVm57skvP/dXOf2V+4Sf
2KYppd6yypPiaq81qZUu1PxS5hNqQ6w6ay6IFDARHYWMOMDeCWz1GA57ocgp671y
Qn2wBniysNTUXIeMl3E4Qz4KO5Ys69AOdqdvn85azlNuZnLGvT434i3lEeVxZdhm
7+3txlPUTPUc6ctkQ7D9ISVzpmTSC9swTYUx9Ihju6ckBDYPZmNzDbrRvtHZCDo2
Jn2kyp52YGHrOXWhAe8puB+lzOvBT7ADzWblqX55xfU2cLkyNMQylamPT7y+YRBA
iBSGS3NxbmRzdks0RJ3j2tNOLbwVatiQWEPVqctYASrT2vIFozq+pqZbBfkyWIre
De+uRVjMdZvc+mRO55NS3pSXc9Pqs8U1oORu4Z6CYVCE8/eSpmZNdOgDUhG/D3fz
SLWq+t8GvcsTVocN2zTZGIBc6rHR7YXSprvB3PirzCPxBCaqnuWCID/TuL4g1lB8
uqoNJg3VSi+DzNWRIs+TVcpZA78XpSXlluYmPY+tmsinrlV9E9Ax4jS9G5zXb9PI
+kcRdiM28OolCE0qN1AMnUIduzGreqBi2TLFdiWFXZcYhmZdIMF5Xi8Ipo7ZuQQC
i6spHWsGELJFwvhe8+p8FSaziXgK3tefEqIM6i2a0UaGcOWEoOH/ckHuFaJDRTrt
IhnlsSHJCCfTEovBKdSDWOO+rmwo9o+s6WOWavYBWZYY/9/vF7RLAklX3JRkIHcB
fpW4wxAPUZgdqhpFFI98KiDW+2GOAmyaZGWfY1MwC+aZqNqg9BIBB9tHy6a6PQrU
ZfGSL72f4f9I7hntsNyqWrNjMd/viOlZSSsifAbKDlC9my/uS8KYgWU4a9pvcgEp
k38JWGpCp+oOn+ErGHut5WG/Y6mwGV4PLQyjZyvCmdGJFLzQe4FmTniCcK4/HoAD
wGa9Hzxq4YJSogeWi8HUB7GaZLL+Wt1GpWNV5TOjUuxeNbHnLNKLT90+YnIospTv
q3smYMYMwCe9W6EFL/PVJLmKPdEa3ZjpN79furcasgCksTqhcjeH9CCjEaUToQ/W
b3gths7knv7DIC666ltoD70zFCC3scQt6D2W1HnpJ2+90VSrLuCshuhPc3EGnEzv
CKcs7uD+ntDvCeHw4r9X729tN4hsGqdDtxgpvgEHXYezFrWj9ponW3pcXrZCgnB0
bKOUEEWa1Qj8xPN5Z+/bSG0jFZ3omWJtMZtxKTR2PlswrAqZPav5IgS0N60qgnGP
jD1BvTe1DlLKfBIJaQoDCeWlCfSrN/ISbqpNfvBf+KL2R9AqlvibeHVQpzF0A4EM
vSohXh17rj6KXP0tk2qDw4wGYdRM1WKIFjOZH4C0pYdjoXZOOu9thLKIPtvWB2nG
0VAZ7OQdCkP1a9fDG5HCW+Ypj3BYNb8VkI/O10P0SrAcsLdIFriCH45E1N+duZFK
TzawnNHaGMaNMH0VYXmMa0pscemtLFtDXbovksXwMD3Ei0c98+aztpW4V83C5CPl
twkDkujS+98naAqcMvZ/T06ky2TURDGXyN7V890F4BYWp02Pcf+O1ivj067Lpviy
/FPUJiNfXrcl7h8s7KO10oMovk7YltHsA10Hrpx1JtGRBiQTbcn96x2XLy3g5VLz
HZjtwfzJ7OPAE54AbWXtSPB1gy8RbJCZ+aJ14LO604gXnK41TaVlHBKPJDG7XmtE
c9sZLoLt6lLC47LA5XzosMQ3krjqShfxzShRM6Iwbkt+PzXOh/ZEkSfL0V488XvC
ONqNTd5y6GFctfEUnbO5xRsDNzULu336Q7glXkBODchKavyPqn1Q/oaJDcvBmWQz
U206HGDir0uSXlMsPgBf5Cn0ZdUWzZ4sVGGBCMsGECveWu6exQzGyP97/5OSEBmB
fbI9mX6QvWYyO8tbqBGFsQKeRtFkc6NDGTt2w7X45gphKhtvcRr3fh15mrqWPC4M
j3h0ivXOdO/GraJ9vklIIPrs7Rmy89N1Mj30j7av4LMocp1CGcqZRk+m2ODku4OF
7U0cvmE+nQU4lORno5eENtF/hqnmEcDZauzC02L6zqjqEGhjajJ5uGnJwThE4KOQ
GTLL3H78mQzLLlbasMnn4MocHS6eMeZNxmP1hV+T/x80x8nDtcoxPeXm5hhcpOtI
McjcDWpMnewJ/9V/jJlJx4p0sQ/DzdpStxgvFpDiGT2VeCu39iA0XCzduoMzpjtc
qsvBUy541mnoAdWku7YrsGV2iDvXxA1T0ao8ev+zOjBqwgc+phGA6R7FvMlKbZck
UEOdBcz+tRIkT9suctzOYpCFDmwvEGzPWf7/Rel4obbjJkv1KFiAWMn7O7y+/vUS
YuVnn0xM2Nsy/EGtMd10PDt2Q9JHDuzdb1Q826nzouiqni6OMrxAc0HGVlw/pLe6
xrhhIfW1GHPY5mVpVd42/xwj8UI2UPdl9o344TQ8mCnpMB8yVlFlk0N8V+7JBHTt
LKOBv5rx2tEWhz4hZMibFY15Y+WLroLIhKk55qG9rLoSs6Ir20vquvI71Wn/j5lL
dmbNXc3aWpVD0j7yXU6QShXM1seh4zf034HHRs3qbcshk1pTHB4MYBDjeTXIBuP5
zJOrLO0vanhoLYeNyVNVxxZSqjtEdyNi1aPirZA+PtT1hyUz72djj4kHPjzCfECk
mx9QnCnAZcd1GKJ+oP7uMSja2GiyzKc7+LI0x8AadXvOyrJaVJKEiDK1KVm+C1ra
W22BIpPgB4aNEZ2dZPtMbjO2nV4rYUF6EyJ757PWvtdkZY2J1J9h2DUXRnclltKu
fdSEb5KDPjAN9SFTNEUcNFbbHuGSHIDyEGviK9x86hsREfCpONvLt89COrNeGubY
YNcuRX3njHIiiFamXsbfdGPgsKoTK39NbHAHZvYP5XcfhlhD7tXNVM7YC910+F1r
e0wT8g0eY+3/eA2zgVgXMcB+zzEEnDitPUJKJ5Pv4p64B6NcWaAOtPCyxgw/OEeX
cbp82bNhpU6/lgNvOIPQQgUk9xyFNjyrwze9vFjIcQ8oeGE8U00MbQmIuffK9XYr
oVM7va6yZFIfjgB7KENgYvLWQ7Ek4s2bhnFtM/DCmWIWyR/chezt+G8vDXdGEyb7
78qOrdfdc6TLVgl2RZnUkPwr7Byb1ibr9nJsksFAVNyg8lx7r8Ni8UxhacqZLZrQ
ZuPMld9s0THBLWohRe19uIrU2ZuFrHfbxLwjSILohBR/M3Xdv9b6Eg5dV8eQpPsz
swoOWSPuzhSRW3oq2+q7VUuzAt7n0b2T5Wt1kgDXdu192ZXNVwiD74xXhtoAhb2W
mpPs1j37FpNgL8WPEEDoMQ3aS7rQv1rdpceW7Rm3tTcanYVtO/5zm8JfOfqgyKQ6
a79QMF/O2T/jeaEOePg9JNfn3FLfW7x+CJZD/KoA5ax19h9WifnCCtceMdzSzbLZ
j8Qv9Ohc6j216VOawwoqk6BMvzYukj6freAXx+2OFenhNUG8sDBOVL834/D2e3UI
xjHWYKEJK20zSiJXpOF5Z26d+zMu8smssioxiECuZCfydzjxvWb+BYgpbdws7+qN
h7B+w5Kps+lwsnOR4YopDZ07gooOpCjsVXsge+57oOJKqzT3L6O7zcWwtt80TQpZ
dIDRkhe51dcsXf4zDEPxMRKGmeqYD2FYfF/VFLycRQ9i0PQcD0gbBlw2efbjERbM
LQv4eC+dwlL9SuFiSIHmPIAHTbnh/TQcEOmUyaamB1ri1VVsUmo6pyCmyGpd+hMi
VE6OlqKTEs1FIAqxQun6StWodzd/ixUMIuimqEsAZfC1RGwxIj9K+ordgyqmvnJj
ifh6fXNbSsrf2/IaT8pFs4MTXz0JOD5yoJ9vigUlMSZLreZsmJdF/fw1gj9FDnWh
khNyoTxtQssGKLpATBRIRZW1ic+oRFmydBsbxpvXfKM0qWoUup1gIZzugndW7urs
4bAPZLQyLCy4s5AeDQVAuQVGd0SyUnXYjkkC+RyazTDLSjF/2d3R2uUn0Fs8HFYR
0iH/1gPq9Lg20iz1vO2lX9dtKI3rw8HPe3BmJKUH0Mv4PZCOMsjLRxFZcGA7zJW5
AQnhWUkCS74avUXQxTfxKNBPJesLZAIjEdoMkhXFfcA23/+l3inkulPChRwaSk6f
MQwphzsloR3+Ad2tBoUX/AHjxgsZdSK9EWDvTsYAFZaydV3RdM1uQZPytgozvzHR
wzUZloDt+3PgKtRileF75hYd/RIHdCybAcQ/l2ss3GdVkyeXCqJAQdWURKpcg3nz
Mvgrz77yT3mOju807ueM+mHFK48Y5wb15tb1hGl5mvaT6ccHGaFQVrCZ2OPEwun2
d2lwpTeUaHBpadVJM8p/j0wwpKUQRSB7CLUsYflV9bCQ5iBwB8r5v8DMCk78UJkN
ByhmhOOYs5doRGkJHC2Haq0nJUD1+s59dfAuR++RsQf5SG+FFCw9qNsswUw1ZOMN
376g2F5D6K5PMK+87DYmX1VfrvoZRmY0kt2GFPizqjN2lEcGNlq1cwEIO5DIEQaS
q1MIgb0/BHG2De8uwfhdHjbaAcmLHqt/Pn5fVDdqMM4AzUYZUloPfAWVc5GcLLPp
+Us26juuH7KVmxQohyKRchIRGRM3c7+umVhLzygvBYTAoi7OJYUIWxk181ShZTwO
q/4hkgeiRfM8+Kr9DtrWYU3NrEzEDJt0YM7GVRUTTgYoYoeUVlnMchhoyRRdFjJX
PY+v+K4loFPhTli9F81Y96rHyfyWJmSVtUzjwiVs/wP8JunTH2YcieTCZ2ApTuhS
Du836TVrMctDGuYcedlnhD38KD2uivYRyXTNQudm7FlLdAejbuu8I9iPNx6/7DJa
TEEEDO7TZh4fmugMUaT0h0uvD8m+/tXJAoPVHpVDIuP5trjGqoA5tEJu964vDFo3
w4XVdrtLITy/3/ZRVKJlfZ6HERxxlkWAMatNy09AMuoirM32RZiF/ZAoiMx9xsLj
R52JPv3u4B6uF086mKeyRovPMBdyRjoZMi/GjJHChB9g9pJfRHC6kY2RFK7ULhT2
r5ezviMFtBk+b8KvQZr4sZJb9nu+a5OVn5Qfj58vijWhyRpn9CHVcUF9ILiqaSdJ
ND0Ja7upOOJy2qtnM+M/hGj19ReEiuTZbz+gN3N4RPqrXbpRilO/Rs6Bc5jddxpR
pY5bs7EsY9yc14K5HpksLleEJiibolGiIW0nOFUj01oILZGiSAWCmxG3sFLkCTMG
3k8NpSpf4WL5Atm5hUlx/xIQIBCi2YOrmyP7o/S5ni8d3tlMTdtEGA8Pg3vcsQTQ
mY0tmeL6I02DRkQi8EQuuxWYYqeb5XE/OHkl8oSWI3vwK6iCZfsNdzSHCOm/E4x2
Yf/GAbAanAlGT1VK3GRmdlHJIAv+b0o+sSDSg4xkpXMZtKg9/Q9A4STS9j9hw0FQ
hckf+l5XeN3LmtVKFUH2sW+8FosAg4cf2TdKJeSWy2deHNYxVpy6B5Wh7bOI+WBe
Iqm/95BHbmazwOlxjUEOZcNSZ0noEj1h6fGS8saPIUjbZkU2KReU03dmt/TbbEU1
vLb2SoaBkxQxD/G1TttSMgf5JTsHhvtA3iGfZj4zsTrDlA4ZstlsveJlboZ0mJqY
4OOHKYqmzy36ll/QQfVPQYOgQQMcfa2AfIrT72rJGLAT1h18kzZ22wYw9QlYAxHe
1garKuMrjYUn/G4ZjnKtk44L6/TWyN6fxHe1KbVAwDq15DIuemKCYlmfkIfa15lF
Dr1wAhClaOM6kCmjwe2eNA7+ieD9k5c8fABfif9XnZ2Z62CjFntav2HP7n6/UhfU
QFuhug149xZaxxPp2kEsGlv9nawu+UCJv0ziv2ZIMJGxCTFWaHCzGiUXH6WxWqPo
6HjgnX1kU6KEYNG5MHHPl+xO717j857uWmOWqoHAC0jd+JMh1gPi2Ky5FD0pj/4E
n0uIYtH/skp/ijhOvxpDzDnMIRYdNnMqXA05dTIr9ApDGyoKv/KIPSGt737g3O91
lNodzHpICn1uiojpfm9M0borVxCgf4/RBXdyNIUGhrrl8nLPMFNeBS1eu8Guhb1W
TR4rbdviKuD4JnhDevvWdemQ5SYnSsqR+I3KLnMfNFBvUIISiE13ofrj5vyWjI2Y
yO+KoaVsdRsr4DUEBw3BG1aFWI1RxEOzR/wqaSwwTCQTf1To96pN5wSWwLLz3Mul
8mMzTFVdpxeYxAUVX7TbZEPhLf2rOV70vM485d8Cpvy1TFVbkKnkAeazG1UcHdUe
3Jqr/UrquZslgZaUvwHmGDNbrAmty/aZcqzgMeUEztjDuY3mVau1WXh5ReAjlqHl
y7iSeRCAjy1sbimgugYK7aStt//MI4a/v3o3MfritObTiiDGJEkvr9p8UobvBujR
KxA5JZFa7MCR/R5QZ0AZSs4LShn/CkoqTX4mvicPrNh9VfGuUS1627ZOaA1wSsJT
m9EnBYGmyk80YHa7qrq49tyGBSQ/qQNvU5nBp9ySlCTiaYgjtUUdVKxOnGRTl8QG
PiBJTqEErhrYI2NM/QDd4qlwBca3o4HZnPBQk5yTlkg2NIwEf+BJgEatWqa+Tn3B
6ywX9B3hKn8RbSZ4aHpp6oUn0nCDiQYfY1J1yq50G9+V5XVhmHPKxnfOqo4+Q0FU
xIljWZFwd3HL8JXoZFIw10FWaj1tl39jAO6MyA8k08+M8CsY39rOnn31zwPd7gLc
avjxcw54JtSHJhHoKIwbghpFUJzyuOaDPxBtzEiBYQTAiyLRaStz4Y2WL+F49zgS
YPsHEnE+c3FLkgDCGNrgYzxVWeAGH3PsUZkl5VlwSpKtjAvdBhD3UUJHNw6UwvUa
yD+plSwYOUawNw1xonRGNfmTxBO5pTArAmW3ny68oLMDceB47YmyBPO5NN6NxB9+
JrqP0vNDnAKvxY1I5BTHtzr8XurHba5dq8bgvU6LRWFCM+AKx+jhaR9iTM2anBbv
lrC7YQ8gO6A+DBSDKbZVIRnhmfa36ALMRza+f1+dUsseUk/aI6xiInm/cdmE2Z/e
hgc17PthDq7abL6I0Rw811FXaDEHg+vrC5joFVjeco8fzdPHX1Q1AXUnS/jJMcPD
WU7NJrX8kp3iuvnSfQ/2elQmBr4zHprEnD0+LpT3MG23pTjTV/yCbo1iP+XkmMkt
FTe7wonxAc8XpczsW6skUJq/OOPoaHVT6aWKB4AzX59voc2DJFtTTBeCumeWcJo+
9MxJAOe+L0BAM2fvU+e5BbLhhBQVrAk89pK/a9t0QdwccfJTQbdcXwj4ecV2I/Vp
fzXV6U0+RL9tFJToCfOUVDsBXAiDBNPnmhBhpUUN2e/2TQHSSidh1Qyk8zhlim64
fnlGQufJlnq+V3VM0PkSW/FM7k0Fz0KjxQjN9/hbtIdHFLmaaeTkGIYwWj2jKZOp
X3BgyIgikdWA13YTLSBkFuQyT1TBYhc6zNSYPC17lnDYcUg1PJiGi2mg1/icsVel
cvNW4F3QfDhPCoa5n8JwDILmvt6vaT9SaaHhdL+lsM9yNFCa1l7NTPcnvmJa83y6
4eoi35m0CdmO1ffft3f8gKpH6EQDMVcl5yxExW6FBuVkJWVL5PZQZyrTcmynA5t/
TxN9KM3ynkN0idkda007uA2cItLLfnZ244wiZZL70TCBr3ytTZEZrIyEc22VrndH
Yh42Bfew2S6T234NrXLlA+ox58+vpwhZ/i9bm6VFqmEbab+G6VuQqQ9WAAClNXAX
IoesBiObb0WA2dpqPhzOftcAHgnICIDp93BSwomURzNl1UsdzbwlB41t8Q5ck+hg
A+vd6up1m89Qumz+4DPPre2+OidbLH8/ywj2p5vuBQRwi1YbZoEezyaqGhXNhB/c
fdqXNmfQO/dJX9c+A+sN45e+uP60xNlXB+TPv069fReVIwODmF+FufOHBa2kh92V
m1a/V8J4Sjj62Uig5vG8LSwxa3Taixfy8y3pZRfEsVtXBB9EEgSDTnEgzIY4xapB
dsfo56lv4kIJhoAa7wVFwd/sAIJ7sQCEI4Coer0neFNFtzql5q9eDBr0GWu+wzRI
Xh90nFCTYXPJiq4ui24KTaze6bUI1Qt5Jb4xZ7KCqDytZu9NV4ROr9P1x4ptkPZQ
+SiTYdyEAvecyRY81gLoM8f1tmeh34XH+gjKQUK1QZcbKUxOli+fhLKGENubjT6z
G6xNhafw7RLOLlYyMrpXFQfslAUMU/VZWIBenUmrRreZ/xpPrY7oCcjmWTzzyWi1
bmPXg8SbTavda5/1yhObl3wkGmn2gsE43KLmWn5lp+A5e1hCVAdzNcGtGdoOoFu3
lKLQVt2GlxXlvEKIQgbpa1F723pQD8HEWSKWFy8sMvAF98/T27MJOa6ONtJJjqSN
wJBP8BxXlZ/Tg7uHBxcgi1OVMDW25GHjyYrn/b6vtXHQVt4+zjqKuB9MTYlCETGB
S4izge+cbuPa3GKbOBO3GPXFk8nV0nDpCKe34YJXAv03kQT/RrVQE5DDzJULbOmo
h5r6BXbNwZj1NoTeinageJZng9AvTWEaYdvU/ycBZtuwNxA4nApNHeDCUtEQ3U7A
52xP4srbmr2s0TJhpSio7t6OaIPCs8NBWAtj6AXC37k/IDUU3kmHbg7+U/vhO2aG
LB/1ejhChUMnU4IGHGAL0sdpbxQaXZPUDVKmVVaQ1hpKkVmJdOvs/NtlhdclAKpK
91LFNpyQRGF1piTursfqrKIUCamAGS61hd5PKSKa/xpvIGDQdowr2HeKOSBjE9Kb
+D92prdye+PYFzX788Lz5y0TgVVLTXAWYeO+OhU5zX8zT0IHa5jTFbQkSCIQgVHi
2EBJ0NpBoZOVq+kH77niv8puqMR58E9OKNL3WET6bPBBXS6ly306WYdsm9NOcxG5
J/H66Vhj6AUCBeQsU9XoZaQzvUP8Xfi8oUTaYvEolPWvvPMc4/oTuyehJT+nDhns
uLwgNOix941v50Oz2Nio8KjQqkCvsNI1ZWq36HiUIqVKeI2CUWdLzyV21NJw78Cv
wsOLyEKWSDjf8R0N1Itoala4xrmh8idNZw9XvzJR1z9L6fP98exA7p5CqFNu/Xsz
4BV/nqtomZW9C7/6n+Hpifhmd852OI8I/stpGWsQE/l6Ak0dLYYH/5MrBZcMy8jo
DTiPOxWl04Gq4d0xJMU2kDb0apaTTx8C2VHFb1SSrt5zXn7CPj2GU/SY923PifyZ
4tmQbVej81Grv4sBb/emnYCmnKgebDmLQm0kDdG/te2aYnfkw6B87HBxnVwT8VqP
7escHxytJJxDfQZhIDj9g9c91TyPIhStOxcUd/UTae/H0lhc3WoLApd5SjCvJruU
hUrI7C78GbzN3OdwRzKaIdYsbqaO3O+/lGJvvxAYNraR3pMpcfupRhdtEAVHQeV1
8ah1PQ487g+SWyJVlqCGT2+qB+n5XG309aEGk09c9pJ/E3VesYskRlwTmeKnu1zG
xQLiyeGl6HW8KNfQ1UGyyk1joxVAtvhbPM6NTGZFXYpFUMYEZC15nzjfQziyF+/a
AQDCO3g95xmVBdWsCpwmSvWo+I3bNVfODC98oKYupbXQhF0yncM4T5H7tuw2V8xw
gfDaHpUr648zRVXxJWyUKkMk4DpZpwjKnmmXq48tagwZNz1cBPbW6CFaF2O3doU4
5IMlHUZOXqj4cLi29IH0zl8xK2dpI1/NkkyEGIkl+UGnvBfQHsbGi+mw+psOT/VP
kZOEDhmw5tyjGb+ea+Pn6LRbfPVwgfMglFHokpZ47ihUjTC1uvUp0wmwGPAMcGVl
NmKSwSr0cP0oY/at2XLfZSvqihy51ZHt7dpvEKUpIQKPJoX7eXnlhdaMPcbYUYMs
QDXN6KCBvWCu6u3s6Ng7dk585S5HBezgrLOoe2fIvJd3Au8I0/kcGDrcTT7YlHty
+qoPiilPMSWskMRXfOmj/q+y0ekEKNNq5IPUjbVrQBDnaEj5cyp5r0HfH4vLi8VN
UGAVrQKKyjwqOYbOZxRSmIvPNoc2uK9hS1g8g6t+nDyGXd2kUH6qiicYtXNaP8mM
qtJDJOVD7gtG8T2caxcd2+jLahfqIQqo0k+lui7bRxS67KJuOZkTpT7BT8k4reJ3
93ygarxqN6YZqRL6A/z5zRpzJgOiQgz47qSFcVnYNaK1pVm0tcah8VZbkv3TetxL
UuPwc4nObtN9/Eg+JuzRICjZdj/IAiJCJc3ZyQ8zMWQJJ1FEvvd23CU6tfbEg7ik
jX7fhKB9rXt0KJtnOCUvvchAcexwsgre+UZT48ahKthBaJlHbpfaVuIpgJbUBhrm
k8M82RordjmuaHJBVdI7A9UH0k6azoql/HNpOTOYwnRoCXfH1JocJjw3qlQw0tm9
FayA/8plWZZsW/kfgsUFa+r/5dgVVlDc1Kr0Bnq/hejpvGhtoj91v4z7Y04sBl6f
YnsiXCmBsDVWYfFU/b0yc5VKxzbRTw4YSc0//s5dfToUdTgxLT5q4j3E/rZgBhNY
At3hLDDPgSwfLAFR+Ythit90OM7UG1XtVc9cV9qOxs+LbSJUwZQKx25nLQXZNjop
EjplFVy/PZaX3ugCesGPeaKg0AbmBrrZ0Ozo6JxODnjrUXBuVaP7OR7k87CtY1fK
4QyYAP1XSQNayA5m88ftvfYMouAFgsxFlbHvjjkEy2pZVPyGKVkoQxglaX75GJGK
r+pFuMu0S4AOk5N/yGcWyv3UOdVxgxP4EeGAusvDEolXPGvq//VoIu2Qs8X9HU5f
5vwsNed3dEu8n99j3mkgp1Sk4P1ZSg5NUIyoEfESCSGafh2jggU/0IE+erECWuq9
fi6jqqg0jScRIJ7jAlVHH8uH1jdwaOby0Hrjjl9SwKCY1pv1jdIQJUj5FTYFaTbA
oC5dGnLzqfE8lwiRLGp3OzX3OVferz4HuQ5gH50p1x1CJrmUbwdvxmttILN3NBcz
MD6/q9fFticOXE5Gkah1DfUEdinmrfq3+Z68srMKxqRgW2fyVPt7dmEbXZWyJdPn
8Ju7tgpcvET6VUo7VQk3gic6QAFHQYofdVcsYhagUa86WY8uxARFwitA9fbvKsNH
yeucyqFMDSOyDcxUc+HtmuTnIphgaE1oHAOQ1mczSUMOWSjHABtRiOtULX5yfRHm
tgC3lAq8W9cVXpC0UUXzCmN+B/k/uHUIUt3okG3pVwdrix8eVf+uxjNZzoW9WwqN
OmjkjJdia66j2A1aTBJCLhaRtXzeB+knyYWfQoyIYjNhXPZvfSufH2fKvlcco+EU
2v5MBs96yommVmoel8OlkzDbMi1tosnC8727qgTLz7MEU8sGYm9E20Fy40sdJsJP
pCwq39PEp43WhqfzTP2jhAMgb5Kf+QUBxE6/XiHqNkrIWn4sMsWOBMMkaBjOTRa0
Cf2bhkGTQYFyo+pYiLS1xSCQ4l8XOXfwNyPbmZOWNd/9JaJhB5TXS9JTXmBtWl9K
LwMFGMKvXWPqcCf9yI1zaJuh5feXGzs/9ISaM18AmPya9yYmgzkOZat54JKL18q2
k1vXpwbFYz7u8OTNaFW6J/W+cN51Ikngi5Qm4T9Wl+RuWLwW6SrTdHQk+rTOq2BS
Qh129cTHws/XLKV3bWUq3uQwnoE8hfZZk4hREXCFu0026Z+DlSjxCBIg4I73I0me
G9jN6G1PCNID2rvoT3iZlhJKnEQLsqqV4qZz2Meb8uJW8rovdKDSrlo8fvgdwvDT
YmpI0KJbTnI7z+mrfuehs8n2EjSxCi7N9BFe9c734oZv7fyCA815gvhjHLLjAF7h
TxbLJ2B0tA6mFiGoInvrJdxTkzcvP86jD/6hbGMKFZyIwHJWT+1XNWndFyNv5FzF
KuU+g5U8/458zCsPC5sRNS2TCBH+Uoshspf7U3jSBB/HTGfBgnN4ihc2t06be86W
agLITxgoIs6bfnD1r+7+Cbu7ET25OUe7Zu3ACkBwdcVXFOJY192jRlPeWdFH1NI/
wBlLELKFdveMO9I3wsb1LOWe0o94BXPcAaX7RluB8Zo8y6oc3bX1Ko+HC4xdLsqB
V/XS1T+Q3RSBblGFvNAH3dIunKejYCvrAj5nIBVia6G1UlDPTB7nSZDk8baoU1eu
ZiawbCVPdVuuC5lY1s4xsgjz2p/fB8F7pa8JlfUK+Siqy5au3BMkiPPrY7WFOP8j
CeEvjL201fXHH3VVsznmEaLzwVgbAX3HzDjoUIs6XP9B81DueKdu5via65umtuN1
PSGg4YMTwdVpGFXFVqLnBCgOCKaV1Z/ufc83nrbbx4d+KrUTJT+bsg8ePFhWn+rH
9tAQ6xfvHBxpj/9yL0SM+r0hO2RygEGOBetli+SmGcJmcih0mP1WlIfh8CM0ijIG
ph3HQ+ALwybETDQg/AJ3aUwskB1+ehj5nq0ZOLQuc2YyC2MJhNYrRIHQUWv/cxBI
GNfudWFMdsJO8n8qFAi7O57et8hBJ/4eODtG3r6hGc5l9h1bWN+j9T7BJt2dHdLZ
eOQw+pKfzSr1siY5fFPH418/yXOl+774WGWU5FJR64qDjjmJDvoCvjHLlnKUUk+2
9nUAdFFTWDM/AOKa4YBF2HO4EKCRU/5F39VjgNMEx0dGeaqpuBWgYXdSX4Snfozp
BIouIvp2C0If/Z8Yxo5RwFl86snkqqovCefwJgLEjRR9dyA8nZIAUOojxWUk8nIN
wZl45sUplZFimF3/egtJUudlyXoPUAzUXSCttMOze62inAA++kDy9ixitPEEIFp4
6o0CHRyus9kR/mqyiO0pGSMm3p5RXFICop5C4ayqxEjdhCa3bRIACMpvfW4LG42f
Bg4VMSkcNhzeBOiAeNcJdr9z+5X/bzo15bocxNuDIOClcpgzwsdl7Sed104/FsDA
dWLjQ9dnB/1+MxCK09njS/3q1o3twp4GEirjCWdP+ZOngCg8bW2eTeIVO15xqVZe
7Vgv5UczqHfSUSiqf+13e1vyql1dqUKbUynSBdnk0IZA08GIERIqj4y8hQSrTc+r
2EBUHMGS2aLntrfet4nZKUuJxERpr1YFEcjMWGLi3wF9CANHS6ksbwgBMI4zVRWH
7pOGZOsYGzGDTqRxMiDDXDUmAU6geprcN8DwohvXHqXUIRaZZPT0yaOVNQl17f7m
1O/ennthFgppNEwbtPi6uAXq4JFCCJ8TL8wFrfE5zrLsmU9CW805DU2tMGTnXL3S
y28ftnGkerZI4zo1XGtsX2X8bUgllVq7Dmc0vXEr+tQjGnm4LjfwjkTdsM9U+H7l
H7wUNxm8mTabdoi/T9sb/1eQBd7pqfaXi49sOI57cXtGjk3wU7tqT9FJCqVDAcv0
fprw4LdL+f0ZMVSp5l2rEPl/vGwbWNcWoMt9sNaKv2JnSTGWkibxjVLeMoUPv0yK
yFB8V/+yU36BAwKsUssKPP+1C0FMpJv3+zpXEwktRVjFFbzhBO6nj522+xb7bTwU
8tvPmiVxxI8sSFqGsyFDvkJqFxC3iHGm2CU+wBHPYPrB/sd6mm5SHseAOdlGPFiB
bYVH2Hvt654Z1bibBoAyIQM33lUCJ4y4ov+2GZ1srJHsL5frLWzPXGQvX3uG0AZn
1UYeYMcFfEXxN6ykIjVqUUcBvuMpeoQKBymexSNVYRQo0pY1yf01sywPaT333Ngf
+xgoqUVrWJy8BJ7xWJtD0Sficr9rHynIABTGNJ9V3+UCgTr/ywjOEuKQOB9XE1BP
Aay+E2qrmNzkKiN8cTTXkVIG7OuRtcsp4lm5qKXqCiGkWapUwrVww1XvseF428iv
hr218Xq9oSfCbNXkinSKumqJWK8MUUXsH9WQ6nEPBpiaPJW8yzJX9hdtluVSH/ca
g1n3msOk6nZPD1osLIvJlwTgrGlP7Ib8Uz5ArH5Z/Ql2cO3Sjz6xPHSEym77Zm2R
ALTUubjVBlxzF9PfAoayfgwgkhOzGwRTL74y62yfVMiuQ1LbaFnUZJlp94lpNrvq
CsXVu3+gxqglj3UeJhKAVyaFUh1U9VMe6pMk6FrHcSWimhpPV9TU9zee0U1gH4Kc
kgIOsIPto1Q19ajxCqtNk83KRKsVMPd/CjMrq2dtygUBi5pI+3sOEnClSR6hkbKJ
68FOtcaX4U1vLHYbaYbyL/bBheamPj1hlb6J1K+92PdZJutFI/hcyhxiyjLOv7LW
tl8aCvZYfl7qLpi3hPmwb0ir4v4Z8HgWt3+zUxgw4mDzYNXU4JOKX8tBs7UYbAV1
I4dPIM6Xk/wLvoB0B2ZZlt4lfepzM+PrMRgkXRn62LDmoL/nEKjHA0fW8xaW59JI
abZJSZsDuVR2mqAtlUkN0GZNo6eDaIAQ7HeQ0Xewizjt0X4QAF4tajOa8ZSp0GH/
5zrPnE/LklSIYrV6Z41aTymVAgDThuIZpCuYGE+vloPvK6ZDDrelMRNhZAdvPClp
VIbG7Jc4jye83w916qTcvF/4CQhQdZfgdo7oPP++BdMDHcvTjNoLHgoBbrfxEwhh
81CafehvoUyesxwTBrD9sz9hO0+3roy+hgsz/m4JE1lE4x/CZFdZya2C3yigC1FY
koOXo9GdX4/i9dWPg3TXHpkRuZS9oDEm7nIfXgTV18MdhSKrgVWJjREglHH58hmX
UM6Bi6MKlMfzgH2Sf3eeUVjSwXBeWoPmUmdVzlbPz99bQfXCsYdoogvjeSKPkhO7
YBl7NKx2NnYw/nOEJPj6wJIxzGoeVJtHDq8SzqLUT0WGo+5PgMfaJbNlguUZGm66
MxwD1syHsG7JNJIvhlAkPxvduoLu98ciuWoZL6T/8IZMjwSwmjA/JMkRirDxQj6S
etQ9PyMomVskSY36xXGe06V5bJPwpVMjVmZwNnjXeJPh2WDipkpRIGsbuF6tQp2l
+4PX0yhNKf1/HaI/4Ab5DXr1Jwg6L9/YxnJ4rQ6sJN5xveXFh89ArmSdEd1QKgHv
Wx4aMnq+i+fNIFtUjBxvyry5jcHJauq0NtzrXNpZCnbIgYktNHF0YZt4hFxlFgWt
A/ohzztNC+FMNlpapM6y1YvWAZ2syG+BhoRqC2LrTtURVRk5Vzk2J/yEy25wd30R
kD9hTfGgUhEM+7IU6CPuDEjtKvhgS0dj9ANCSbpgq9EnKQvcQDDkbO3bxwlWDdyz
fIsUXdU2JWRz+xdV8uCmX056ch9n7HQ4TH8f/oRv23dnuy5tOosp4sTNU6FcnmYu
E8MLZXCRC3utHK5qKc/la+EdL2Qpg4rh9r0vUWceIU0zOh8lWDUc4m6dkZv8HA6I
nJKOBDRDCmz8vW+rh03MeA+X0hcDFNlmqyAfYcUyMBxl3Ry1nuexHoSl+rZACR+K
mVnHPpN7yvIFdx4BZVEbv9677p+EJePLXVzKjwv4WjuF2OnIgDrxgArof/TS7XoX
mPHUKQhFZ0Qzrdk0gOmEbrxH3amfP/+RwwG9gnjYjiKPM/hevszMGPdoMK+W3Ha2
K8woPC0NKDPAj6dmg6w0mhEZxNK6L3+3rMiGha7nVr3zGk2qWfpUWMnc2ZJTpt7f
L2eHrVdmKAm2o9LjB/eZkrCSNMx0RtLD5ZqQMAqFv5/ezQ9O64sEy3SXFPIwQZCm
Kiu9Ua+fOIEkPTBIXtO/VFYane8QVJ7P1BSuag/PTws6ybEzC4FgtlSx3+KfeYER
PeEPPnp/NI3Heaxcj8IvSlUuzF0LegcTeG74ut7WC0CHyviHm0Y/vVid3e5TLZEp
fs6VSTA4/3Agx4PHTjjlg5efrvMuBKqQ7kEQ+YvX1TVyPUqRVNbhZSgpxw+m9fIl
7ytwtB5iVt5w5jpnDDEJh4fkr2H38OeWMVy5VtYTK4BvT7Un96hMhXbSAmE9x5Qf
j28qWlQWtO5WC53aKyLBfvTxieEIKbIVdVPn3Anrkc+ltOwQHFxvZ1n8KkI9Vmjb
m4g9MuOWqbgdvhMnbrHOazPqKx7lNiv8sZWgKm6n7IJd9QcZu53qhxgY0ApcCPBy
bYyjB6ErXZiurgEmXrAY+axtL0/e12BjfmJLZxtx0Lzwol/XIrNh4P4gAhoD/PKU
IdXu3zRSUeFOQqDeQ5TLc6Xs8poGrnlWmlnv+4G5FpLNa0g7j84ozPPqtT/GIYgQ
dVaLdsFogPCEpkFcEiJwCPo2vDN6H1N5PYzRh6FkbxFDpmccwukRBETNyTYzMhuI
dl4nZ9hKo/QFu5Q0wLphOmm640Srfw5H7XHkVTKeNlqkpeJ8NOQxG9rQW3QGQWKe
bpnv1L95di3LD/A2eUCyEw/Ulr4zHv0oe0UUBBvOWXJra8ZPDVZzbs6VxpxseL43
5iZWB83hR6GW/sys0u9w+r22+w9c+8Cxu7yezfaZ+MQCRjTAIHUNlv8vbmaQozHu
nM455c0x5l9fwXlXGqo6N7yiPJLt7N0J16muySdaLxEfrjtKnqURRrqCOujlOane
rRFo5XnXwA+BqYCDLoEPwd5btgQ+cmQU4pr8t0A2lSMUu967d+oW0Lnk1YsR159L
Fszs22y5ofE83ia1oV8/Q6ETh4bcwGcw9TQ98IXxoEkAbNwo+X+ZIHGxpMvvuWWP
GAvntksrav+1eoG49diH8KQLFphPBwTppSZkccuRS7TxMFn6nD4mC3GRGlqlc74r
7kxf90RAY79G5T2PRHKhLcl8d/df/XIX5DqiwNwDJJtG+8zO6dygyXo3BJBBkT8w
QW9X4w3JoQeJ/YOniGP5YWw5p0wewjzRWXO05R7ABQsOnQmn/Fl1NbLZTOQygjWL
cNUURf0KJXWquN90YiyfPg8xb10vh7w1xLRFd60ZPkw8vAzKssmOmL359b/QjlW+
0TyyZo6A92IxryVmyIo8DYpON6MWAAEaR5kwbWMIV8vzoaFlXxiHXCyChAUECL4P
X1OO/OxGxe66V63sbyxhJqJZqefMk+fmDa0n/DSEqVcM+GxnvDOtf4gaSrtwxzeE
bj6CHJykAkz5ByXZqFJ4clSdFdjRQKh2VAF/QU2RVECx9LVnYviYgzPtgQNZHI/Y
xj7HXXXV1PQQ4fe87zmee/Eg4gaHuckyopcvsxZ2U3/XYwESvHYs7nU2Yq0zuwGL
0iFbTPMnVQLnBnCVqk6uNSKfLDDwgOAaGxL0KWKyJ3WZM1E9vf9KBRBgahmUNqMS
332L3Djoj6APLIYA21xPbzMoQNTVP3MxBQdJsG9MdRhgZt5TbSzZJgQfGXUkCHoH
GK3PSNc4rxTkCL+XFAARptYZb+P0h3qkBCzjEFomC99rB2PRZfann9idgt3BsnSQ
7C1ImzUPDWD8sCjginmrVV7LiGD6q3nY0TM6K7/DCgvscqV8gtrz+2az1+q2ebFE
O7jaVolmCvQJRL7jhxGM492Wshvq0B+DwlhWnpEbA0l5tHQvhXr6G7b6ODewUCiK
b4hqG6eySrHstKKPxc2lwAPq8jWiJBWXazkUsOqcRKmR0yKMopZDGE7FKwecRePi
eaGxPjIDVW+ML62AhXGCkqxK2DZD8x263xBKBqW53t47b5Uhg15NPWGIyZZlnUdj
b47jFBbBsaUQqJJOUSpzFcdo0i2RRq/XaIIY5+XslpT+q7h8H87IEp4q0/4XuIBw
IZAJBG3o0dj8OGObPjmEf4AzzY9DikajHJ5vD1qWmod6+buAk6ShmTZ9Kef0iS8Z
fVUSQ5SQQtlxi9qs2CoDdhA8uunGOiid+QRLE9sNQPCThhAOb59t6qCgrizWBm0p
L77/6EPcshPv6DvT2CSl18hDVO0/xQrdlPzwZjfimiLA9pEE1ZbAsso/TQt4A0zx
lSSaqRXfaqQDCx/S8W4/TyyyO+xWjjD9rHGBocCy13YbmK3FrUZj00q5YX3isWst
WSSeYBLpaWGTFUnHzKt15LCyqR897//Na2g7woIn8ondXQLnCxcSua4dDqXwbM2o
kZLTJqRIr/Qp3Xu2hcsYGdmg1GE91wWvB49wI6Sv34GihC+JOUJPADZMoiq9KAW1
PFFPfKK0aC58IHeEm5wsuJKSHD6UFttfwT/LuF6En6R+wgDbnS0hUvyOImMFLrJ1
bb3BQyNl+q9YoNWy1Df4jtSx17Onuvbv8W08LnNBP0GIKzLEirGPWxsLNZFIJt3x
ScVYZg8/txojAZBdWC9X20McfaxOl2sKzG7zxRS9KmbFfZI1qPRGchNfNgx2HigR
dKXiapi6K417FouZsIeD2ltLP/mva1FCTdvJWW4Lrc3zV0xU3WcNz2gc7hNCtn1j
4Wh/arvcUYRUTBX3hU7XzJnJqoCDWefKCa7+llL63IUmRz4h4XRFiIs//WLQV4xm
gl6DYfFKFt/QrIOm4XcKpUIOB83WHEFyqXzsM5R7Rwg6KRMx/R72aO2cy7XqU/wT
KVGQlyu9CBQtMYjm6nOaQ4Ui1byJ/l8P/bmXomcfqO1uTPV6yPmMYa1zrT9pRaz3
j0sGW9Gfju0IjdZJELkcX9jt6ArYxUYnSV4v+qnu0CDp834ZckKLSSygG4vDaL6H
yItrLQe4srXbXKJCp956oL3y857ohdsxuwkGwA+DtO4zsbuNIDAwKyX5ItZrAQ5m
RZIYglHsJt3Bbn46Fld6xMaMOxhIAzjb4ivs9UTRFDWsqtUpnlL21EemncifcroS
6IzPoxM9/Azpmsw1yJdR/UarsCgdP/Z3ddkvV036V7uzZJRnMZdXBFtweqYzb6FW
N5Dnl5WLwFc/Hsw6/FknyRAdJlXIUANTNeo9DIPwOQd38Y6BS3vHwmWWHA2u2Onb
eTMAew2D1aDvNyXjUrI3UIhLWt0gOJrlvgUZaeRGPYb+KOkjZqrdxaGbtgTZ/BMu
qkyGPq57UwjvqJZeLdKIpFBU+HjCqSWjeO+qiJBE4Al73Vj+3eFGFqyK7pSxxCmy
rnU7WBFzyJDvRKc3l9sR5pTW0XN9FWinSZ2Xr+SE8L+aCNV9FRD2KCpaeiI6SDgW
B3cR7UU4KSnBpDtG4KQGF3XUSHvyTHQ6Uf0GLWvmpYBikt0WmIwXb+ENOfKmQULE
vqXt067zi5wxmBBngD2zoYHTftu8s7vziP6UgQE4ANRO6gGJhJ28JO7twcV9/AZR
FcObWYSO+tVCIsgCNQIv7KaBZAm4g5ks2iYjB6ybYoj0rB2E0JyepNOwZJFzsffS
rmKApaKqP5uS0fsFkSmJeCHTo9kSwhNWbLDhvcXnUacB00IFnJ9lHKEobIkDfL0Z
jRM4bM4O4xXSVOD7Dmbu7vr/VWysVwuI6BmHF3cdEdf9ONpX859Du38gQwMObAnb
cu0/08giaqsDN75lr8b9oKUxS/wxeNx4j4XT83fwsCod9tbhwZbn7jC5Jh+IdTF2
PZNmgk0kj06FUoDRKdxnevdITArEMHzEhKWHzptZMWUF9+BOPvOhvPfpztEM+ll1
9n2TAV3sOWmEuDuSU70hfCR3jff6DPvu4yvpiiIJc+bW4Ryx8GD5MMLpBLDDIa/7
7Bh78Sn2zWJQ3pvQQDpt63OOs6WN9Ym7mf0r8PJhs4wzAh4h6oRntdPIF7a4fuSO
4/DozXwC0/IdKuZt+BgzminPKthyCPPPUvTcB4w09iou320F+5oT0AgebZG51ucp
akXbSweYSLzN0WAXoUOT3vTqc52jX/6t7SrMdIN9VF3x0GRAD4S1yNMP8pfJqEyf
e74t1k1hGosOK7iZhxXnYWWvnapcp7t4RC8zSNC4pRHauGJfA6MFS1qBoT4rcMpO
4B973k63y3vrkmkuoYUz2x23XkRPIwD10w28rWLMjO/63taxgmU81apfx4k47Y9m
E5qvJVp+TboSDlJ/rKE5gDYP5HtZY5geblos++U+mbgz4dGRu1JqJUR1zYS7MaA7
iZ/e1feQKGc6S01srpV9zWpqrVGRC/9pxNF/pABCBmp6etjI0xxkKeUa7NXFVZpm
hCQf3rpYhFMhyw3GXVIPnTb/FIZQOCopPVPEtiAUYu6G0IK5vvyjjYLLB6Oj/mHl
Ct8sCn5U917vvwKd0RFL3K9/J5coeeLiOI4bkiILKPII6Fhy9JVf+IQWtDUlVg6E
AAVN5x+PhZaner7d6RmbSTbowDau35KuNqfqw5Bmd+T/j3sGunU1/fknDTajxRs9
txJYl3DlQAzY6TOuJuAgu/yyRiPYym9OMzLJWtSBZD1rINaWZGeFVgjM7H3Ez3kD
axtxUR7oFT40M5cTmHEUJQ414p3BhyZXm435nTXv7avJWjJYYhmxXdK/+UHSXoBT
ZeQv/ICMIEfGg8qUId13PsiOHJpuZb8UYB3a5pkB4RoT88HkXyk+8DGJOGV+4EaX
onBiBIZKsMNVRaIug1agF+iV8i03z520cZWvgYuBQKlq86qwCuQxLlnQLr+MP0IF
hLKMbI0LSNdQrvntgo5jZJ9GFGzy6jqKcqvHiLmjVd0XSXQTDW4Z1apExsNDuVu+
P9HzPFK2odiarg7oLA+rNHeMjDjhOy222HkTd6R5KxOFo9yy1jl8lIDN3Uv6aEEd
NPKYbiY3xtAS220CoqwdMCsTyQH5tH60PfiLVIfyddE/ntaeVbjjCEkU9qAIY1IB
urt3GQ1EJoUg9A4gHKZ/luXe4zRI1uZJq4C06NZG7FTvZP2hLfOPcYSjrdU8Qus0
jp+Q01NQIVikD/qt7kruft3hMIDMLNyJYMx9emPst4soxBqf7CRwprdETP6qtism
jL0PrF/DxCEUtKJo1hyZBM9Ubq4Yh+c3jd9I3biYrfBz18Qi8xJiK1/P5XM5/9dx
jS2uBzWqjvATmc7KrrKki2fmwkrCRM2dtFIM9rpHKgwv7YWS8VOdqMEKW3RPZv1q
lnyG21Rws6NgcnyY0q0wC88diaC1URsFaQkxZIGVG/M8e9yHDzvPs6ZHcilCWwj0
Ho3zDJ//dfZtsexkg2Xe3Tv5UpN1LLOGcTJ5tPd0r3iXalXMo87XP+x+3YKgIjTT
cJmmtTpODEQyLHcK7w0IdO75Ql94WMANiwOxcSdb9QoKVznPfMn0dAgfidV8oLKu
kZ3Vli2I/UOtkJH5mSpN41uO0dfGZGryWUS8dbXkf6h62Pc3Svejydjp91V/JD92
q8opVLEQAQO5oUDzA+CVS7LuWaWbL6cF9im9sfAs7V5COen66iGok4zpOQov5dl4
/QkReFG52H7+EjhiOjOQxyyUEX3hHFUMGaY5K33tqlqk83DEtD4gK4VsI4wZYTLz
qKGm/tLFQilOEGdetw2ISDMoPkd27k1CMQJcKCC5DfpiDPsJQcAX3bjdu4xXQCRq
Tew5TipcGZXpHaDDDlVZ9n7JMNzm9efJw81YcRB67rglzsCNOeL2MALwafzDofey
wNPLtQY9IRM+xRz7nMlggNBm9bsUhv+a5cHGQmOmTZWNgRReqzE8jwvX+wxWJ+Ef
v02kDMM81pGF4LnaJH6c6r700ztb+JW5gmYRRWucGst+qOD6ydMQlo7O1QmfQh7k
ORHa5Mgloesl12JaVWbA8dhIs+9PWrzKEPg0hyhdSKQeOxYX8W83LuzbaZB7i5i8
FM8uXROXqleupchkD60WzkAo0wRHGmhgoF8cBs3KcGpEUr9j0BgPXdeecXo6LyPN
kZ2iYhf59tgT9oEoG3V/9zV60rid86LTN5HyH783Yraaf+fLLWpZfDXCkDOJgTz0
J9GcAAw5YviCgMMoIjGUiJtjDK1B9cnYqQDdZdzMGY3zxgjPAfRGjosJgyJLp//N
UHbFMHCHAIBwjYKw/hW2P1BZee++xVoAo0aYMUfi1lxrNMWCXe8pXu86JPhnb6xz
yhlVwheR6BJhJMfiO8i5rLcPb99wu2FkcHVqpva/JUgKx5Gyzai62b33QcN8Y2Gb
cRIec49KB9IISsh20DzEtVUK0WU5XaVIA6oQfLl0iZ3+rd96mu9UUQWvVsa6BIld
cq3QwwwuotaYmhtJfe31dfjhPOJ/IDOrcAJESjLGBaD4pawTx2yZt67vZZEWgstR
xFk6h0AQFtbpoE/HuRmEv8fMvS9GWmFckhorDokKKvdEsc6R5NXhG5sqJnJeKQDt
tONqwNNIrEq26UTY6Pd+qakCR5o0ui7CMvUvtLsGRQomwQDNa+1/KnPRqL9vF+SP
xqN181xb5pu7ltTQH0Yt7uZGnxhu7ruFXtkSbo9RHPwfep6HvgGJvPjGyCv8yFOZ
haEsH/xcIfsLe+dk/2Szck6nri1xAOUwdeRysP3UH34UHg56IYQhGuCXD7u0KFjI
wbLmL1g3znGlQF6MLC9gBG+GXAYl14exi7xUYPSe4tpBirY02+nVeH/ebYKMGreX
GWcgpDFmuyjH4c9xup6KBnHoDTn0/gC2knQv9ZwyBDWDMcP+PmnRthKRAHGoVr2e
Up8k73aRSXA7hpvLc/ULtziNENvAiPctVX68yGl5b0/r7kCm0n2jvPtz1B10vAIi
uZtoSapgIa5BkAlbo/n4kVtOKJC+DuRax6SKiXbUI69OkskMnwj03b+pr5iivxjp
vEuYRbyaof0AYzX2OfLy7sXiWSOj1+02rc7Djs3V/ajdz4b6PcXiTH+Y/5t4WFg7
+Gs2RO35KXAY2EBBEStpuHHIdAxP1/kJABGKdoEfJMd5jet0vzgxq2x3UgWwMRIi
3DWEbgSIbolY1DEOP5Q/TOIfUYCjAXgo97N0rMAc1yEPshesgOWBXKqVAUfE3bfl
BWE5rTPdmDpg+uMcgAl5OinJsh5gjK5+WlDJNOMU3SW9YWvx09pzZiUtE3ic8ZRX
8sq761AXYx8wRQCMY8GDCF8z2ZbotWpvPk2tuHQx+4RNmpmWwgLXHHRf4Q/udyAI
Ohkn9fRTYEXAH54Ts+UkxAPgp74mebMefr+uniLpcoVsoZBjYpMaDNR/3F6md7K9
PDP6BTzoqNGgBlW6TPsDpXQL5+meK8WKPu9bBhX/h1GiSx0KT03LwS2irfH7D4yK
Fag3k7VmVAk77MzgtrNhNQ5EDFEu0kdA/n8NXJQXcDruqkv+El63PjCcL/DlIchn
WpQ9AIZuR8de4LxYVcOc2AMGfxus33UNXr0IyvRxGO+l7HwFbtKZUW+kLymhRbvv
BejENBfy5JWAPyDaJuRKuWxsZhPJvXP4hNXVK5oOIzC3++O3LoUV2pSy70gaIpUI
gxClT0sMPBnz+A+Cwj4iIirXkzkroDq9zgpdyRtJS8+4QVs8q6wFnsCvhILnR8+s
Z8JPdyBsXMnbo+w5It9FfxUgLhNzY8rbgEL1BSadQAoi20LK6cuOW9ewcP9bV0Ul
qCR9Am53dwAtc+jZn9mU8UHxra5IbvPwvTaiJNLUaE0a8iBbPw4JGwbaH2v7yTpV
ihfhuxx9mHvsdE6GLkhtGjAX7bmxFEfTDT/8d7G7Qmec2onL7o6+Fw9C+t3595WJ
pcLTQptb88TpEOCrNrMVvcsg7xT3q2vBRGEIabBOWpdaou22rDmrv9Qqu0a8mtC+
zgAJb+IgOKjj5VJosEviXAAv5lTE/HDR8iZSmyqN996yOzrvmDMnn54NGCfmVv/M
uwLk5nTnWHPgM5EsPkEEKWdBvC5XECjEBJq1iGUemrSQ5qvFczsRDeTHty+ePPGK
UJVg3dCyCmTWNqSxIOtc8UlQBrT4Q5nSMsFX+Hog0cREXt7/AYVkjbCoK4t3H3lD
DfP8iz1Q/kB77RG0PMmZlLAaYW/VWpGQZnKl5PXGFMXbzyDOk7zuYQAUYh7gAsZq
P5CWFXM3ioj8gzEUFJ7jO7TB7mlOmIWLdkVTT9uDghPIrWiz+GCsdV2zPhkRFxfD
S7093cH7dS6nF1q/940ymRr5RmBGBsqNi6snUxhZfDVIgeu30COdIQgaTDkrcFaj
MZyJkPGJRgyd01EGgxRSkqSkpJYTT60ifIq1oNx+lBvkNwCmsTBvcgqZONJqgjGv
R5tC2wtnhqIB/Yh5/GA8/JkGF2EmmRsp0CerOBKw9uBBtFy/21D78GpLZSAzG39Y
miqhOTM7Q2m8dn/vd/HxVhm3DJrCGbhzG+VWC54vpwtprZ3jRKro1FstlxDUb2Uz
EwkpBF5KVn2Lf0hmCpUzFp7wYsiQJDZrj2Gl6skb2KdIKeWPrfoLRGL6U2rLsScW
sZ10l7FJkqhCyJgLA4tnAKh757RfLEBdsneK2FCnNPK3+/z2liKugCDJlHyXvvei
kvM2Fq38qs29rDiCeiRWrBIPCBZfZoA8xc0JPN6hxa15QG2UkmTpZH7dcjIHPjdI
5H5rzKGFDq9mq3B4wUwl6Az33EebsurN3E/28NCaoatKub+p3LmlVpZ2qKlReJv6
I6RDeW6Uc3BshDAv4B1TCS1Ke2HliyiHHqADPoGhehr1wZdCNCv5QqZyAXRC0nE0
HVfWrhlLKngdRvesb4twu0gNGUMyEFzpvM2Eoux4WZmhNtrOErzc1D8UvEf9ySsr
DJsa78ESQL4NUVVEU6UBF6ZgBydysxgnowK1sMJiFyOWVbBEV6bGSExJmGLayO3m
GEXj1c4OnRZPVqjejtJBJWfz/u1cGmmzIpYTplJIUHVzaIQJLh0OoXkQc/37fPD7
v0cu9pJJWAqHpsCJjCsg1p4W8WrPEmHGYbMewxnh8qIaNSrMnPKkqxB8wwnqKhLb
HUBZiKiMvpZGL8UYTk4Z2AofQ9E7wgj0JYDGqYYl4s0SkFSZbcihAG5VwI4DizV3
MpoXHIwkzIDlB9rxj/sG1uTCjDqVmlxgn+C09WgrbjI96OCWbeFUETcOp2R7fvq7
8lLyx79Q5sIq8/oUhkf4llcjDjmmLDYVMnEw4i8pocdalgfD0HypbRyDV025+WHd
bJ052qbtnwJKZyK66sJXU5mfHigVdnH6DS+2qywTfK6hapsLyqWTZ0J9bB7z+eUl
IloiTkLdbJt6AJVzsgw3G04uodpIuqbaJO2dyEv5GZI7tTdICCf2YrUK+1MR6vcw
b/tpiqvGeT6GWrgInaAUs6diueL4iosidMDhG+jRwimNX4NfezkMOa2GGifNItCD
PackHPZzCfz75OmXIs/xwvzrXf7s17UFOVOWOZ0c5YLaNoZGS9X+dViIwj8rPcEo
GlL/9jCGbWpq1qqGVr0UbLS8tF+bf/mkEvRtbPqnGqTuA/EUfpkrzLGFBI2yujYk
nnUsnPS7a9z9kESbUgTQ0wjpYG+DOnKGo7o6X+JR8pBnQ0t9jxz6WuB2GMt5+sUd
LQK9rFgzAvmdMoIMVoiZx5/Hf7wiGH9syZxAnoESp00uCXco3cw9w90xHoI9GoiL
ErtieBKY+S39hg+cGpcVfoUN4g4Uc4SFPnqD62MWenzjY1PskxDBb4ZCQLICZV9v
NJkFf+qhNfBaA9uWSEFq3WoabokukCn4w0Ph0VACAIoS4iFoDjcpWCnbLWMP4MFk
T/fKZENGnrwZVm9AadqQiIrDiB2567n1IC1ZEw0YMCduUZY3b7+U/HZdkEi/pdy4
ExptjrAf80PcNJRtbBrQE5MEMMHUBhQLDQjwt0iP/rZtggo5ypk9SqCycZZevWP0
B+L06rLXCRwkN9jkmRQCzzGaLqShjfjYcZadHTgy2ZeS1glH0g8c3aFcd6VfCn6A
QjovxJdVfmdJI1XL8JeeqJ0D7Dx2op34KTeRTMgyoZiEXVrr1QJzXrVAWQBMLJ2p
EDFKiuMSIZg5jTjeE+kbl8u0WxuzbtmBDz7QzM16CkzIFMzZlXtLblHk+ImutRVQ
PmJfWVObFrcaROf+vqJHCjAyoAbU1IHg6OzZgHbps97o2vnGh6f7GuJXewS2TgW9
7+QY2mvS94w8AnWdkGIYzi0h0lD+6xRJEk/69oN8SQAW/bpeG5Gk7I4nPr5hJVSD
zCeHtY08FvMN8su6hNgN87Y0vQBls/bly+ajZHZ4dZYr4NqNMz4Xn+S1pYa+UsYz
FRZJDCwdkwGqIZz9j39WLZz2JFXCiTQzbUl6wCkp4SXVjQLF4qaai+N6PIR8SNQC
m2UXAm6O9j3guMLytgZes5cfOp5uT4XIVAXvVwKgeFx7LICO+ef81QH3o6YzKXLG
a6g+wL5S2BXXQYY8rcPSX7BMu54QLeMVMlX/eB20q2XkjnpQlcOXXS2MQY1myc2t
szuA3j0NOADz8TTsxSbceaNrjY0Mhc8lk/9NRvbfVX8fW+emipHptNtDWqmQxZah
0FVQ2bU9fA3MKPZ8PLDQyipcBf6p++1C/ZZ90aVFH2WjZ/ASgfN4vmAGByKPZ3ZA
U+sr+8mGrQJtM0Mh3x5um6NMWT/JiyGu15fapWisQ/p1cdsf9nIpu/9UxZB6Mz2l
9R7+au9ZPa2IhsW6+TUYoOOgO9PIBJMhfyjrvugMs5CCEo+XCIbGT2ODLfBToalo
BdAv9VLCditvL+KN00ptR0oGWzENMfnJVhN3r4eOADFluYkorkmFyZrN+9dNFEwq
MNdRntcl/IxNqDLnZWPqjPVl5MKDYdQRvgT0suqq2UDCL+uCgnr7n7018b8uD9nz
wSmLNjnI5MJ7O8BLMcDIMj/ZEJBdgAL3gN3B26w7Rsb0I2v/E18p2I0hfn1ASfed
N7XQ0NMtzqL6PYbdripuYhkmK/Im00geTSkTXjG2IV8FtUq00Z10BsFdYyDCzmms
iNZ75nnrnoCs02PSmoVH5xOKFdBaDcGbGrmRvTW2znxEw9fcPphdsrhDkAozAdTC
bkaS5cn3HsFDGQCK/Zv8nRoOy1ceNH+qV7YU6yuQ1WdUEHcSXHNbO4d/FV45Pbn7
RGKrN7HU/ydeRRTLXLs8NQaVux3XfrMlMXl+TE4/lRGS1GXwcmKtmKhIfT3gOFQ1
fkxT9jIGtoGNTutV3phRNsA9mTrH3wY6thR+RFoyyJgHSVo3J8vkNjomygvm7GKl
+gcBMmclyAbRW6rO3ynyxQrjCfEaC+7VMZzX6uD1ls3lUlKYuRvQ556Z0s0C5A8O
CtJfaq+YSYmqVogg0iIDIpAP3v50AfPUPELnbX63w168pa+xHbpFCMbDT2HcQ15v
7CKOgZmOzEHfzCLGfioPLb4MPrpMd3XIWuG/FDsDDUVkV2VMW1mgxvV++MWH905z
qaK6EfiDzYxtL2kN+7xM9ERFDhDwf8oadngsQGm0Yo7MUCavWXRK55xlMiBIuPjX
RdJH7C1JiV7XjIj/ex6sXoOqdYHywp5htPInzfufdWgYCBriPgO+96z/Lj9OA2vz
KaXcLTkE/2kAoxdJ62/d0elz/c7tiibfEPvRlzb3AySVeY1AjkXIWyUEZwzTVT/9
i9RD4viXj7agWHkUKGSOQgzHqHKFwzCP7Cx8reGwWG+2OjCCRItkslatsRTRDAj8
SV6Q5t9Mlyg2s4gJ1beDpgKTmRv/Ew0pJZkhy9SaubUipWZBZQxj9tsA7PhzoluN
PnTWHbxuT56dP0/OOJNmVn4LfmlW0L9EE8biK1I4lwYgg8Ao96yWTNdi9NFzCUEn
YQoEYYJDGky7H/ormTurdcv/yF+h4CycC6V4Y9U/6FAby9WE+Xt8FNT+e7m5zXEe
dSTZuXhuJ1hmhE7jQEQUgN+/APhauLbnkIlLOQF1lNOWgatquTgLsnSINli+FO4S
InVjmb95S5CclfFPc7ZmM/QPXUy9v32aAGkumquhHI/sstlgTQVRflFX70/vAb3N
L8engiJ7UJ+RXyXal6jE964dunyYDVs2Q+nZf6WVPET9UH3HLKIw8G3yGuB8V8ut
L7fBBPgmOlSAMEQOcK75NuoqtcyE+9/HwlNtUFJ8MUUx+WKIAAkzb41ZLTdv/+PS
SAhnWvx5YeAsYTBFM9R1OT8TvD1dv+lJdApP2yiuMXgLZv8x/PnbygG0TsUFIjVy
qpKn1gBNk8lai5CTstsxtBPP5tgc7czUKgSeN8bHS1KhHH5eDSfsZxu/qlBPsWr8
Kd53zCh5cRyJZlDshlzY7SVI50u25MtdJIzatsO6uLMz3OkWppZ4WGCXoDuOC5jm
sbkMW7zpzD7o4Ooe6XbMN8IdoD9U1BZR47Ii9UFcYfh2LAshh8Gih2zXgD5fsgpY
URsrxk/BOGe284dmpZRo1qvmLMNFfC5fvInX9cUf/vycNpT0NE6EFjphKO0yAqa6
vVEECOFSG1CuPT5YXEp/fYSeXQ3Qo0Ek/a1gyjtlP+BiLKMrsqT1f46ZTUbwZ+VJ
tWhrmJhmS3uPG5HHm+fDA2u1eYsHjE2dFeR7VknEUl8/pRKEV7QYbMhKmWjSGDh3
mhyRtczonJjFX3vKbpeuUg/4aTvmIC7ps9FsTyZDldERnGvg5R8as+N3MKpcKOnS
h1c0nGEqBpXrSNIrUkLI7pNRYQhc8DPZ13TnbwxGBdoQnYxq6DQZLhFHFLlM5ddl
/RJCP0lgBbNehAt4BAEraqMuhnehkT1ZNv4m7PJ1fZIvw6nwCu0ZSzroM2RWSh5S
4XOQU5qM/yRS7mhd4Jlt9utrcwXLmtY57mnAmNP6SBz8NdRKhPZ4ap3Q9wI1lIX4
34zSECpWfaND78Q9c5nzI8gcZpqUgfbQL67m9zygZIaAAJx/M7XITMwY2dI4WD/N
5fQscaXjR2QRTW8BAc4D5Kqrd1E6rLmmElZLKxKi6I37ErMiQXpxH/LXcO3C4tlU
2Ni6tleaiTorjwlcHIdkqbwLrGVOeEHqEcfQPbACv/VneGRHjQ8JHRsbcRz0DCXk
dcmhMOUkjim0bz8wy5zeqnLQOaGNP4I3k/DN3kIvCtGfCAknfBxwflyQuf3NOpNb
wONZIrn7Y6BbxHTKhvqtlkjLlymPqG07ES/kFe3jsHi9W+Ey7vNXjKr4O4JvA4Hr
MZwhmydSuSWXeUhepYITZRVKhsK22aG/tgIQ1lOQnMXhhM4tf5SdMpBwTZKHfwEY
2hbRo25SwluY5sC/qetzVDatb1e99xFpWs9In67olpmngTSLo2otMj4pvDvAMoMq
PXnlMdRINAzZXhHhf7mRpZzOWv9SQh4qp/B+ZjYjGCRiRF6ZpO0Y0QqOYWLv/j2D
hn/9fqan+t3S622Pt86KcK3ybOHi0zaG4RGgotc3HoTkXQFAFqdzdp0idQ+9TUD0
WgQKQx1ob8t+/ietZEi7KquzOU+5GEUtYbttcDvb+M3wGMCLj/SNL3/tSqc9AbIT
7jmDcGd+WC9HPgAgbIC2eUaJSEFf4vGJy17tQ9CTzfYH46WRLYgPq7CIbWtjstBA
ZolyASPSKM1Cqdw8LYI+nj1sh2oV+BSpEcNNu7GTIUHd21LCeRW+V5kkVMySuVPY
QS+HTZUIN/noulAJd63P6TdcelPF79ff9zqDYQxVubhAFpfrdxXWGMkv1yTjuSVb
x6XFHGVRcGKRmX2kRIQ7Fe41YEaiqhUTpaAX0qkjIQ1p/+y6uD5enuuioRF1b6Ce
t67OuFRczkxZjTfpbLzKVqQ8YPINuSku/eq6KYFtt8tvAkCEIvlPms9O1vZOYPkx
4fxc7WCjU+P5kN0ZaoV1ltmf1w/V8cJDfVPrxWq/HLTn+1qMSVn7XK4E5DzO2rHV
oFcdcvAiEacZkZUmVowBK+sghmeVGzOzQtwY2xxLgEtIb6LfI9XkTi4r7Ze5/hGf
h8z6ePQrZqXhUZDtKb4tJs52CnZTw531uMo5USREQPSskFyQtd6Lm1ONdFXKU+pH
jg4+S6BoyLbb5rvjqfA6oGo9pPLUTqOgCdwDVhF6LtAkU2viXyH6vlfSfo/kMUbU
gcgXcxTPQeXztaw3TAaU2jLSqTNaWyoHyZCnoX9wlgF5A8F2tnEmDqUoIy8kICi1
ds6l49i3pObSXByZTE6otn9/QgenU66rCCyhrFNZGclZnU+vfFAVBri4nU+V0nPx
vg+q5NMZttqFQ8GCY/VNTz2Gla9RDrkxsJjevgybcCAYCnPRya8ndsvkJeRyimh+
mt5w2h0KbtXOSvIKBo/i4Qg55X3ip0wuSflF5omwJvR9p5CNLGBgjm8cBfOQrrLJ
jH7iXWCOP1KENX6Q2g3pVJ1uqzEeQP/An9Fgk08Xo05+RD+UzfWjTjh0TI562H+D
HTbvHEUMjobv7tKey0HsolG12D7DX9AEBZOAVsEDAahDluUhF3o+zWNdMI02F0rO
h+/67121kdGxoZfLFZtMrhlgCeb564DrHKZwHXd1r/otKM1Uf/LWlq4OFvYr8r0G
K91NGepQ4XiXS9zZs/K/gbrLFX4ig5LlOS37WziBFOhEg5MN5lkyEMQP3JiWAGki
A/Z4btanSf3uR8hVvHxuPK7DG4ppOoNJ8bsRSM63NJPq0aJa6c3cUCx5j4bRBiR/
CszFOGzEJN7AK5r4VO1V3aYZHCRQ95DXClAztCeExZqlj4fE0u3ecl+5nl9eFcqY
XXTNnPCSfYGTmAnrIJ0uMdWtF7GZSVIKhDQbw2PRK+Yg05HCol3GBu/asbl/Le0U
cw8u2L/yzIUsD+3onnNhYN03j4dN3y520Y81filC1Ld9vr3zA3DL+Dj3Wn3jWVM+
RAUmr7nhwXV6QFCaRzRlmHSj1T8k/ifNNia6uMbeq9Da/lmtX46d7SnwxfuglkBV
/kB0+bz8zgUCKA6V0KzHU9DTQC9Q/aYIoGdPEKJMnjoSxNkt7D+PcALdpblJXBEg
80Ex2ui/jnDojCzZGlBJTslx807lypXEi9im8j+qB1/w7dNMaG2T2ikcTXthPs4Y
0BL6WDQIXjkXU/cOZayDA6ipvAE1Rn4n+XU2ietHwJYR7IK4onc+wyimO4+/3N+j
NlNRo6AqGos3VMS3XO7c+lRCuFT5iVDS/q/1a1RwQdgFtXz2IOgYUlELMIKP1KJG
aPeB+Y9SxNl+L2lg5nyl1IUzKKCUiQJkpa2Ti0MZ0wJ29IcvjLvSd7pVaV6sNuS4
Ag728eADPsFTy/D6nrQmF7YMXJIAIGHXQGOo+dRG09nUf/e5iNKizigtKhDQdlmW
1kN/Cu3o1OqLQDtY7jPNOKQCwXE0ZFDUSXgJyBiZwhIhTOdZD0j1fqSAEt0ywK0k
W++GzU8HqoHyon0ZhP53cX11OwDBl1V7a/lyytIoZxtDjHQL0hBjlwziDHsG38p9
oJ7uNQ4v3KpEsO0igoQBmrS/LdSlTUSyDVwkKoe6p01IOqNrA1gFRzOYMoZ73+rA
O2BMImXf+ctgt6EEZrSk71RPC8E9HEoS9IrFiUDgUYSh7gcB4dEgYBrFvzIz9RMx
Xs9Ux9y0jxtsbxObCtBtNcvQxp/IzvES/mK/fefwBwSrptdZOX7loAkXHMewghR4
RXEh6WpOAyk5Ao7gC+LhE46XHgin0boJ5rlcoxWhx7ti4fGv/IgFL/HWYq7TDRET
F4cQFLHyAT4W3lf5EsKpXF+aCDJddHX83gF2BWIHvaMY7acYefce+gQB5bgPsvGW
TUh0XAxdXnkrzlKlZG4rMoUUkGPfNXu/XQH/qdCHRCzoAbcUd9zVhE1/PRJd9EhG
1UxuMSjoTOK8Q5nRafmICTddFWwV8ZPY7Y4dCudY3XWOr4/X5dGpFoSc31UBSVVV
xyrfT2+6MBtyx0LbNgfMKKWcjurnNqXTr9D+7eEfC2mRSlZ/7TbctMmWhZ/noBVF
MJQ76g82GaQ9q7loOWnEUWOqAf8Iig0SKea5NB680fd1E1rpAd1bYYXu9eMJr2AX
r8lxtOKZqzrbws+5pwaAP9RL035p8d8AToQpp71eAqnTwwphqoKdU9OSEq/dWvFV
lluLNUslvTbROMuGzIMR+hBwz3ki83Hu3ppG3u6aSeBugRaFRCmJNU/xT3BJ7N19
LnkhF1OOvU/h6MoLTUR/nZ58rtIDu+LHmxgrOLDOz2FZoel8EJe5Oz5zdscOeiPi
bYPcMRxD+BKCPH2sPd888EHSyQSX8dxrtMn5Yt4rDnHjtLqtv8X53o0cj3EiPRN3
VK/hmTxqIarOB9CoT6recWDgo8c42QJEqWzVSjqouGIIWVkTioPO03LnGJIW7d7X
szv0IV3kWJ+00kDGBFvvpwtdlY2j4Vb2Aeri3vCC3CaXbCj+kObhb3s0Z4JaCIRB
0V80ZKUmXtw4nTNI+n7jPaJVpLq4uJfTpxy4gw6ys5oGWf5EMGfJpiBWUaCnpfGe
1EMtCBr+Gvpuk2qXOhJIUzCkF2cimlmECDeWfl9JjkTuK0tqjPfprpqeVWYp5Zgt
Ruvk8062O81/3fRwDYKg3KchyA/sXwFYrhccEcTWz0QI+T/EGG4YcM/w2qVhGYLq
w3fP428P/pFRIetGvIQHA5BbJUyzwcRLapQKr0ho0aN5x72jLVB+s10SZuqKksgf
PJHdh8lzjgTLw+4VqJn/wHpiT+Bobp7HDFPctb8mcNgC6hjUYEmzuG+MqcW5/Z+T
DmztZPvH5TanHa21+BddTikuO2MZXotzDNrw7mgyLVScv++MurTUIWX9VCSaXTMw
0lVc+dgrfxuEXbGBUr1K/vq+IVSN9JPu/udrWpjgRbHWDGwNOri0Ol5CO3Qlch3z
rU2B2nF1mOnIpCyI5Poat8BViCod0VPZh1jj+UuJAW6WxT1NQu9r2xekl0F8WoGu
E3xvlM8Oyib3U0+B2UVwxiq72LErpR6FeEjv6mQMPZ5S/3Zpb6kVU4SSmHPWUlnY
jdbv08REcP9ENECqB6RK9R5um2HXj6BqCWOGkm7FwSoTHBOpOFeqLeiztSZrdIZE
Bfc7HSvCrNJ1MzDBDwJDweQMuXVcRlM+0pZvTgwAZAYqFVMFtFlz22uEbM/w1XOM
RfCQzfpQub02AjWgm6Rj5/HyBptanla+xifmUkTbfMzA/uxAjIj0HIfWtk8LmgG2
XFGBsP9hOP8IBNN0E8boeXxNsiFGzZsNR1tvH0z7O3U0VKePeblVUzMnKTIpHVSo
Lyg66SmgTzMKyLI0MHGuwq3EGiMVJwCxVUYhruRnOdRdP2JCIwYvmnJL0u5/Pkyl
HQ/3ZBV4SpHXNh0RDt0kkgynJiOzvECkbCt5JFQXHXgTk/JGIbkT31Cc3/qNFD62
gKFi1Vjigi8n7bI2lK9i8+JaCErI8VQaLFGowrFo2bVUGkR1YeFnMGo8PtjJX2Vw
ekvezS7kaIaD/mL3PQbmjH5pJWhWVeDW6iuK1utFH4q5yOjWbJXJOTMo0p26aX9J
n+BPrGSxVuRmm2kUQ7//wRLZ4u+amdIriZWRRkOZVH/UZpCVGNxbcjPmAiTd+2U/
/0epHgB6BMY7a5yx5HGhc2uCFnq9tg8hVH5v7OvqNu7UC4xCsujUJ2hJsxS+XLn2
Nu8ttNbO7OztfzTnrwvvj40Ku6aZu/rkDtwYmpTxLpm/8bXuXPo0FedQ7fcGTeya
QRcWBrKGQUSTH/wvdpjRDNxjqppgb54Aw3PEmSQYVZ1pDfgkvecgdPp00ttXqdgS
U1oqscUDxc6zKFVemon5lR4Zta5BRx3pCP0at1zgCzsbb2yaymJBaIZMYKu3A6OV
sNtZCEo6doMvG7ewYYSf1DoVgkiQRnd92p3rc7F2tWcf+p1LtKnZjia1XPsfmfCU
l4Ux22WObMd81v6abZNylwPuVZdoEu+31aB0fyi7SJdFP1OnpsflgX2B6xaOPyoy
+BFnAaFCMZ2bjp+XRlhZAqvtRMwZsxgQmRAriKrbNADcqiBLd9edvEcBCwCS04Uf
9QuZVQpQapNHkPVSzJsF8/iIBGFgopJJMZCcoG6WrHBJX83tzXN3p8lYediEbwtx
l38/vlQvv3q5mms408PtD8UBAm1hEdHo2J75FVC6Q/53WgjacIP8bX7CRbRFn2yR
sp/0jigwVV7YOrZbOMDgcYetsX7n2vBgxLnYlg3FW4VNf/dcBOSw3eRwxcEy1jpp
UWhfQwUFDKB1AZBAoN9WEwmYrbwYy3giL07C/Up3KTCWtsOeCqhSTTyP7xtkwSOP
JXLi4U7dkgEluQtrbQm4VBixL6F31zObc7m1MWp+Usv8wwmrNZCmzpi/GLX7VSjq
PkF+bnzJT3/gJfIZi1tGUfyZCvvMVavWaegSK84sxVDWswpbKq1EbiBSHaPzlw5k
5gnVpr9lSGuA1DD8RD1TOdMvnQJCbhJMYgGw7egKJR1/ZT3ZXqXBFHIOfLf3TauD
x989r6qba9/53k1hZkv5N13INpl8QJ2t5gfqaB9ttbdw2Za8+TiceVhNTqNaE1Vn
6QEMEoYzMRPl/w5PQffMTdsQcX+Q16n5Y9ZW6rd4+4KzJjsRuNtpOpr+yqRxW3p8
NfcfWEXtskgrUGg9HsfSOUgOLl7RaVmyOVL7WmdXNpzcWjok1KK71G9Uo9fnH0/6
qmrwV557oTN1noztqEIc6Kz6cBFBJigPoh77qYy4yPK5G2LLwyU9Qe2UfnXt30y7
WdvV7Mnj+63A8GHPnwMO4WEtLnvSoJZB/RUMz8u+ZGLvpykFC7oXOyiCm370PpOX
en1m9VOFvAKCE87N0IgvMRAbneWlq3WP/A4G6YQQnflYDbBnJvmDye74mWKB7+N4
hwuvzRcOnzd6PDkMAKcBjpHTivb3ROPpr8crViMV9G6tB6cPe0myrHOiDyYvF9rW
QSPNI/Ez3N1M+hnWSPQ1rgSVRvYQLjXGNPbPQQ8UC/xzCOirS8dMtTc/vxK7ER4K
sTTHOSZx3nSzUrF9t/XxH/A4hMtld/d0kBq2QFuQU49dbRjhCc3+SRrR3W3U3fKO
u4VOPFT39IRYJ3jtR+k/d5YNVIAFWRL5gAdgJ6RoS/YoIGw8HkK944ZK9fC0r66w
9V3ULYYmTJmuG4b13CUjQyhNSxug8f1Qy6zZNsxmv30k6jQwGBU2+cYK/v7m0H4D
5X9QJVn0/A1A/5l1RfDuLtwLWGtcSn1U3iGcWYrqHrSLOkciF55DETnZqmLQwdsO
HAFYKSevQ5o1AeI01+UhdeitSkTyriPDMa2Obk7Osikp6HlAAUFMq+5owXi41UNL
i4xr12ZNf+fKzteUz6rhnS/O3G+wS40di2xsDC8Tw5BnZdrsMC+cDJ0D4cE3upzX
YA19Jc7ENrXz76E4VUvDUknGcpMo3u8dg5gFF9dPtDmVSv6E9EnwrG48M3TkWkri
YzfoK5wEVbW0cms+eKyeOTaa+Uw/rKt58Sip+4MQj197677ZvMLGr9ROkaBGu+gH
IjjwY8rmoiQlboEIE+mn4INKi61XEoH/wQbxL6teh9rNORFs0pHH9o72DTHgfjhW
csv7JK9ZRb5iTZ6jVsuGrZfLM1Q3kA96f8AfbftSWUM8kMJCbkSfj9YCDQF+nwOD
a3LHe02ARmVKGMIqdKyrH42pkNXmjb9ebTqrtuFFF4sEgzOTxkqviOrlqMnFRb4Z
99gDo5NcrkmlAfhfXMXm3SevmwIUUF/imxfVRql77ZP8Xa1100VzwWi2RU9hIICz
5blyVnb/SfVqCLQolTcp+Agq2RJfdDRSTHGgNyTfHk+1EbWFJ87Cj0dps/z3OIKc
1kIRUpdHJXz5aYndh2/prK7gBVYqr5IYD8CXztIhpJJXz/tHfCS8VgLjnzjXDyQj
61/2PUVJC0/lpoYdpyIQ5lBEA3fD2jmX1Qe/nTfRknLFKX+4Y6j87qnJqkgpD8og
siyoYBhV8Jh2dxuYWQ7Qf0T/AYT678MgZXNUMXlXTI2Ro9H/wYwqJj9+O9uN8WKh
K8PVr5ntztV+rn40XESHHpdj1tFYU+UnK2nj1b2Q9+LaJet7e+vTc5anmHVReNDl
sDUXVQvFSHoL+E/1LDb2oWQ0Mmkqd/Eg9MXB+32NYLs+bGd8LxBHS4hLDBY9P2E0
+hHDG+AvH6E6C5DQWfgOSpPB7gElDfsqp73zkELn0TOrazeNSvwa4h8uO4OUlIfC
au9/+FKt4uGySJf6S3pp26+w2DcrIuH3G0SSl/PS3LDsLT6IgwW8SW+QIOxtGSqq
/wCoJ4whXh986cNUNBS7GekHu9DnAFS5+mKkqQgX4tdFUP7T+SsAwHH/ZXrISKGl
JfxwOKDquNzrR73CuAiEYOzRr/0G3Gec4Q/0e1x1VomMjNZaHj4XbF18yx+K9N0h
2aa3beot/8G+91jxHND5NKY/IHVEBSAUI0rGFOXJWeVaRwEYnGpvKorX5zKLJmnc
spSyFosNXsvKNQal9rd15MlK1t/AV4jspBP9pD54Mb+8+sYegjzKe9OjemU687Qm
6cdB0VceLPCN1vOfL8vtl7Snqrf+LWtnJCo+doIukQxFkAsEe+VzGAVsqJagkEWB
AQCdHu9OC+DpOm+6c2cTaS7Xf0RGUMmRETl5nkgM+b16wy+RNLCUlPzOfR1Wk7gU
3KcdjGU8logaOVJXLx6AE52sR1ho2SBpQ5h2xL0+yYc/Z4tCg0y5ZVSYq1aDiA7q
nq5D4apUqg3ua4ahJoWpjzV6Xx5RwBSV87XMJVGjSD8nbl7K6gbsN84VTFbIuo0D
9GkVSAgzQVz4dmMthO6Gcms7fwdsCdD/jThfLe4fP4g/yWue3YYeO2ZzGPC3zU+X
jAkh1nUJFgYwZlLEvxSPEmCUuYGh7Ft6zhRqjXiloIa1CtF8y3kbTUm0lscLYA9L
fB4Md42fEmWwBr4Aag9clVbx1bjickUF6ej8ggo87PIScLlENl0sSxEMMCgrXIhi
sbMWvZCYJnzL8UHXuIO3CxB1lslII49Qrno0f/04W0oekxs08utUvHJgtLOzzb6E
kCKOnYfqlrQ+WaskiTaQdBoihQNk04xkCAzxxb1wC4WZHp9dt2KSNi6lbzhzJstl
xY+mkMBJ6SylN1+NQGdeJbtuESKbLxswlbdiP5OV6jHYaklLqz+ahZqqForWuJwz
56EKB7XgqZEJeiTY1eciO2M6T4sBxZUYuwQTS9OitrTFq0xLP2FhNSYDxOm/9UlT
DqHjaikpBqy//kPRrKFnDf7ZxnmSxrTnQsrs/wCdWzrr3wGQ+9OmnH/WfB0p5BBs
L7DkwvUqjT4fSm20mf2oGfbAKtEBIAM/2t3IccThiq5RACcxXL20qkjuyTk9vvNx
I0J58CG8MGWIUHhbl3Kur2hXzxSNYCcg7kfIEVw2/vnTuWmhGUjyGRXVg3zonEBz
A9E53TLN5SV0SyOC9zLmyLQTkc+ANZSBxu7c5vbDqsU7dEfMRR3zJCGv+q6hTumm
gbAf0mn3yRjo+xGwZAYYjHyUfnyGprgebc1NBwrF69MBCIKq6jW00W2f3Uv+FVgj
KI0JAJwsiwiecS2yVt3Q5Ts1ZeR8K70eO1P8Wiu2CIlwULjlAbySyGv9WyDAjLdb
e5gmwV1wDqZbDsYETPT0VgRTbZo9mRjes7lyqQaJD66PboGLgQiJflzTE/YfQHEo
I0TxZu575GrmD9yq8qhs+JkIi5NCv+/tOKW+xrZcS+G5XaS4V69Uvupgvfa5Ce+l
rP/kzbhei02Sk3HBkguf+5RZNhaXRrEsLUUmpWELjmHDjNsouaqGEAJqScRs4xZf
Y7O5zRp9yTM3gtcYnDqRGAEoFn4/4Qt57YeFRBzjWUkXjNKumxshHKCcjrYWJYiA
9+KfYm8LgkTmneLL5DFqd1/ZYI36aSdlr701hZooGLyyRiT0Xd7RklhlhMGNs+BH
HOqiZtJdIScjExVOqeNdL/7lmdgAHHDq7dMZvJR3WrXsiM4D7OG6e54BownMTnPc
xLBWghITxF0Z1y1KxClp++LYBhlpklB+u0aDlVFSLqeg4x6JH/PTaZ8rwEejHqWw
Fe5W+reNUtqmrOb+ke9WwQEiAWWI7ZRIwxo/T7dJVMgb9OjRrzeKSCRTGI1tJwxb
iTFFD2zRClks6/US9MVY7dpAcUZ7NC48A1VU2KO7AmJ3dAGiTKHjP1LlqGh29Xt/
FN1G2u1tcXNStZJm2DfZ/jMMDKcdjguYLpFgJOe0O9mIZUdww7/bs8rxfcHUPoWA
lFILgibhMAvvUZ8mlce6V2RzLdcBLEWNsipJwkeTn+R8vlN+cayX3NiueygtuIwS
++PGa3cNe0iP0ei9g5vRGkBNEMBOLbW5wFdYDWoSHP4McTTe/HFZYBkC/R8JPGGD
waMtNX34OUhKXGVIbzci9GRpbUom1ACZ6Fiozwvi/fTzmcwHfzWTl1/Ofy5DA7UX
pWaLqSI8WyZ++deExSep7IcXP/zq8ZGDop2Ffym9NdlgBRxRRhWWr46jEUTIh9l0
ULG5bU+qJcIUBjhHtCyOcoMA73TOBeMGu3nQzat2uxi4OiaOpwmWr+zNVB/VS+mH
Oer/CGQnJh+Wm6S/oxpnMvZlJA9NLjLePyYENp0Wylscp4MQ5+7nJBSCGP9Bc/X6
AXmuB1hVUbXMSMPOLpQYA+YykUcxD4vkcWYciiUEOKJ3FEeNdKxHAnDx3wxex3Mc
5Gs/bWjHtGV0lMLrhoPhKh3Jm0uN5uctcZU8JAi3rv9yI4zp5mbV8jCRALNvuyKc
p7IonjVEj4hJyc8H39UEb/r+nmUS6CzjcS3dZvFCn1MbFmG2DCzGfj0rJbMnOLRd
GeIEX59ass3SZKAhuu18mIRfBUhgeyi+JbVEFSEijb9kLxmN05MFuZmajXeon5F9
PS6H88Toh30b0m2uroaPyBQIXc7H0hUqDKxEpv+6Q/OXv9coXkecWiF4ejJkp6pi
3XdNDWc1obOHogbFm94UTnj51ceqZsJXE8SLZ4ScSLzVf3iflVM0BnkxQ0G0O+Ze
/D0suSqxyLahkyLVjZXig0cfsWX3IKZCHj28Y6G0VnJa4p2r7dGelZ2nwjN3KBj1
l9YHHlwMgyJ4cfgVVKTA6zLCRBeAz3nFViP6tYvdn5n5M0uOozStkMa4oL6RUC9i
hVE5l5o9QQ3UGOO7CfDt39zt5+fowV3PAjv6/umy+Lw/BI+XcURGvIKpea+R8u67
Y0DJFnbp3wTbIyTF0lvDqAg/ucq9EQlr3UyJTyD7z6BdgR/02ITecKuF+aFrt/Km
ryphDIckJkqtR9O5bocqQG7xM6Xu13zTAMOQl0cdVSeY7wf8PdgnT0pEGsORRYcs
EEyIwIo3O8W9xGJmXPaU8H7YeFw8OkD/v2dRkJLm2fmdyzUGlrJqtza1DQQ/5w/g
zMkN6xITVAaIQZ2RTIim6tUnQkX09zNV/GpuBB8Pijs3C3B+5xOoCKuf9kNQbw4g
k+ArC6A6s1AseBzAhEnCZdGOOHUda9TJ/MU1Obj8PNC1Bqv3BpC/oQ2m5vSydND3
Wnd0I6aR+2yaTdJsfUlwaC1fu/Mzu1vVknAY+HIAdZw+6c8Y0CnUE+CzNc92tEse
/W+DbF3P8Je/4HOK1YeErLIZI/jMOFHhX+K0pLhOR/vgOF2ncttDB2l+uZccHHga
pUTMW1UMSZGqleQadWmjdi5kkUDax8YAy/OYbWNAlIj3iysnEb9rXzfy25RrXedM
aUUuapErpQTIKqZ0EojrNrIYdY7eM7C5AR4rAGDrwcyYOCo3xDEWScCOCFcOT28v
NE7laX3XNCiAazMOaJzT00Tcv7uEth1qHFCiPXHxUGhOG3VAEhmgzhy69m3Q8sS0
9Sf790sK6i2kbVcryQmKUCQR2XiRf0O00GQNzeeCMR9Mpk7PMIaOhUd96CCFCgTd
qW73I+IhkKyN+th1uFcL7lctvzaszbswXLiOGvZyeNSmh8e61Dexj/gyXdkPOTFh
LkN/50hjbn+4me75t/MnxG/WF3DvxbySrUpBZWfK4KS0n/U09IDJgzzYvluKo0ph
SFuKx3YSxrFVvklDwIorVAJUKRFjKIpKPZ49wuDqoH16d2UooEaABKsue+ji0olw
hVq8X+fRqDRGixLkSUczxDMLtJV1k466nic55w4UBG9tf7lny3IpbQE573KGl89t
AfrZU31c9CmG9152MSnOiMs0o6yRkJvVGbjhHG7DfkFpofJT7VoTzMVA/mo3AFZz
OUAwvJKNWHpODGjtdwKJ9K6GDZD2UkwrVZk4mKeG2iKuKyHdWohN4JMXps0dfeQt
A0dTp2v8jTIlUe3FykIrb+xDPNfVeKGqU53dfJPTiR2TihUzUM/A1PBv7anTL0tS
cgVJtMa8MNpe1suecggtPby8Kaj1dYlCw+rh6HFCUxOV4bN6mqHBpEYwruTDRVYz
b22F2JuTXJMh8PTOtyZ5IkXn5uWcfvIbKhhNLUJEpE3CiLf1q8fe83CjryYryQ4f
3fSf4Czv1/XYLAtCuuVvTxLXBgupLpHSfpDbwVKEwQtBhx6kFrls7jKfB8d8QIS5
OcdBsqsFyDbRetkJUjE41AWExw6ASpWoFVVJKEyu8SgtsBjvgMJ0eqDX5bauWWVD
KOQZ/6nvKs8MiteyuCoBhhGFWbz2agjaQbqUg19PX7yZjW/TVjwTS13LsXGUclVt
FbMtGfKQ1pMYZB51cPeRQTBZSxEh+R2ociMY3wKsfKkxGHmVRg0Vn71IyiJt/dBs
swP+7/AsUppVjds2HNxGId7OCwrhxf4S3+ELu1hyPGmfoQcmV1J2meCKBEuUUBA1
jEqhZiO3E3rCh5PUnvbMWKvOfeWDS2DvEjPZmowF3NDiCX2ce89/DURRHgfwvO2M
sczHi7D6PSooVWHQ2m9sWm80A4EGyH88l5eY4LVuVD3+2QI++bkWAZcX5vwhaPSv
cxFzsT0YNO8XwN/stWAk41FZyTakGFw0SyfqKqZeS2+daQZWuV/k7FYQXOsBOypt
PVOx+7UTkCqaSGHkfjXFj9hem5MsYEkDWv/lH6JmYw/dUgPKIGLEnIcn9t8mnF2R
6kO+ENxBdRm5GGV/CCfgTpQNtSLQoj5eBneMshgnkzO8XGwi6COnTZj7eY7iq5cZ
ew+hsWiVjwv7/YxY4yFLkh01C/o6F6tzZn76W7AwmeZ9bdAJ1uj7J0z344+BHZHf
OtdzdXNSMtl2rBCIIXH59gC4X18UJ3r2YLdEF2ZAjOHr1xjzLuwBNsrPnv7rTuev
eAnOhiweO00oCLycOWwb3kH//dchuzPHxg7PHNEJvddr6TDEbMHZfOZOqN23LWox
WOkbLzP2Aj/QY+1AJMNjvBD2U6lt4tOQrM319pesADFfRLIZKO6DCmFpbdA9Q3pr
EwdjwbqRvjt7XEFdBnjlplBcEzo54FabXPlVWMSoCtIMySdwlU6dYSCPv5eqaWYd
aiYywAc90LWUr8n8FQoswqcbzoGC9xYSpUWdnJsC+Pa8p6xW8vBh5HrAieZtXHLX
hKhn35l1NTbRA0t5QwynhFjUFFcGZOhoisRd8jzCEAKGBF+pMUAG6y72iM7tePph
iGtPazWg/Noiqg7IBB2fZUng370t2hld5cAC3LF9DNtJE/N2SeeSUeufbP4BoUlT
JuKpPae5e1Tt+7b3JvTInu4ygcko+tDk6Bs2f2Bu2YoKthARtgEXfvvg0vSWQIMO
MsLhejFzjT25+9Gf30KnVEdRrwwyDYBJXFOJ1rvfxgzskUurox7VLUL6j9WHyyNz
uAaNr1jx6EKLVF5zniuPvYQKPL45NkrOhqAEV/L3H8VYhXFw1W0PILyMhNgsMgQI
8rsHv6cOhwrEPvpx1iZidxzVoyY3ibSG+neh1UtHAcoLPl9ullubtnAyxzVd4Qgy
tIxgoPbz93HVc5pzOoQquQ/pNo1haC0ym8bvCfHxfQJo9Q7qV/xm9XH+bJwtueRo
EmyFTscFHRrFqZYjVOfxTy0Zeiuz4gr644C9jbX//ZZ+mZo/XTWeWvXtWh0GQ/9i
DEP44Y9iUozvRMyklk03Rcux+pWC42e7jE89JiaotH9iRo4YlBVjTbnGM+rUAuVM
nm7D8lwJq0ByZukjGAv4mBlcGyyDlRAqndTpRTXNNm9EbfoSpxv6URNoi6NkdlSq
LMDIwNMex4iwLGgmbYfMmK10i57ottVAC1txJLla99Xu2wm4rIVXKCVlSmiOKDhM
W/IsLqrmuN6lffS7A+lUSP1YAEuH1UN0uxdcgFvbpCWShWXB/JqwDnPy6aopEO9T
r+G5vBmoUPVaWnN2QM0KKsgnrXMTXkaRN9ybJ42hTYXMBX/p0bdfP5npQtxe8Hez
1/6cfr66+En0Yx8qHhvnIx6pwT5TPIw/jTQkoVyLv0GO6Pp0Lo5BrLh7/GeHBbdZ
BvMZNAGEjHQ/qZWUP+UBIE4ApnRZy6sB+/+ech3YYfqT1GYnKhUkFpat2yuHU+Qu
puPZvT/WSH957ZCz154NS9k8wf/hxmFMKRNGxyYT9MDlDVtfVcESnI4zer80DDWp
vsud+Hw1vafOOR2bOL6dcml48eOHkUpmSfXI3kvEnpTbTcOaJMocimUl0uaKT0wq
QYK3qxsmQuUJjD/7ajptsOTcCS/yheBXfKlIqv5lH7Y0yRY2XTFMx+eSmwTdatDe
Bdqg81HhtNDUGW7lGbvUgLaTm8pq+557B7i9OyPUtKczwDjOxTjsR9JiFz0UAfxE
MRBXrgS9oBlmxeFGKGOwaIWnzi2zrrj3Fo038xyv67KCBV/1VcGhv9BB7UB1UYR1
FThCUxYR8vG/DTydOHCPv0wECZw70bos/0VK3nkAFCt+69G3USR9MIH9pVAaqZOf
rPjN/hZjiYWLrzFxJl7nUzKGF7a9paGCJ+qBVla50i/9zlrlxgn7WrXoN4hCcmJF
tqGheIrGZoQS7UVUUJBF+JcWZtut9saiH6MariR9adX6gf6zR45bPSbdFqlrDjIS
Ob4q3K2mkSWdKIZ+92oo2UkWUjrv5uTPBFAdZpGnmABSmWi5liAk/Md6phGAcnOn
hV3rBVsxvJFkuhX2DSpTsJt8uhlWT1udKeYAk73jA4HjGPRbA7bd2nLiGyuZbaZa
aLHv7uyWjI+7nxmKhxuMa3kkbQ7TA31qW2FIfI+o0NiJ/Tggd3E7IkW1o43lQcDY
+oILEQfBkAH55aYYh1NImL6z/lhc6O+iaS9szH3oT9Q/tvlgkNRLOfYVqJlVnvDn
BksZEJF7BcCh2szeEFTfqzrveWWNzxshkEhWEj3ZqPbxgj0Y5IONwcDS/skzdqUj
+0PCEM9hkGzInrDkKphO8bav2ANvTEKBPTSfflc+93fG303eJ6CjOa4XlM2GH2Cf
iyB1sMH7E2GHrRWcNxgKj2KAGc9wBttKkErgteK6E13I+4i1HMRHSwHYU04MEA6+
7b9JDF38S3CtwT1jbikCYxo6bWetoozk0b6HMbaQvwqubby3sUn4t7jN742X+fp6
yoILmku0Zc3y01lDBSudTfLKHfmECVRtMqNd6Zr8ry9SgOFjwo/np4XPu9zeWw50
/ti3vlZkPYovBSliTgVJP5EYSOAuIZ389JUfBpICv1YsGl+UNoIY46gYWq4zAzgP
918DC5LF31AVOo7lCWRYXiCpI5nThFwwXBXPgk71JixfLVKfMgDyzk9ZB2dUtbN3
E5giJ9POPnjdpRhRONUl5xusDGsQz1PNyrnPqZosDaAIh6aI5sH4S6au47fC2cns
Uy2tVBrg3NEchDH0s3C0n7jwhf/I8Rkk5A81eeJlBlwi9fVFL4SxxrgqTt082eJQ
1u/dr2Pxlb6WL2XW5AcuTxIcrS5uHg5gNNybsm3n8ZC2BzBIhbO0DBvwlKugAoPp
3oDPCNUWFVk9KWun+yn55D+9URJJXjQ4KMC3UsNtquOB0xbTGsZnsaOiZkdGI0AD
8j0Te0qObVh6RU2iMe7EoeyKHVTJJiJBSfJQoSe+lm7FilYX5rgLyOFxUDS8GQBY
+Q/p2FNtqQD8IVEX18qUICZ77RkOgKEvLjfMyQQRrEZWIajlRsHmI6f/g8+ti5Og
E+ReVm7C3X2YikAntLUFuE+P6B7bwMqZEBiBsH6IOkwpn5m0bUILQTL44FxpRixu
ZwKlwsYrpyX6X3RzG4hkzepeyYCVkSNtSSpXri9eib8bKqmXyV+KPf8K101xsZ4K
zdTi2T6iK2R5cYuzhIuTHpxXausGrnq4RGUxBMyt9ZGbh7Z50oTUQSvaPR9enf4N
BnGUcWlFbqaGNJSXvortNjYVarOnb+m/53cXVTNsToU8b+RZYqLQeVTFzNghqx9f
wgOqnCTfl93yiDL8JJunTrtA3BDqX0jWtzJuPcbHuECT1VE6STymplQYKeCZw9VG
+Aea488Y+UAhPyf12fgmH35RV4jZ8CFZG7/fufUDitqaxPcY4MWthKvWKbF6KsWX
JkOOC/AP+/KF5k4TFuU7dx8jUagejy/j0ueNFkaEBM14ubiGsC1nUuiW5eacRx3c
1SFDDkza4qDPBwnBN8XPDAy7Vblmwh2Z/S1Y0gBz5lY8jlZpPiq6ozJWbGezVjku
B0qaboOPD22uCG9tUab9m8ysH3I1mpyqVqxq6qroyXel9XZrDxOHoQ3IBWW6as+h
16Z88aZx33AJmWaNMoO2RgF3yu87UFwJd4Ivu/FoR8QEbstai/YJMFLrcgjdoUXO
yNpBxwYOs9zWYAAw3Zo3D6tjfEMnMpZj43TEobb3/xIo7k9+t7w3EyA75vBwaPjW
wmoC/TcPmK9+Ax2HaPrmEM6vQdmTDh/vq3wKf/QKl0u1OZt5bnElwc1rH8qVy2fa
ZSZ0kzsJPLLlYCsFE/oTgABNThogEuqzLy1MoWLwETLcKfd74jxH9IYQROnJjo69
cDk4nEJhrq3joGqkyGhnARJ54MeRUX9e/NmsTxIQBek7FrU4HIIFRrwGHVae2LST
vZK9PmIlS+vtVMCqiXjxBLqggfdnng9yoIwjYNnn5jVBgV4vZ94o1v/EQiPD7Xrq
G7d6k4+bDfmyTDvPro7dr5zyGSvKmt6ZHIIAYpt+SvE6tIWTrf3PyxRiotBucpTO
DRYSMpl1m+g2cDmo8/vLBl+X11lPKZrIE5CMsQHNwNRo6O/MSkfwx8petX/6r9Pg
wiwV82Hxa0YGkmF8FBwWNMPNDE6vPmpUQ53IoSqF0o+y4Cr3CGMydpGG58Wjcsok
ssv9t6YxcRlMNODcFEa06m9QGd6bt1Yvbb/a1U8i57NGGgZ+IPn29zcr67KJmpeI
d0xDutnS3EGrF4TUTl4oHfsrLyJ7IUvRf97hob11Sm9X+ArnFORrvHqTG+h9OcyW
EhkTpqjzhYGjoH3AxPEg0gfOVFbjr7skPC9T/HEHs4rA2LgJb2JGKIlVeDGZiHoZ
pBqnGg2Q4CkjhnOqhlmDdCjy0Jg8dkU+sDT95NstQBHNHuEQsZ+Liz2fyj9P4WZn
fmLnV8Ix6xRrPosONIH/F1pRxAjrMvYMQ8GEUDCB2o4y2lTcV8c0kQdWAPk+Ff4v
QsE8CvIg9YwKb9+IgYIdI/VbhcNn3lZlPGcdBrxuP4yJV1s6usuSUT88+Xw3gcum
UeYvYaOQcrG7m7oEQOdLT9and2+WS8CJu1w+hCrjYYbjonmkWQ2N63itfQQxmcmk
tNq+mW1PhYTblY2s1pY/fQAlQHThu12vmQc7/KqURi0C0g2C55CHtuFdrywFnsMD
o+wZZhWyvVw0jM9A96EGKl7f7oKZrXcrdWk1xc3n0P3hci1CW8ep7o3eiwGvEhwx
wquAq14TVSJUQl0J+UkMC+m/oKqDamD5DLDUFe9fLyTcPN26VeLKAEmCknwLtWyn
5Qmod/eu+qc2QeFTGCVW7vVCdn6jcpp9y06pW/C1wHYe9tF984WLPQYNJi5pxrSw
qu7LPzGFugSd54qeswIOTVyRw0X/0sMeUw7cw1+BObDGHwikctwYsmMhs3rtmGOX
6GpNkQBbHBSDf7xl/wJ+KpkuQJXuc9tKK95behM+G5EfINKz5wfme1C7O263oS7h
wSsMUwojps74/n98ioytAqVHKDSLge975kfSSo3pX+ffD8YPoGEDFMZ4qUaGkhqd
0++vMFupFyuCzcqwW8ntMQZ7GLHhpmsEfbKA1CS6FFgClGjj77//+nGPjanM9zTG
Or4zcY3UvHcuuLPz7Yublzgbw+SL8xB72hhKiZWF0HBuSI+UcNwMjcwBPFywWPlO
0/tZ0n/JxX2H1CUTpXPH4FwCBfuW1ccrk3J1HCuElqo/vd92P3YPlctPNmuDVjqo
FS5fgwizeh2dHhjdLM93o+mfP/r9ZjmZ0Od6uBwuX//MfHa2mzDNPwyvkhMiILtD
YPn139A/77pPqh0a8nwrCUNJ+o7YxYnbXARJ/MR71A95L9jykR3ngqiSFdL53GFw
Tjh5C0LGFXzNLE731V17vrTco8jW6xUqHTi/ZzUT56pQYvFGFVuI3TD9DiY28Flv
ske4z+wft9dETia1IlW6E41NenbZuwBZB3TVhIwrO5D4EBPmQNJrPTWQJHxokcal
gC5DeGcNAa5N1kvfe75tIsmWJxjEXo3kgDBKUoN70kkwtWCWQeXi5fqqTFuTnH2F
yEYoUz3kICf7ZJoO1uEwJWRMo1I2+XZCeDBspSe5S0340EnIlBU9srxjqDglMUTV
G0zzXVwcYJUub3DGFlzk1JE2wXPNxu0gYZhUuTy+qr+UDoPeoriSgtcPz7Wxub2i
d6z7xk/+h89aaoR5ZoBW3n72BtRe1a9rE1aLOs9SWCkqdsKkc6Kfp8dYMbfIRxmI
LUQL/rlQWUGLjtaivB1xYe0WgPQokxPgW8+Dj2cDnrQB18otx5YRDKU0/NIsGJsq
3T0d2l7PunKhE7Dp19aT3qPNOVy6RLSd7NKiiZVxa3PD7dVYPkJpf4rsNVJo3mtj
Ag2L1vao7JWkFxJWBCpvMuuSD7ktBxnMIZT3ill3Xmzg1UfR5u42MEx7O8S4qtCG
3GQJUaqoTbD1quGkpyyWzm8w/rjjk4hKMcsn6fAPzC+4qTxNeCTDsZAVuiAMcL6Y
JR794lfu+wiAgYC9hyZyIjXGEfUVSRNW9XemBJxeiaQhd0KSZPPxK1N0TjdM3pL6
faaqRvHsgK7FtPhu1u3PsIlZIsWPLG2ABV78XfqZaiNqqTf4bRdFb/91ft51lJMy
xtqNJRS3tgIbUgUuj/B+vNU048VLIq9WiltGotOY0a3qynMDxBL1rVbcTOh6N5TY
TcyZTNvjedTTI9H8or1KSJ0hyQo9trVXGiL6izJDe64ObdpEJzvfpG5ITZT7oQJA
Giowrmo1LIwLLkMMunSTYuzjDQfuHZTf4rGZitYBDEfku1y/9FTxHetXs45b/501
3oNLELRi8TCaM0Jw7Ud9nJhTRQIhuJBmSDSm6lDn1184/ArsQEFOwTkzdmM6G64b
PQNdZKQYdhOh0vyH4GmK0t7a/zDclG4nW42Hpw4bMUCfRMEfh38Mm77+ffNqfBQs
b4RCIwXGZPsSSkUUquqKDcd91zBFXt1MtgflJ1isaxVqAO0VZ/g4n3cNw8YGudOn
XFcJ8l7SjV5AGfiyVJA0PCmD/MxsN7mPts8SSMBMhoFa7MZFGyJu/oG26xJJTtA4
hZKCLkMw/euN8nBZMw5+KO4Ncc5oXU54c9j9hoJ8CBsSfxAgiagcBHqSORKV9iX5
oYlBI0JLF43s8520gTCNkzj0/WK6fwlI05m+qQJIzZGRaazB3wpqyvrHFp9TUdl1
FZCBB/qTsK/Zxp0iILbl///Yw7kUGYoMR2ulQn8uAWfKPpI1cIpkST8C9h7Jcfz/
bCK0Ds7kNoCGqBrw19M/XP7ZoSYSxYCbyJOKMkIB4UZ1M0saUvE1tkGclbCMutNY
KDVYx1Thy/xq0ZHA9tXEHITeLwQpWKWj+GEEbRG6F5J4PD51dsDGEwZ5e2M8soY2
XBhvc7pNIuY4I5cxpUWfE81WxvUCLbchp0vnejfHZPhb+W6cgzZ8huXpxbtCzNkA
GMTL+cFf+trezjcpr9sB1pXMDMyCijaYHztnqTOYdP4K+xlUtLoLkKAv3hLv5+JC
3DvfMtzBcuPGHoRlUVgC6Y2Q+KZHsPh55kbtAgYgK//AVWqdoXMUSsk7dHW7mrW3
HprhtuO42nBWQjsjjWMB1yEbPL8vRDD4w0UxsQs3ZO7BG53DWQMwlWjb0CUoecLO
x45r/TV30kz+7XojSqtAH5/7TdQbawybF5LHtgis44Pxqs0nGWjYtSfH+uvBeI1/
WczIJERlRVv8f536nSZPaf1XIxKb40L8VwiYV2mjhrJ3fyFWXCbpoyTOc8111Kca
ce3GDE4da59+tqzUYNrpWbsir9vjpKfteAY769IfD6NgtiuJHcBEerPuIHABwBeF
ZytdLJ8J8jhxMFMK3pSnjJ60t3jUPag+eL//mNjka16nO8Ya1jGjC5KQEM5YGUtT
So6JGZ9g53SqxzkH3gcouUW23t5Fc4//u07h32YtuV5AxKhMMKD9bxEwXGAHOAcX
2krgJf3BdsaeH3CxA28iz9KzbfJOnqw81k4D57cLLI2btP4lVGhkvIkYRzfAEWKN
344rw3yXKIUfRhbtT1XvYn9JnZKHT/RoQNrtcIytSt3khAyOrEuk+yCYPHXrkd/y
JkMx4BJ/46N9MbauI9LKmMyITJR91x3PxbOSh1zaMjO8ONnkSdNOWIjgWPAktHJj
YG2zp0fREHVqKdJ23sfsu5sXh7GTfywuCSYvlgLXRnMS9fpr0B8l9j1hlkh8f/0s
xjJLOVWJZBcZ1y4BIu9bcVbI3McQt3VxO9rC0Ml7iD1RgRL3pamFa3FG0SoSQ1DU
YaqY0GEyOfnmQnSXYCmdY386O3nImRZJNsv186zlNIzn25JwhrI9l+qu4kTtomhw
X7mycVDP8IfzRHNP4+auxOnsXSh9WxJcoowgnQFKeLqpPbZR8WTHw/lnUmsl0rob
RMm5XkD0aONsYhXBJK6ue8bZagkWaT8otXRWdwR1aBVxk6eou3J1czG5UbCkBzWV
muXhMEZ084iXt8ysykeBGRHY8yvmgMpH16N+Wi9kXwbgZTCn9Fkzd93rbI5erkqf
iXVemH4Vjrh/Oerl/1775f8avTJRdmAnD4MQnNECwOr3/wRDmrzeObLvuVxJppKs
QHeyQYYTP+zh80Cg270dNVpWSQkJHRqgdEj8siPb24lgC5bUHFbfuGmbu9Gkv24t
FFf966u9sglE5M3CJ9UMwQISGsXjnL4nHxpZHuU39VYr55GiEcvIV1yWBBsyVeuG
vvgmL47PypxMeeuGjtqGaeaZoMQBWsM8APRpXc11KbDWwck1GCLr2hRaqS8ihDFl
BQ9Gg4mYZuYNoVe1vKfr3SAW9j5pmbJdZ8jbrJUI/1biu9Aeegt3AJvDdcYAlEmu
G59IgK78PVICTTshAykbjZx8QsoQt+Gt4JHOiodtDJNVNELPI6ptc7et/o7sSv10
hbSoOkNQzr1Te5jstFAS81LIdscNHZ8MNsrE+/wx9Iuwy3+mJDGAPd7IBk2CsTP+
BN9uXoIa3Ch0PU/yYjUcYft8xrspq7UebeP6MTCP5sHP4PdEOAnQl40XcjEsdCvl
VFkaSkN7vyceWMz/ls+/60AzWER/Gk8WkvqzKCnZPQ1J+9O2oPl4mZ3ogM//Zuj6
4vrvVsUowPBCJQGH2yVa1NcB/0Gn7h7WD0LMRfFOL0wBmxsnujPxLadlhCp0w9iA
x/vkJkq1hnhjvKBdBWHOpPpLrN2Kw2THYrALspgDWhqoe4cW8nqQ9oUuBMSEVn/b
a3rqhI367cPk07xQZejceVbZ31WgOMCLAhJqfBruXRO7RdE5OkL6BnYvNu+Hm7Vv
n/w5aodhXYPA5CLvoYoQlJ/iW0Wick58esPqkk+ghNZIdUc3FZrKxtZOU+8ItH6U
pV0w5k5FTgpREE0LTqIF7K+NFcoZH94Zd1depQK5z5UsNa4g3hCDJ/56T6HY2tx5
fPOBv9/gPesz7oxPh2s23EN4U944rOhPcF3Ki41bZ243Z1/q2aA4Mx3df9mteNWc
bJz2XofNCMXQfXnGg76wgH/gyLverXpBfhqbwcygx+Fn/IB5QkUZDoMwiQnggkln
AfSMkilOX74PGwP9bGGJ1ZkIqW+hXnpvBIe/PnzoSkETU3w2vxXTfozYXHQXevGT
RPT2W1ZRSsnZbQE/C9WY3rWS2941TtozlApWw2JIWdiv+ln3V/fQx/zY9YYDfnzd
5PWdwpG6SQtT6qYiMkJPjKJJ7bBe9qjpuzP4vXK4IPPbsdkyZi8XMA4LaPIQdxq1
WKTRFJo2MluQ7Ado/s7RY4Pc/OuzEXurhR5/SbSkcoVMGR+OiCg9C5pPH/qOh7MT
i+PjFEdhc2rqdGJy17faRKu3LztNfz4fY20jMKR3vuek8wbblD0z1NXQWK2OKF1Y
f+zi67By4gMDGKepfwySp07p4rUlRwdgJn1M8h4bb+5rrEEi6+KY9id5JVcZyMyd
XNta2W7Fsokj/J3m4cRTOfjfwh58BAiOmSgOBG3+HQVy9yPih/ryyqMRb1iNufkK
rQUJe1F+yVFavZ7wOLos99UiQV5itNFWTn+YcrU61/BI5MvsOkaW10wAmbAp1Dzw
+ECbQ9EL+5K9mVftp8AxJZU1mv6UXQWfMOP0NRqP8kAm055Px3Tb/nURmYHve1Ae
+FPMpeIXxLTqsfLs7iGSPtuSOn/oOrVgKmtu0DsSoSA8uH+F4fHkmMbP11N/ZOxU
myWBJHAY5arn/Yz/EoHbc/tpoJBeUoY2rABtSgwiEmdJF39k5d5LUjdtWTAiWxBL
2Cafzn9EWXfrAadr2259/52o9x/I5YVss1E9cnkO6t9A3WEfTzgAJLX+ilHa3G8d
YUUJKYcUqhtjcxz4bZgDZ6uaga+kEQ5LP/FL+8xzLkRLQzzZv81PLNqERcTbH627
iomyzSHMWeKsdrXPEHKgob5aELxiRm3vKplHP23BTW9JCfu7EdhZjXzmfJhV62y0
V0spsRJ8JbWvhbYqoNJvOnGONUpsNFZEiFr8DEE5L5rquTGqM8l3KgoacPu60AU7
9w9e+i8SJi37uPBgiD4GrS6WhgQ9Z1kkyA4P0BTXTvBwNHn18MAMxlHV0/WxAXiE
Nc51wcVaL6/wV2X9A1rP61t7ImFX4IMUS9LGUGE9+4feD2Z03cXDS0Aop3N9fwek
jbEbrLyM3CY+CJVtTEQU1ujSMwc8U/g4X/1kJuMsdMkYTswldpUwZ9m+LPqo+gqG
mnDd7J2Gn8mhXdVoC2X05BuNpQuFG2UAc5Ajle2fencLEg31ivxVL+LmbUIyyK02
1gZxAWA8FlvYDb+cT+KEfdQmWzZaOYer5BjS+zxTKws/XyDujdXFJJLHmigGsHIH
9MD1gq7onLk6KqWj89ltMTUNWdblooVBbhH/wHoMfw5+7zSMylTMJ6qOo2fII0oD
oW4C/oRebqjhs0g4y21F8baRYTG/GxbTLseGG0zerJw645MLRZRJIU0C41Tz/A/o
oxzVROn9yVwrsHcYDvXoQGqVCa0SrpbIhFgvZ/NxXU3laWeVro8OEKV7+x522591
2+oE6Nth0e43nX8clQA8gEMgzf+IblkqHje63XM6dFn/F6u91ECl8CSOH/BhJrB6
M9qQb+n4oTsJnmGwLdB8vn3M4ywhbmRwG5CxuoXGQ/6qysx7nI2ScuWSgRtByfo9
IpbCWBIFBunARLaY1XtnZvqTNtwL6fRDPKX+Rxn8+DmDX07JiXyJBjruHg2JK/Lp
FA8oSMJsIJ7g0D7QLWBqz9yVjd0D99/RispaAyteSclV7KJdguPrOYtChdTTSToI
OdKA1kF4VMgh8PpxP0DpFlaxVj7kNZNGHSpis0jGeEHy382Oj82GqFIJtcH4ByD3
cyjOLuhvWg8AZroO7edkTI2/eYpnqtpPFBPCAQmhHysSLX/q/TDm6TLiT0F9EZ+s
7uD6SZJ7aEUhnPpaM1F+1DQk26pn54sf/qixQOBElLxKHrcPzoRzNaUfcf56mvsT
mf6cP8U7H3Lqljbh4e1dUi8uoTWcduSlpBf9r45CjuZFXJ3P1sWW+fT9wxoZmsm0
WAHJceVVYo6jLzZ6x300EhsXpWNBbbs8m7SnHfTwU3PfaiSZE3fyPUpv6NtnSDH8
2ALUdSSI2PGAKcsgUKb/nLB8hEbAG2JBG7Se7xCc6Shwn1L9OR0QDfOm72EmEvFp
+bUGU6T6QIHBtasogUT70weeMoHvUaUTrOF9x/zStSv1FUMxlGuNEn2Tmn/IN5l9
USEF2zsXkcZMKn6HuPEThkIXE9E+Ra0WrZD5K5CHyTjway7KQWNWldfhGj9hq7DU
szkf71bl9BDEIJnUoyqCT8xd6A7L8KSJUPgXgcUob3IaloiSnPol2QOEwvfP3dwK
bsNvGEtu6dz2bcrCGrBWTXb9F0ItaMIaBVhQIhsJdmPAR/xNxlECzjnc0far8dYl
b0Y3NDdunM9AopccB864oM2iQl9m9PhgUjAkwc422mDQGTBTd30D/gBBpQ4jeEvy
QcRGSEEnzBAmX6sSV06KgTy59w3CaM1q3RN4zl4Pzi1KtGmqJcczdycpfuAiSiRe
cHucNOZYBKzCpAdaaAFL08InbvGHd+VjJcUnwjncVTpubfStJpFKzQpbjiFevahv
2Hd4R+3BfiRlvtoqjOHeTksbqBEOkhqMxVlQ6HaE6yvjrQHV8gtvnhEKNm7z0ZFY
9/FZjetHOwbtVAZfkl6IFHeqQ2tSX6yDpsZul3i1eP5kvwerqu+uSfba9ORbnL9n
4oG31LjwGExEsUPGdP/YiDoITHS5okh5jyzXt9pBaMSkfr2DZ5eA31Al7yilpCSI
k4czfWxJwH62F1em7+++gqVkt6WkhGgBRTT9UdBjqfZuZAUVxgGgjQ099lrQOkz/
WJCZUKM6+1YDdb/T7SVshLWRFFXoYHAFKC3F2hfxiJtwtOXqvuaA0tZf7UNSamj9
WjJxGezkQlcWTr2jWL5TdDZyXCBgRLx6Je5CzzhSCht5RFuCkJ0H3D32k8MCxV0/
y77TGtA5op4qJgv8nAkbMGyeqgXfx7PJn1vixKweRXWIU2e12R5lNLzAdR221rYG
QNinskZD3E48G3jiZUs8bPUq5E6QhLMifSd3u2ahKEl8UbgHoZf3mGLKp6JKeS4q
eGH0wgg2ZgVKcbvMxKbWg0GBh74Ay24Qq48AoLGFPML1mC8bCTvlgCp8qmIoo81+
1dhVw9xX/qmi7BaEgEY+smO5VcQrj5jT/m+1z/hFhm22V4lJl/e0X/JffoCKmJJ/
8vNjXcqAG9fYUeY2NmMnTeeBgTt/ZY1U4K724ImVfSDnDoQnDCsWeVKNJrSAWJso
DqR58rIuGIkZT8jMvH/JVoK8hokp74NrdYvVHRax7C4K1sjepDteH7RUj8asDU4L
aTUptMNHHCyxONn++yjcPB5BFuChCwYrdgJ3gnPNsMjJX45NFrbQw8721aZxp/0J
eIMVX5l7CO2mVO+pb9UrhkRDJFyvCXj9xc5iV3ybjfDk5w8Nh8jEUOrouIbZhxRp
3ySU9KWgQTyishJ3FpqYqnQn34thslGCoS5luDaIoo0H6fRkCLUQnRFH9DA4FBmm
qSRFHFqiZxsS+E8zGpC1hJXniuaaMWPsVOX9INe4gPMvBymdSU9skIuMebqylJpm
J06G0c+wPE3eZlxxjGpueDjda7HndbS6OLlLKzoIqrxo9ZBZ0ddIxtGMI2DA4KNP
L68DliC8w7VIxX8Vswg0LIf2NXuKrLUrP7lDr+XJAE8vMAukncSLSGmXuybXyi/j
2w9NQAZUkf/E9/VdppV6yB9cohG0kM1j+ggEBTtroUsKk1GCBHGBWl2X8veDRxh4
mftTQpVDS26a9RQFUUoqRCAx30kkgKgdV71pQywaMTSb/IavmlgyEzqY+0LJiOvJ
tWAd88fY4m4O7LEejU55lgUomzD5LpRdYmnzAwiKtLex+hKRooDwconDiUB7nwUk
HCC2y3BCH2OSQwQl2H68vBFfGD1mS1OBAllTg16xMjiXPh7xfjSi792ofkxnXjb/
RkhAoqR3WxrmWUpSEXKQeoCpN/jn7LqGgafZiFQ4HVVRmMgTvZrttyG7pYcWEH4a
cjajdzWKwNSNXuGDm3fPVJgX2vDKEJns5xe5tM6NXAeSehq0XmyEtRMsScuyYEvE
5G6dRYTJfFUY6WbQBb/eK8Q/c+oWTOT+ndHLLvO8n3Ra1nTsaSj7mqwDGwCzpwYI
9cdewzg+G3PwtFKhqR2GjfMsfs7QK60daFaYCCm8Ew6F8AC26mZJ8MeUlaH7ayaR
j5DdcZ/YoNwFmRtGUG7anzxsSzzcvqdkPw1SB3QjOvpZgR58RN9CgJAPjMFaAH/L
l7RC5yfGwGrSHHpuZVEFO6hOOJ97kFEYvkrhTbw7dcxtJEDBjxodsLw2Tyaq8E+z
dN+4d2TcBoS+F/1IRjv/nM1cri6953h3DrHV2QM6NMNXltkxLg/aR8+0YqDDjZD0
ohTMeXsnXs8AWHEHj8mz6rrBBhpg7rufh+uR/K4iUFwMywju8WDn8AvZD6Y9hyHu
cFIfqQ824Wj3FVJQGaB3KtZnGD7+kf2dNC1KSPDYmFlC9DiUfIzAx14pQhGFZEGi
3M5GyCgheiq2qJXg9k9AN1+lPLt4aBJ5DPLYJ9GNp3ZOdsgLh4vu04eV0JU5Wwvf
GFIJAZraqQ/kD6w95LCJlJDsMPhm47xNvyNRpgEornibVROoUIxvqhhfcvf37Hvt
2pZf40Y9j4X6NYajz/VB8zTHxgYyFu+Bvmu7IQDiv/BH0VO+T5iuitKCFj/01fKf
153JpQPTf+efjvfa8an0v68XMqrq22t5XLOvsJX0pqN4Tu83BMzIwWHvXQw9I2L4
qp7sCxLFNG2eQmQ1cg9sLyoZqUGsmybmj3W0kbwSFcayq8yshQEH5V2evpnXOjr+
KVw2Fq7YWpYuKyIz6YM5975o1sD+EB1nODFHfyK0/syqEMaHXhjzdi87Yne1JXyQ
QxZ3pKI/44Xbwbj/0lI22Gok7M7zXXZ9K7fH0j1N0MqaS9VfWYrryH44MOE7wv/l
huvMHeZv9HtuQpwJAfmflv9M1GJ4cDSJaYPvvTqItv9kdbqssS7GxG0MMVoNXqhw
0VYhawpf80co7ReH2sQzdnmDTJ0MTJY+bJK3sV0MZzMX96cI59GBFKdSpiTjixyK
ScxuLYjhY5l4MRIz9EhDbWYMcmxnCn0N4Uxagq3iGNRmOQGjmcgkRQ8X2DjU5e4t
dGwGSfIyQcQpqtEpqiOf0cjCfmaGGtlDCiw4vZjZ9BYXP3iWo9VADgcu1QjAIbv5
rSjORAgbTfnuNe6V8S6bw6+/4PUsp1uvZpjSZFjnf6hIBZsujipOB/8w5M2gX/mD
PP1SXAkInK9X93GOW8xZJupUJS1vQGk0VWAmhtfXB0/GrnYO4HNeOuuxlQolMYIE
DxGnNhs+B737M+RzGEV7NCkY0rDfJ5DJ+IJduBnU6WTQr0u/A7tq3IIDlI/rgsyh
VrT5LZXtGu8/Q7Kxw+ZMNpo1ZJHHebLDNAjfQmU9IRaKtyhPAm9tfoc9JFtE3rFw
qB5+v/UW/wQE5JyHvySlTmH7HSrB89Kc+FyWNwacYnk6Ajvk3ibck3tVttHig9Vj
vMRiHMyrkPkXEO4leWOmc+roU6E7oYqaKnAXGw+9eD5Nm52SCOqBlfUoZ1MFxdZW
E9BeU6qp2O14brN109fPPkE6rPqrtNzEQ+u++iT2cX49d7MWeKPFBP9YeozKTm4L
0LVHgcr9UMA/vQ4vhHRL3WNoCRHz6kZUY2j/+n8ioxIBZRyktsV6MKn0g53Nct2T
c3gfQSCMt4bXnaOZOOM0IbOdYkHb6W3c7WMHWf/EbiudAHdox49+MEZtRRGPCE5N
Xj2AXpz0x+xiVJ+g59h3x805cRPUpA84a9MB1wf4E3cu80DgCuQ0RDrgqfXWrwYW
WpVUxQGxFilV0eH59vq65qtoalJHcF9OSiC1h2a5R/QnWnt1lp/SzIJVFsYkeBFP
hUUh0012vNvXVi/KB0Qoae4P8t3LgzIva/AnFk3MBuiSJdaLpTq/p7yCK6gloCFp
UYhtma4N1qAkoeulHdIbAUwiHAm7IR62t9/jq1a3LrM/QBOTLheuNdxc6lWMoVFO
G8ViTWrACER3SexMsarMFvgo6CrsmqhpxAdn9gA5/fQdP87lyn6j3X4TG/M1fjPH
Yd/ZHbsvgPppIuZZ8r+6UiB+ocmkJUOhcDTcBFZCtPFif+gLnBQY4lfPq7wNozrQ
ZEc/acqro1QPQ/njQzfZaZSdNzZoCuQWi3haZ0p7BTUPkHAq057hq1STpTyvwhfB
LTaQEnFYOJS1FZsrZ+n1u94pn6iKbvrS06jDhf1WOEl5X4uOxCLfQFjE1L6Nx8wx
0rUctmKQZRG1ulOz0tABvlEmu/Khov6HqQp4Klr1YcKIKf97ZbOMPQoqQkX0PG90
hCJgowWfFH/ZRAZCGNdjngCSP4DV76YGT63qaz6iTOb9zMLttZP7HRZmpzhjDchk
t7SoOXSXK/acVKB0Y/gzsQeGloo/wqlOBWHEES17DEm+39Xxdl5HSfoNZ0dUQptb
L2A37MuqodcDiiGR+sXHpgr+sH5OUtxKnPTvTxnH6aX/IXTF2EnJP2+HlK2vBvUD
+OVTFqptYZwZ463E9YzRWz0zKs8UQhSsHPbXO6x8+/ytEr/Mh/1tHkw+YRjB/ti8
lEq2Fg4e1053Udw8HVazYndCfgIdzCRg1WZ1moKXXihU+N28byp4qR51yUbvR4Fc
2pMfjmmbzz8WZhckAvXvkyPecCjBiX7suOVNUXWuzuaFKbc+7GkFFtBTddkDv5WG
JgYH4+7E7wy9QCkLstD3P1fWxvci6TC5CGgcEHAqryacxyDbOflkTuT6CCHkJpmC
NH4/e76Mk6iYwUumE9HE1jluvaYUkskCCIzXRhoPDxKZLyQr2Nb+EPVJK5JLvqCG
EW4UtCJ4ml8BcAnb+C4sEN4rmMsae22zMkTVfKgS0RrL7c+Y60fG/MF3w6kXb/VX
ZSbVzVKSaA29TsZCHlw+zrDPCmab7pkISmMMu73t29xziLtm/WKkivMGMVPt0N7R
A77h2O/VXDVQarp43labRjhe+TzEbDH7toEKdYA4gOuodoR1PChBNvy1pb1Ufyo3
BWh+bwmMzs38bTrVbdXZUquoyYwiTc7/lY/zNryjcwWor0oki1BAlwZHf/vQtWVI
bEhe4VnT00SojUoMPR9rTMrRPIJlA/tCJLZ1/daAh2WGkrWPBU4PJJgACjLgSi1F
gzlrgHrgZNq00g49jJIdoZolxzEhTFV8q63IPEMEEf/Wi20MeGUU23AoStg89Nbq
EmGmYeTjqIzjbO9DD9XSuxTpp+9N05P4G8MJySs3ZU6nxXSW/PKIWXcrYVPjbrhS
dM+N0ekf3jyrOrIk3JWhX5gr+Eko+aOVClXTf+bGDlawb1+T8Z1YMQJP0OmfzWGu
v2xS4m+gJucvYRvqPB5cyHLaCxo5YgSpVDfzxsSI/wp/E/Lv4epfUt5DXfbd6GJH
5ZvU96Ou9tPSDpVvdlCvJTiaUXMYUC+Z/PEgxmBZT675xGGnxHDzlfDkR8KaZx0U
zKue1UXDODP70aBTHoVQFFBwM6bXMCs6+iRDKYUSxatxKMpBYl9yrpcfpU1HbJIm
nSa7FhYk1uT26eD4/XtK/XU9+VI/pvxOCp5GZdzMiriScDW3+a7pX6SsPZskIfYE
afgTNZBee+K6STjKBeQhNej6v88m3L3bB0AyfrJ2LfYv/LfEPfpw0QLf7LSie9VA
Hef2laP4oDTqv4AW2ydv7DRakk5/wR82IhHo/PwvDqjvTeoubB8WBSddBzfWk6Kk
se61efylTTMnicjuv9t2/p+j9ZBeh3ouxJc5RmpVcsqIs9jtcSJg73TwNSr7i2FQ
8YikxoxsbehVquSTdlXLYISDC4T/dfSqw1wn3C3dPpHmKDQ2QOFWZsrzmA7B69sC
vfnCgPyCsw2UtZkbFeeAwwxdOJGiOM6oWSDKrdIu7SJSpFClSPI5ySO3gyKV9E33
FAzzVA0TSYGMcbve/O4enLs/yWnkAO+QG1DwsKf5rbZNBVrHcfSZCCT+iDv2TaCp
Yh1K3miTDIhkEFR65qwl9eTTXspgxGmGlNXP4awZKcyD3BLyquN0wsktPiVirYL2
WdSjg5dJ7R4IF8nc9Ad0hI4iKo55kOUnMdx4k0o+khiqCWSxL24uL/lab/rbaG8I
BibERT0PEpXUAXBkkOTD5dAaIFyvsMupWUMhGh5v2so7keOgZcJIrSmvM+2qTqjc
xGGKG/09pbGFPxzYNICuOOJZHaYb3iN+fOuSltluD2yk8lBHi9hDwcR+if7KGCj5
t4oAIo7BbtHK12hHNWK2UrwGW4lSmJJctfKxAt7GrDoZ9k/pdQgz+jTvXm1J/2Q7
DFmXb89E8yfDAhLmIxawm8ebzvhrAvHGrs0o37KsR7k5DMDUf4VifSHKDeNMzImr
Pu1pp/BXEUVWbTUfMhxAq7Vk3WrRdREYlVIaF84jIZGDK3vErJzUv7sz+//revXS
bHqMBf8a3F8fiVazxFpsjSu1/+KC5z4ms40aZGh8vS7A9WcyWvMAOjBvPHXAuGxE
PsW3CWB4YsMfq4nCl8Dujx+9gWz0jhA/OfogF2Lt2D2yDmZsppESfIk3aK/wqmQq
bdDI2IHopIV97xiA7Sg01aISc79BI+TBsbtjPpqW5bgq/2G14RVp6KYoqBk6sobW
9s35ivu97mjIchZ65b0TohmIVazQOTnwv9W55ATZM7VVMmtDD24b2z6LngdJBHuj
C9rzF2rFC4ErSz66b9uWsdzsi4ErH0dSm3YPKwH3zdNBrDecA/0FplGft04l7QKz
PNFC2ZJjF9Y4OecBppARbfVhugKHhxF6kkmZJvmW7PRESDF1DdgbTrDu1fdaum1K
cEQUjGIlTA1I+uOCqMIAf5XVEwWDUyWW8Vs2y1ssb+lWzyKVx8kyiu87yy8GN0gR
O7tsYglVs4RKlq9JAQqVndaqBQXiKTCqSQdzka+RkFC2+RJvBDIbXQ/0IfGs45Mz
G8zAfmKtgmDOnO7yTaN+PJvvNiC1edIQB7M97ZVN2W0dFVe2nYOxV89ocXujpE8+
hY4X40fh2EitT+g7FKzeMkpGpnrAZD2LdMTCjPztsiwNaLZ2T8/bqZQ8XCI8z48N
pbUTRDV+mcKmkfSH0y8HIj2vwZ/6YGrl9rdZI3WFLpZeyICew4YgQiJ3XEkQXKTG
bD8Dzc/WcC/OZtzAvyVRyxOysGRwH3MP2oPF2YQsp3COTjWg4yneVQi0m8UJHGV0
ej67fKJ/mObeF3pCJrDuA6XUFbTBiAj5iDzPXGQVM7x9MBNKdJ6C53YEOnMNzdOF
am1Zr1pvj8OYGgR+rfGeYw53TSPJsbHaUmV2KrTIuwgN/kev73JLSMjfWzp03Qth
+3wjnIAahdWpRsSPdcp1M0HX8l8fnWihECkMtbKGWT7PSYZHjq5CDwouefPTlT9S
+l4SatBMWE/cQUVnk46YV5hBKtj8GxrODpPJWAQVJcyC8VKMzd/5FlGtrIW3g2zT
CU/9aEf/7iNj40JQRkZd7f4yPtmTZdfb730hHQRG/hpbTgldgqhDqsbYZyDdrim7
2zt2asCNF2O8GkBBX0NWGy34pB/woQY7hQAg0liWMxv4bCeOSvS5cmT3Pr+vyG+7
EsxT+Ug/a0/RtI4Q1qNpjMLZE6DtYsoTvOpArL1rnOMMHp2+1dNBjF/ZgWWLGaP8
3gmMYmI3Ld8XoPi3CNSR+a0Jy6QBEf9SyiebQ1ziUZ9xAi5+7VtrHCIa8nwCIz0z
YT7VJ8NsfEFPYZCVzJrly0afXOCLCEjn72C0kr4Cf0g04NsZS+feRtURNjcanFpV
ju6U+KAdLVOYbckdPtSwHtwKInVkCjTjdh1Hgr0T457wBtF9Tchqn/DHaWUnWNfG
sjF4xTp4XJ86AIx8UWmBlezQ1jU5GVpgOlBWxb60MozP6Qu5wP7zS99qSZOpeh6M
jx2dz2dFQ0wYlQ0VIifb++y07JvxwiW77rx9Gwm1GyX1ni4/NCUsy3jp+qDtkwuU
CXydNEwnvc2bZIwJYeG6RB87wH+kaNZ8ScMa0cE/0bwjxwXiy7nDkA2FRJiptccc
A/Qe5rtVrDXo1FAzoQ1jeRIhnNyIvDmpeP20D4acbxkPKFl2ME5SGvfJvLG6I5FH
2QqzZVE5/LVFKSbFyjaaskagZHi924DJ0N3g882QGjDaNS2pyoplf9V9GcQwUNoC
esao0jL/EKjskrL3Lkrqvtp0DVdFQCGwSKYH11aoIMQ48B5dz3oy12poraYt4J7V
ZqjkcYwvXNb0B2lyNrHQo0DN4a6mLC1ASho54yACvW6AiV4qHPF6xs3g7/kDfDVK
U87PSRnPUZRXWu9U87Am82BYDflehneJsyR0AoX05pl29ztWsDbbagQCUy/UhkSb
LnUlHbmESuAFQwY7noI3brYvlh5kOZ9Neo0OfMTP/u6jGtRdlq9a2mPoPc2uZmTY
77xrTMBHyJadSSkf6d23AYf0yiv7GCyT+nkcKr/ecd7pH4QSg4B96RT11F30mmM3
r6Vu5uBBRe0ZD0sGwAO0TrMIY3G4MW77A5yS8KcIlRg5GlbfYoTKK8NWga62LPPb
So+aZxnlLiUcvK/tQtG9VGM77kD68Q5v5zbisb+aSgymR084v7BNJyDjdriQAMfi
ZX5SObOy0Gzuq76DQIm2mj0wLgdkPC5VGCcjHWTvLB+ni2AYAI+uFxbJWuIgfyU5
K7Ih6QqS9XmlQa5XGwS+SrBPab9hHNv55lk+9e4XUOiD9pM16Ev0wQGjqKC6Elxz
8dSyXOyu+r6XpCZYlb2961d2lvOMtDPDh22o6Um1f6XDAEHIxki4BnmHy53abVbL
0KvzhdlGFYhlvtOHmst+PJwb6zZchNmLvL6tQAL/iXV0bE7SPpgOLQ/pQ7VoqdOT
p9gIjwICGKPN+Pzlp5L69wQbKRyLeRlx8h106Dsm9Q0ZOvFgNYSeRcDNzEWuaFXC
pJkmVzRgFusDTGFoXNUJNjmO6HtfG65OMs8Jbj/gqz8hH4jwAJvoanVCYnDl5Q3B
2cQ6hI47MpUk3QSll+hKgDGzYQ2d/5+ucIeoeOS1IVVdsUJs4q1ul0zNxz7G7b6J
9tNz/3l7GITo2hwIk193RqGpyz6C16OeIKk2usf33pGepCwDmLkwxml+63W1j7yV
PjMzWqtNwu2Uz7utFeVFFBZIQq3O2yrQxnKgMhUjU5PvgcYHOOdkjXCj+jOt4gq6
Djgw/h4fFsEMdei+itE7mnKWoz7GCbY3LD+FW8sIVOi6mPDGZEd9FgYqWePG1arB
ZF/kKebJu+m0XgoMSp3h5w4ZqDUhjftgd150/5s0FbeAFb0Qihsu7VeEIdTxchUq
aDBv1bu3S2VnAwreHRm8TkpLuyIEndBDALu6NdvW+SWB7h+IlTlpb7JjLqC9Luw6
Q9GKS9MDQf6vqpzed0Yvt+dI3chZrTu9w1SfRcse0+lHSpb46Z2ldqfCskx2K9Hs
cMaw4ssPXNNfcUP0tDlfj1xiCThd/VSHairJ1EUoqPME7cn+Ja0rqDjZX/RL8Zm1
+4WWwOPMvwEld+fBE07YecGhXywRtVusNZrT3L/RZg81A+QCb83uKYbGBYGo8zIe
d20pUPiBNl4FZXD1nh/M2dei39PL1IaZQ9erc99j7MJizxucs9y8zpSWWYeNMVDc
Z+FbsI9qEFIkBpltlJflhz7FaD3SDHN4W7s3wvuke+7Tb+X4DqaDnvh53JBny1/3
izt7LFPhStnZpSV4KsHsfd2OnyN0AkQMq4qBZellFoIjqXx8eJ/vWnDYt32fcr2X
Wc2FIjItMDJDH+s+pV4vLvQTKnBBxJgoZk6w0+aSaGov2ZhMrzP0ZO8f9x9riU0l
tX81Zt1KJvVxXrzSOxTijBV2ARrdak3BXZOMA6rAe98El5+tqLo06TU390NeKONg
MTcXK75EmYJZuh8bfg7U1/Dp2wd5r/QzqxMCnzZ2e3hzf5CDwz3f3KiaVIbzhUVT
/luRz3ua7BKul6qR0oNUW47HD/WVmDEu48RDO1Ichrrp7RBQFTKrWEwT/HhAZbwM
KcpHe5uFvk5GTqzUo6P3FHXoPhTgK8WkigW8CKKcwn8XMnJeozvcoYR+pcB2EAB0
qn/gXD5418YgBQFFVzNIQItgkOPIQbBblFyE5aPa2XLAmeTD+6lH29qMhDKIpgbw
2dDzG4r5q5xZCWW9639BaIqbmWbulZTTz7vnzQy2SjQCl7YtoKc0SCVg9b9CJaeU
vvfuXw5iCm7xn623OefKKIfp6ShCse0bcXTKzfVUWacTGB284jXobd0rwA7qKMnQ
OftSjAC7zmW2JGQ3V1S4m5ExdXAPDd/0eR/OMdEReE1vQ4tZPJ746k8FfuOZRGcd
5Cv3rT9+j0o1yK2o5vB9vRsdrMeNuDS4e24zBaa09eZ8g2z24K0+/70UoNaaZz5o
1AZ7w+OthJL1ukgBJ5QPu28c89rA1GlhlguE8CeIExbbnTngCH16HTF2esjI4Lkk
n0y64eEHioDiI4Wf8AcB0X5U19hSewdpyPwVElvuc8cbcPaS061G0dROH4Y2bc+c
mSzDXPXIMUdh3BOnUXvtyhe87ZnWhVTFj021j2J5jtnlW4INdsBeuABWMa44C+fK
LS/ZTug0VGzPhjLKrWVzJsSIwmxBzs9DOwpnnMI5XvBcFt2Bds0NWeR7AkFEOFSw
5B3nKZRm4akmEzfCeN4as3xj6dHI8BqSyQ1R8B47RBSJ8Ok82W1NKcjwl5ZHEI6Y
+ll+kp5HU0BFExiPnfDY7m4ZniBjkH9Sj+Y4y3Zhm70ON6oo0kPBBxfakJ0dhKXP
DQ4v/5GKVGkU2EyWqxGKvB4+ONt1L/YyfA2Ok43nB8I/yGyxc8XZ8zn/jW+2bx1J
8f7sipVXt0HcPPErFAb/lny5Ot03nHZdlXILg6+mFnJJM61OV5mJIK7R4dr3jVaF
V/jFjV+x9MdOW1BwK3LhH9C+cGw436afkrZgt9v1CgqSkE6Tq43JXehaB9Z+D4F8
KNkNuAHu5t5GkDgbckb+VQSgZ1qpYiCLOm4SxaFPtuxEqI7HbnHwdXfp+XPC4TVu
6UTxeYMusGs3z7sjOBdNmM2U075KEm95g6BQxehY8Je18HgI5GRLF/e5YSenDpW7
WIhv0sKk0TtjhiMDFS3TnDqvuz6QuZfA438P309kDcP25mi1rYDeyylIk70w0X11
6OQv+Szd6GRz/X0z/+xdJTIp1yhQraEnn88K6yW7Gq4dGOQ6kHHwQ642o2OUD4KL
uHrFocmDxHZd50Zggu9kl1vFcJpNRheoQfNJuhZ7+2Zc+zJCwPDTXB3aUyk1MC5O
jRebiMIt0bmByJi0+AAvgn/qkEvOn0nb8Qp6LxHilSJoM9Lw+E0a4STD+gw8emUI
cH9x7M/AcxacocHvVPIUVJKy1ygL9r5oCq2LLdk5kldu5O0N3AhO+bQ9ztbWRT8M
CJcnUiDbAWDXVpY/EjfKAnFUwWiWjRQ+M02e0yTixnbY9YhQl/+pN7xI8E4qQqt7
Jb2buHyoZiyWYXHu96BjroDUukDG5sYLR6cTrR9UinM+Ctp37uRxPe4pTh6TpwRi
QpOQH6GXNBGbediX2DRydfM5UqE4NDah1Qtgp/CJpKIRr8Ss9rOSmXeRVzOh2djm
oAq/iBB+zqm5SUDheEcgHcTpgSWfrNle0/kWeha6QGUz8hAf2BbgshwhIugp8beh
RkrfzGR6RN2BCrcIlr0O5feAquh+bsK0E2CYIAdldCBWkrUTxwoJCCXRTd3DUB/0
mafJruI5CFV3q3Yqin7n/+jfYhqQHyRhJB7w97kWKvunn4MRt5k5qKvt+H30epc/
PW1OiD7a76golZajBZYL6/jmUxi5BzjrQs2vSEwQF3ziXcuJelR8IRq3QuzWt6Db
b64mx7xv8D22y2G3tg8gF9ipWVdRkkn3saDj+rWAFaZrW3lbG1t+ZrhDsCmUtWa1
QH6iBx9MP0WDfWEZQQI7/jtSscXB1AJZEg5YK/3JhrrpBKJmnJ2nFBcyb29x9BAr
RS95xjJY3iGJL9VvI7dcVkQDjSD95jtFJEP8pZgCV7av2sGqXGCg+jp/iioz+bw3
7+lOaWnjh3ktjjaO/4UmuOz61aK+HYtpDpgLpidouvYOakY5w+19FwjAq/yfrIJ8
+aIAqo4PU6xB8mKlYlzAalfPo5Y2koARf3+dpzQLD8t0yZ72sNGscG0NYwd5yTRs
nRZcwmTA50IPW/tOzQl/7f/RPq4puNOM1iAa7Un1l7UX2EYIhzpGr7UssBrA6nt7
UjcnZmjSMyfJV1Ze+L6vi2su2xTNLPeWYR55I+CGmnlLQIBz+9L4IhwgDHt8k7+t
akjBWw+O3jenYEg73ztMO9/Z7CM/oa16uHvVYL3IayT8zO1wqsVTXtbO4mhxNowc
0AeSF+bLuUJJkmvrBhmwtf1aGWYJUHEtCSuEVBBVlpfeDd98uI7IOqE8yybL9FZg
pKO5QoXlNZFttcTdZ7jJdUetkicAHPa1rjj8uWz8zKZe42gX6bU7QokjrK2aYITT
LNjJFhAGqxM8OayQUr7zEBL8J0gf+n+GP2lEn+u2CiOvUjpEBWi/gXp5EUf9Ok5o
OKWYwE9EqinHVaKena9w7aWZCqsXM+3lr30Ri83PP+3ckYS3lQ/r+o4uXIQRoPXJ
2CUQgmIiNUSyMauiIT09GSbhAikotF9JaW59valtaaQPPsgG5uVqxllokQqxVQsO
+pvryGhNeUg1IAbPhcpewXgWIUkpdTj+tAS+CexnCMCItVE1lI2fC/Ab4tqierhe
clahAYFkOTmHHGbZARReuc5NAduMVAWXSekXF0G2xhPcEcgX1ymaVstcPq8Od9oE
UvwBlR8DbuxkLB7rtSaPj28ZRdBVpfFgXtLnEjg7ykHiSTQUDgsI0ndYhaMWPUEo
eTrmy0AQatyo0qA0fyZnlZNmTCueFmiHg4orf/5E77WnojwNH0HFXcM0wXlMJxLr
EoJNuUDDCJSLH2hZHXwfqjrrmgGm8M4n1m456hEi+f2vhcO/NVtJDsmYeGU8hKXj
j7lVvyKqWIoRcFKSxv4p0wra6uP74pZ83mse+lf540O/ImRyw3O4/kzeZR57Ezi6
zPgQX0MRok2Vor0WEqFWPJZ6WBxGXVPHMCTH42Y5I3vj5YZPwc73JzLDkuDVfp9s
eIS94r3/rMVWuxyaJ08sIwYz7N4s74g8M6GIxoSKn/OeFLHSAW052I4257vFG6BZ
MxgqI3aqEsv9DbZtIBrsIzJhBO5/eMdWLpFdg9qxJq6Y8QyF4DYhaR3vIdufHJ7w
qsemgrcHSixfTqfqHb4bOoCK9M3ZzYYq7ncleMB0jIxJK7ONSmIr5fHj88bNUgJt
RepAaialEHa3EzZruI6C3ft4jLy3BlEP8Fi4+Hg62lscgyo3G1YFh+n6tQml0FdN
SdZ3cV455sx/eB24KEMr6d7b2Pm3sZv3yVZxECuM0Bd/5u45fpBda82QM92ABm/D
92GKbbwcMVs6zfO2ZinAloRFKVCMURwBVkX7XsZZcjq3+HKz/6C3F+dQ5mjCWsNH
ChMOrVmPikqZYTXrsaUhtd++dFEZutzwOumcZV6dQcL5S3KXB6hX46ZEFJH6nBJ8
2dGxe6PGdCGWQkzkYJQ5npBK41ynanjYfgCIOKOTAiJKlskW7Hzt+MVIx8k+0r3u
E4d0M9dHSan5T4Trr9sB3vd3jP5/d3WnmVXqkE95lX3yZXf98f+nWyYk0GFWyowS
zlyOP2QgH3o1bOPJou1yYZIZSA0HgVtS36JrKtgis3VPrC29Fag+wBOT2dMsTs2F
UVJMAXjhK/STxGnosGTca9TI9B8zo23ypUHXU03COOeX2QxqO/ZYRVbEv1GnFLsr
fScLLZFtzFxG7MStDeYq3WuTeHDMkqX6YE4CUQ74KjrW93mCSNrcDzy9wJgSrKlS
CbmJaZtxHJqcgOoR5FxlajbR6syxywJ7bV1KBkh+TrxQXKSuIg35vVSI9o6mMRPK
iDLkzQF+LXSlahIGLYH/kL0oYmj8t0k+qRBHIPYz01h4R3bo+cxzJXKk/0otfkO2
wp6tjMd/sQffyqRLGdeffNG50k/OYqUmHjsvN1x8BbNtZv/J6nmc/bvDjF1tZQpu
oYwlaOmC89PoZEOBfCBKsij0yMEK3ZXRk+BIkdiJxbD4KGmpAoFMuurWzUgBjIzQ
is4U2zJHew7VypwnTXWqul1mtdR1g5XJXb6NfdIq93XzTV+tytMg2J2y9DrsZFAW
TlBcIyMkCkYVM7tf+6ckIFvN/RGZMtE5PlFvnXD4OozzIzL1gy9cODPWYYHGOIyh
j7/mO/r2Il+cR7Nzqyl/1fhTwyBtVKw/9Ny99MkKu55KUgxFYBHxWqpRnB2+ijRi
r/rrMDWCnmm9lqKzlWgPxTiq0sbF6O7PvZaEF3BFGCmBA0Uo3iQyh5estBF8/chx
Cqru6ozVjFGht44E4fjYkE3yGKWiQJb2eWtIsZJKlvNMgdNWm7jeIb0MvE5ky0PE
Tpo+UyGYb3ym/4tGCK3eTsvi44ye7cXZp0C9qtHK8ALdXOft432ZppgdFI0zoH1i
JJnBh4wkQNokaDfTUE29P2eY87dticuxe/hlmFd8T+8++08kO9lp1RbnFR+clMID
eggwzO27oUalJq3VnTL8Wrsfhf6j8H2WieIFtc9FwLbF2TCEzJ9Ok0XiGgyiM4+j
Fl69hkScFDpsmABXTN60B2Gu6asppAIsYB70W92dQk4HG/+DeMkHSodf1QekXAjT
K/YRg8sAzWI1WEVqJH5vI0PQ+kO4mGX7+pvlb8qPlrVsn6TPW9B4hz/WoovWHBUx
IORjBjVXscQx6S/ASnw9rJ9pf53lP7L+Pr4Q1v2QFFaPZkpe6fSrdj1hUI8v5y/r
DD9wS3l4jQQ1KfycuZ9UKeqAL6+l9GchGwSA/TDY+ZLaSAXbe5cTUA+HQKFVCyet
4sHIezaQQD8hsD2FqL1PrJ8qWTOXFQvD94/h1grTlOsYxsdlEQE+cApOAyYjX8ES
7SiHyg2lhJ/D+g3Aq/lqP/25kIchDMy3ThS54HS/U1VX/SgJW+VtIYB91EcMUyCT
R4dPrZjIRXmvV8ucToxdCunqy4v6w32xXk1nUk0NlmGL/06YuH0vSRG6sRRSJ0dQ
QuZdKWA2qYVo0yxqsTKyBe60FJ8O1qfLga1J06TS/zND7rLJ3aG4g2maF69SOMNB
0+bSht42PiccqG0aR2ZWn8SqTVjx+gri3iiys7VCqUtDjDVRncSw4+urSU/a82YM
z4+uIZ5n4wNNoJa82+88htf1arFIOtD0bYFkft9fzYipPyIK9Tgx6eY8fr9q8ECv
h9m54qguVNKPcKJKYE6c27tXgb5m+cw4AJ2kj1UIq9xIFvLqUZ3b8YHbCbU7/3Z/
LIJBzShsYHn8W7hQjxtAYjwcJolk4+LxJnUyhr1hSmTx2yHHzDlwxXT5Mno4IpxP
UNlTy5slye9j9qt1SJzA+i4DdP6Xg0IQC8IsjciKHN0WvL8E1xfmHtHk9CZmdFMC
xx/YWpjrnsHIsU9N86O/KUEyPL4BZG6uEc9LI3v7tdWW9KdQqldizE3X2uSBFtdO
AV6jmxM9Tcv9n0uN+ST37OdL+HGGNKAy2fvqlHDGqR1UFSQlpvRS60IkrpWe1dAV
jXOdYpeSQ/CsRfKPOzRJwRnLJTsa7/+85XREpYTE2Mif9PGOuvX7mRB4iiNsRpWH
lV+7l5JKWwN7+BzJ9d3cmaJ/pb1E0TBlg8etmaeW8iyzlM1bHJsZH4tae/+zQCzE
OeochNiD4c9oaIZbtb8zUD7B03YU9huTJOdJ2vwiBoALIDeqTWXn7/YXAxOeOVIB
MnEkbOjTLQ4khquKC4BwhP4k5R/P+zoMKThL5YNfVQ1KCGotHryBTZnds2+0V0py
9In6/7g0rtxASHSc9ERJL7WB3XvENKWLdoblP9PjZMTvbJSOh08BsOC4/nWkETgm
x8Yk2iUpnbKYor5r9ezCFnLTQ1wjIeNMQ6BR8JgoUrfxCzRMUcBYY/h8bf0Ygfm8
Sw6t5uSOXhMh96HtJIJlVfe96vaQjVTJT+wFAn6rQ7ikb4KJCv3E/OpncUccLF+t
tGDI22dQqZMDDmGGRNpOMqq33Ib0GRKIZ7Kzac3D4HVUaSlZeAr9yziJ1+k8Jo2W
0Ytz+d5GzCdO1z8C2xcnKSOBP61XfB85O77kJln59zu+1XEtBv3FP7tSZzS9pKQN
lyvDHJGlUin/wyKqzJGVrDky8mQakjLM/HwgIIx9IRBa1K4sqJRYl80TU5CHfswo
Z1qfptpJz8sLmPcjIsW1lK5aKLy8CMl9wY4qw86WpTxD43dLTkTufBAJlNXrmSUl
jrTfXKckcXoY/pJpyYuhLtU3x+LnDXp+z84rcSAMZ4ZWnI3rZ6PzUuXuNd5KVYXp
tLlc4mFUDrVisdugoCJ7r5ENEXm3ZmnDiBT13JMkag7GUcUJNmGqi7YKm2Gluvvr
6c0lTPjv+PwOr/9QzZfv4/jEGMnBZjMZxe8Geo97aq0K3fRIIyrY+nik03sWIwEC
4S0NEZ2Po+zcNDE8f0mSSQEL+UmfwJJKwwB00oFUkDK20xKSMGExDyrtW0vkPoo2
K1Hz3sDVpgNCl1hdfNsWanv5SCTNEaVBi0S/fQIlaf+mjPtMqFgvtU+64BXavdno
6l0eUwvNtpXdvWHJ+95WBFlzF4Wb8WzZgq6s+hxGH5VZIsgFUIiSieLUgut8TyXm
XimZ0QWAQ2Y3lBfDuFlxXwIgDbQJh/LRn+srCkhtLgXHpPeavI6WKAFRUTtdVXak
J4du4nM2BG4Yzu27utKsoX+WQJznP+h/0M4BDCHhS+Gk1o2cxE4DdMPyWMgYoWSJ
2B9Is7ApjQVFIwo0nFh6neInEP0CPnutnAgT0NDpnQ7FPYCNAwALqqJC3NvRn58W
zZ6lHS87MEoUBK2OC+B0sksBclCVy8EGPLrMbWDXZ/0fjlO42yEhnzAr5hbLIiLJ
gqwEpJuSkJ8SglEDOurX46LCADaUeTD0qXw3Zpp5KggFR+fuIAnD4UBACjw27gCz
z5MSMB3sdk/CvL5wHDV/L91nCF7SBj/La9ayckkvi++7qixNRlrQ5ObdNMubNROr
htOg+V38Y1ayMwdMHDpxSOTCj9iK09htp24MJgnJISDaLncZdIqRIzk1t+lHrUeb
vEupAp7ASUtt57vyFVHjd7pPZDt0CykODTJS0yL1P5IRomBMLDYKRTV0fifV3Rms
C5xMhrgjVlkhbsb2x0FR+oGFZbQpy1cfKs6yueJn/KqXZkFS1esnYwWBQw5NSDqm
b2Xz/c/A8iuQ4O3XspASguLOSpO/EP0XFCc1r9mVewGcciDAkYLvg4BtBtevqxRJ
3meU7wgLz4btfbJeKWTS/fMD5UuslaqpP0P8dzLW4rPA8r7UOKaShT0J5tj85BAM
4t7a6+eYPseqXoJk1AUCknI+d0tm3l+WAv3IU5F4tvhV1i37AJUsneZdKq11XYse
NByO/R4GtfPSlr2QQ+oKN3xEOS65DHKZl0aicG0vPOPC917lou7wo+5tz2kx5bBH
Oln+FrVfuSQLBFEk8gdpavRQoMjL1cFz239O7DDUP9AqjRgGDJ/QQ0spRvr+lATT
DzsQMTMBcxVDzc0PhMVQdVHbEKcc96kQMAPCljRT1jgNCQvf7/NureE8dQcqSuuX
e+4ZMnlhsKZ/C6x/m7r7SYnrKOCdRmqaC2JqDAztinbb+5qGBn4KpEUnpvQbuc5Q
siq3QpWfgIE6x8sga2tJWDLgYlsNIOvDBtxKoZwLfxbAqNPfkOeZbkaEnUmqy/WB
WPEVKN/UrlCezH/BZNJ+dhVWDdi6/+AUoGOMjqwh505dcCKTeO4x4nN3/ovE90U9
zzhgdzsAW3OIl4EhXAX4n0cYrJP2faAMlzGb3wK1ky9UAUiiR1cXK+6tq0LBx6GZ
kI54zWvAoGp4Gd0VP+UbIpteSiH81NirKbc16+Jp1MSNgSqcNqVgsRjhUSfA8vPS
IQKitaqLErlraFyAe3Arj7qBeBm5V4p7RwZ8r6aczfv6fa0gfOwXrop003kOuQNq
Yc53/vpr/yUvDbkfD2ZS6PKRRzRmE+8ENjqr81WVT46xlIRvPib0NX4H5XDI0yhA
DoexY6lME6mK+8/n/8t+4Hg+UQgr9+SfhW9jX1twp/nAluTlNtNX4Ln0TQ2si19A
3OxGNEbywJlx6/eNcUxb1D+FXo1dQTMs1svTaV5DnjXgXhxFqiNgABgwG1EGXeum
L7eLW9n9+3figjLX1LINGBSGxTqgiyfXIlU8D573ylIq7ETsTCXWOmNjf4DkqCI3
sR1Dj58ZzqRk/3M8tjgCo+qQIo65/CJBl+qrrq9RItKgnicuAs8kGJgyOwJ3CCfu
6WDD5NPivHcoLsN3W0E+rpcdUZCzQfOjGUfoNjwhfD+SDIfvwYkfPZWBJyn9m3hB
mEsakakLRhFs0lAGqoHX6I6GU8MfglcxoHznnHhVYcrq2bPUqJq2Z8R05XiBEctn
8DcLwk3Q2JE/C9EwPpOOO4VIrHJoueTSz5Q/YQUGMRbEPnNkPqm51Ioe3/tw/3Lb
0CWDv7YucRykBuxlzrjHK++/WD1czfeVNvTXt2Y4tiOGE10b2rfAncS/WkiI0Bo9
0CA2kCaM7jBv0MAk1vKdyw+AOHaXuUI38o9ck9fseRoG8QBIpuUTkRGyBTI70hoB
g3fbWPhDq3/kqNhJVoeCoMSdvm/1J4xSkCY4oY8VGHA2omLnxP8E/cTiXR3dYutU
O11e3WT7K27u4yj7Zc9VWpz3oLZPHmXLn5wLdxuqYi8dZMkdMR37HsKCddnYxdhV
gw0A3aUhfKmftI0ynF/NpMsjqMHllmJ+BJJamQmBPNsUlk1WJKTLLAENsB75u+uv
5aExlssiwFhiSwq35kd/N6w3cNps5ovYgcvzHyqNWkz3BW91om11BN0S1w92Pn6l
cENIFjnUHxBHsDvb17MK3WiytStflt8zRQBmzkt3nfeMA/hghTVrALvrx/oqDmHx
xhKY9ig9+3lZwjvSENhYWzM1BH08jptiO6lwvYkHkUho6U8vkybXkgqSQ7Q2iqkg
ViVVCuUk93LdYlEl8C+pTO4o4s+jUlkATQ9AHYTItnj/8k5V/DRak2Dg+CstB4Ji
gm+XQwaRz0SWldWwLgmQEzpJbe/BLDOLcZ++a3mO8YYT+JViod3XyLBkNiTBHhTS
UuJg2xdLzGnvgrvpOGZs09Nrc09wv/xtkb0ityDIU4RquS+vCIvYtgbBBet3CkQR
FENf7nJcGyYPiv+6TthQUOaV2iYPwh8AccBhXe1+6eF2OqSf+40hC9SqCUq3Cn71
ABeSR1TajjfQrDme0y20MldqsR5/Scl5EVjBiO3i/ljZVtrwXgja+0mg/dSdESl4
wKoXrEGDxX08evXqzHrpZhxWWJmWQ2BV/gsF+wh4vVDjjJkXnTbnS5xA97Kt6kO4
xECrceMwca7Q5zAyP/HZ+jqpQkmv77HUaSws0NyL8DuajTZZPmcIfAwA9thvcATJ
G3fQrsWZJsld6JGQqtwdIMt5fXc4/1H1E5M2nTeMbm3xRKVmnGp3aQqizML1E5H7
73Mc4gn1X0bSStwC9etlkl8X3nAjYPIWqrJeHnMyCt9nu6Bm85r4iGwrcddHRdGE
uw8fxlgES4VsDyz7vup6j8OpysC+fDfA9tITZs4qJB2OpXe/VnyEGF+ybkW/Zu3Z
L7Y0M+cselrhwpDjAAd2/YkJ4npxnz89PiK0pHCZP5qkb4hRjJ5yJRA8KDDg8L7B
EgmMo3y5MxRdiJT0nQ3EU+OeTJbcRxz7uGgIEv+BC1GZW2DY2IwNFNGLmwUAgyK2
DBg3t8FQa/II8eQRFcNqkeY1yQD/rI+i66/x2CHO1bDBpL3wiXpwluBYMZbjq/l4
A1IDxixTa7sqTqbmZ6taYcwnAmUC8wmKNWNAfmnISAABFr9P524yHQi3yvgxgVw1
k6ADRMAADb2vWclI7q1EuVUYzo6C9l3ZzThSq2LYtPGLpMtr3wGYWaVFB8oiqdRX
2ym0E0g0aQ7qg2/hyEICw/5yNHY2Oli+I5kWicySddjgZsBwfkU0dzBMUm85XrL5
OAgD+UWtbzLym85gHkfeyJjEvwlQzTocJOPn/gXTYMZmHfxs+7pXpb/cI2T4XFXC
7c7u5KdsTnkFc5fX06OaXuZoiLPLvl4HwXKc6TTRUI+/tnr9EQJk6TfC2miCZ40x
4GAWtnX8ZvD3ncg7kdXmh+OPrmk+myLPxOzAq8AymcS+ZnFtnrUvjJzCterfxnMm
n4TymJToeWwr/ZTO5hibEwmp/pbYG4XYjGt23Quxqf2Uv04siTzUaeInMvKelgu+
Gpi5cyi6pfxuXEULrlFaUH6MHIcdT4bJIioGQlVq4dg/vYNzgBwojNuCXAq57N7/
nO7ZoXKogNS948Zqzq3IbsFrK85U2twZwJJKoNNrP2F6NIEMmdQMlzn2G4o7EZ0R
MDXTKjR2X762tLZL2gAkOnUOfMQR2Tk71P6kHaRp6bwAazoLz2NmdiDcn5Wn/LIr
YvZFBzKRUuDXWW8vxohks6t7Y0FvWgMvjCwPXJJywLwEIetOIlnWFLb9ZhK/4Wlq
O7aE/2YcgHzNORK4XSEXqZhKCgLDz+9hYi6qeVLr6Z/hcn4mMPdwobUTc/Ovl0cL
Tnu48UeBF5R1kei7VpD9odKXzMZxoRTqqJftF3rvBij3lasBadJl/d1i05DxJOvC
6cmWPWnVyjmZuRYexBbKMgDjlJopAdB4Bx+vTAj2ZSrye9gwmJN1bPm28GF7kXgO
fVBQzFKTkRietpqbe9zpo/58ETzbnsKmzYUurejsx3ij6+DFxWnpyXI+zvVzmEIt
uj5mhkgeoyJb/2wQ2XA3vwJJbd3OZAup1V79mVo4z8zVTLFa4JBJ/yyIDkMVIOF1
yTydJfH4hh5bbgYC3dGimo3BYOJlqXuZbF11FJvGCVsQGyRAB/6L9UD1yvu/Eker
JVwCQpCWdovyruBpoIuhKaJqZPpCZzj2Q2dCOYvlQPHiL42hv1WQZR433bldn43v
i+XD+F4Ue41fQ/bv281RLrnDTlQCeTFRPw3D39AJz0TVjfQMB8lyeTd3MZ+gsFNY
ySr4tzJ2PoPp3e1EgpVC6OezIJ46YkKdoQEZpLuNdlVpH+mVpOIU1HieNJZ9v5vX
IZAok6lZO51P+G89Sh68xKIY2dlmNB3IRLeIPDCBzCj26309GM1i6blDlp0BLWyY
FOMAlE3EY/KBVI+cD1HHEhTu6t7FzwEwHUVI9WL2Lpsd2zNQizBXXF4n/Mmo+73i
f1iRCM4MASPeQvGv3zgMAkZ10NwmJ8lZNACxLGEo1411jda8Oi3MUU8ywVe2nia5
4aCK61BBF4DguClshwgwqYJLInt0YeLaEl0QWLOOQsuvHmFfufQI7MpzX3C6DrV6
yCk5qLtYe71dMu45wXqW1L9TxwSNMFh0KdNYVFEBmcqgVYlL4fflg7n6fGiVhbGq
e/UV5LuASpd94c2GLufeUCyi9yB6yrKSaQTbq/NfIQVOQGD8iqM0nQF3wVxCiRsX
OodL1cbHivBEbk7zthLZiXyVkvUyUEPS9xVBrIieRXeWCYQqY68rTCZptoyYGhgB
zvVvSr11gWKEzSnKJYfBYqQeszASnt771b/Lty47JF2nZHhEUWIIactKwDZWbmO7
gzTgpoI8d2s/r5pWGfdcNVjqhApBZilgciS7xBsz6j5B4iC9IBfV6Abbgx8l0cW1
DOfrth5cHTpdjnEUvbOjmN1h80G2BjhNv3RUKREvmmzCNabXrgQWv8XNSxLGLjIZ
y0/UmDB2MtA2zXFi6/X1GbYZ5v2ukp/qsQcTAkp9QsL14HDENN4X5mOfnVWCTM+5
vXjcElosD0gj7zqKbiyTXgssInVkDegSUsAv/Mr0KX8fKOVlwco+N+AnusYRyU24
S/6qdYQm5t9X+NB6rpR36xb+rg7bLy46+xOTLuS4fEa/yp4dGa2x5hrMmf+eOg8i
nHRGywO3h9J1VhFmHcv8NoqAUzR5HbSEVDjVyHKD9v/uDg2F8Wd9NusTRfIM1e3c
BfxOVw3rPT0TnwdzOxGOMdtggD9p9aiP4HkUIhgzfMixM7fl6IuVG4G2yzQkMmxp
8WJMXSmunZ4oGhwbXT4owBwY7ZMKKhwQw/WpKvd3LL+2JW3kgbDn/m61XkOmd6B9
hu4eWV6IIJWjsTnOMMNa9ryxWrJqCFxFWSJ1CyFiWSyX5bznI3puOei/KcxpAYaY
/8I9uo64K35EiLh2q3bJ98rs4eKDo8usAXMhUNysEMhmOz+liofi/M2MfGLhuadn
tpsz1m3XB3xStV8XGqQEB2Pjcrtwrm/Cxb46lSHu4eKZSAn8HRWueSM79ROh3mfl
+jgCag+vH5sNzmVU1M15cC+vdkPOuZ1wxPFrc8NearJj2uQAZW/CN0c61A93ItEq
wCfSuktpfDAYwSupoSszv+li3SGOA6XvZ/vuBI3WL8D47vOkW2hoJDi3JpTowWCf
kaZUOIt6k/HqcM77VRVJd8ID5nJh8K+Q8KnywvG3jNWRCVieke2bxtr+Y8AJSg5y
8LWfU3tFrmOzKZbLThj36ZqmMlq+N85mS7/FtoL+s8QPsqMvfBEk+z/kW9yeFMFI
d4/Dk+PLXPBZicJy7wO6HUTpUw5P1j6bC/zA0dR9dwiR3c1wfkYVbrLB0SnLN3tN
rl+zDJAiS3hz9Bc4OE2zCeF1t3u1rqUnA1eaYrI8vwmWpPFh/04cHNMK+tQhPobV
Wm4fMCeVr3pZywHEJz3LPskpcQIELEONHtF/v0IAfsa03/9J+Gy/TNwl4O/ykv1w
Cepq7C+pL1N0KIUI2CdDB2NdMKq3Cyqgx/n4rG/+yy/5Fmz6iqlTAPT6G8OWGhVo
mbznN54Hc32Wsy//UmyKWuJw5SA+dOK84NmpGzSv1Duvp1Kg4E/isRL1puFG2LG5
oja9M8arY/OmV46p7TdwAhw5sytjJSOCu7MesmhVNHnE672X1USCtFouE3u12Wml
R+ltlL3gddjCnIraEemLRz786iXX8GiVQgc56o4EY4jtW+9OwRNFEP8DcSPISaCp
7eUcxVnES/uWacHGXdW58Czc6cCw1li2GMoe03y/LmRHAXV9VkUWtMJD0VoMnhfq
e50iv4yqSmF0yzjQlOKG/yfZOB8Iijckc8EWVCVUjowFMQ30pqwR9Ze0Veq/juFH
4YWO4Tp4sh0vtjkjqTOipNrKjqvfY0pDzFFNBQg9s/Tp/O02MVJ46S8eP0s3sy3j
PfvAezSgMdNWIGPP9uPt80ONXthjxWb0VXWKy/MgOtVcC5ZicSbKisCSUR63DWye
F4Z1MQjy2juIfu3CGXRZJETlrbuOqRfRiAW2Lvqdfp9OPd4xuFaOrEesQjOYmcI9
+PQlk5EYGahslIwzkC+QCz3j9BQOClqoyxDTTIeLMR21ZuJLtkJ6g0pclg8KAka8
hmsscM9dXKETx1t6YN5nOpZ12Cywqad8vopM0M3uOAKM0KL9rnv0spzBkXzQEAid
LsxtbTROBXQJSMQN+M+WZlL6kJllUWqD+341CXmliZ1uuX6scS2Pmv6YGjc8qUV5
tUusOp9AK7IT+cGuYinSwBFiMBMIQpqpF+nNfR4UQbnZ7kNvdGTNZ/gM9QTIgCjc
wyNTaflWPt7ScRKf62GcH+djsQrw+mNAKOXE1ss8/zfy4fl9YAJkIiahKnl7Z/1I
54Z3l159o/5SchVry/SrFhmbdVHJnku5vyAfw/o7OSIRTWItNpeeHJC4KeatHGeC
fodcOg97jK0l9W3fSmx+OT9F4N+HsQWCZMlfIfYq6ZVrzK/Uvvsqc6mSS76/KjAr
nVBLDn7FzRDmFHpp+AfgCfvpA5Mn3bsKrTF6I5TMltKwqqzVc2PeUzEXWTQg3c+z
XOp/kZuBw7hpQwhBImcAZERaQuXlAGY9Mt9IEdiT8XF3hodLaCULkI9RnOgZk+o3
xWnsiYUqmzjWngJrN+lrDPvnxj/CXGI9ZTy8K7G8gPHLATxrj5sjxZp8Drqy2DpM
hk32P1YlkVJJgbL+3GphWXie0Ua4O9IcpMOWrKKW9d/FHZe5Gvi0FY5svo+N7jlg
D0GrQ67Wl7t9N/WgjsGQclpljHhiA1ENM+qZhHAVo1tdkrJpTce3jSJ+6DIMuxUe
LwLxoNfTiQn+pYNb3XtnWlk4rcnNAGx9Qe3wVAr6Y6belXMFqSVrI7tUieAdYnP+
9zOzkB9U9ZWkCpN++eykxMjSdqPQKAELHVOmbrPZr5hTMUCAWWy4kC6/ubXCz4nh
wnX1/NDMrdBJC/vAdTH2xrNDFbC8+3HXKowNreNWM8GPnyRQ6YSsGKKjCoYOb1H8
3e5zvn0p+d32fMPDDJ3yuCFbpGevb++90BBwQYr673hbvaNlWqUEfG7uaLqGOcHy
99N6YU5xMeyP7oeLmLM6CyPGwhL6QSy0EnTxO/BGTXQ3rA4VRCVeOsE0xeYkCwDx
Mfo2i3L1/ohZFKuG3ylwm2jvZqJV2PfCnpdvjuI+5UpM8B2CSyLROwSYYplx4krL
KWmM1pc8I+ILny7KV/tF0EGRX2zYGIDoGE0FliZbjGgS4K93FJjVD8XfPl58cTB0
dX2ctOiFNCBAb/l09T/RUivY9WboIBkLT4SfnFTgIt/S1bKLXc2FNXpZ5W69Epjh
l1vPaq5yii9ftaZltFRujotK56oXAVveXOf5ab+8+BMapK9atVw9z8zcO2DN3gsZ
sRhv3ec1Y8dkPkdU8lD/6GF97HrupwEfL4yAoO16QNkjECjCUw8EzzGoPvFIb6bu
CfDgDKNg1XDxx2Rr7hoEpXfX7zaJIzxsy31zv+dw38mu2Bu75PlKuzIJy9L+saSU
+BWAT5zXbZcVTBN/UClswRlpkViANNdifDt0oTYeFQH6/16quEdPwuOCrr6SVeFi
7MjTtTqz21lMrs/Tlm5lTEiMDKkg4OwOzSXA1bN7pzt54ivwIdgXLA6ty/v5PYCl
jDrKouJ5/OhGxauGR/QbMIJcCxuoCqE/IXNU+Apm8W2quFJ9OsAHhSQl7zPoOzLf
rXvagxwrBdOOKLIZrHk80hHM20Zr4KcOUYsnaNykIx4tla3fN9+uwe6rBX65Arwb
AsWO2iDvQRz+7pt1TX6ukLxJhXrYy8X6r5zTo1s2YkYt8sPyFlhYgUPacePHAxq5
W3zMRDHi8RR7h/C0iXoFzOU9wZt9yts25IfyFkYLNgGdbsUFQ0EXDQLuaFhKOlc6
/twBTFOozLh/yzICvDEfqXNjZyj69sZkCiMR5LEzqXwU4KcNLx5fwoBuDEfGDJc6
Jhw/dNFZbnYcapdc0tothtVtfh/De1qmAk2Xe13QowQXMxK11vwq1cA8wzudZ+GF
VPnB8+Yk1L44muUFFsX+2VvTzIPDUjc0c155fokEOEhFfFjhbcR1jGRyQ3+F0nwp
bVRPJ1GSkXOtAxCZUhpUyfNeJNScGtLMQ1z8gsaJt9dvZ2jGoOPxjvvTGR8Ry6Mc
F9kTtksmeIOJykR36lp/1xEwba/2fDI0MwAE3icNe5S9QWNYhnpIuQmwc2R4ZCmA
cS325CD3R+deKIg3hulFNJ9lWMBLGIimwcPVGPMpT2DM/RPxmjNYd3VnyTjJbJK4
68s5biPYumV408D2md6/IH0quTbLbcL2cPQh+hgIQZ2k1RXWkggLH+LqIOS/L9wX
u42/vzcYBPiH8sjFKMD2OlrZ/u8hBnBXOAANC7BxRvc6YNi2CBwwdF/sR3vcVzNY
d8X+g49ypT5XBj8XzS75Mg8wahAnk873TeZU3yf0rIq9LW3KCcuB8hoI4oWyanaH
NjGi/MhFpgOiE0v60PWm/Y8niS6rlCskdopzm0qtD96kdE7vQozb6QK9vX6r6OP0
+GXh7CYP2tgtx9W8AEChR243cBu2uGKo3btxGctSAdxkwHPEzsV54IRpVtZUGXGx
KB53y3rdGEIyQkE/qq5Yup6N4Fi64pcej6b6xjbJPq47LxVskdsZImEKQiPJUzSm
SYuzVVpy0L8iucL6MTOgm1v/plcD3SM5UqEt/gGS8nME3G60+m/1C30Na9jM2NOs
GxPQcV1lfY8j1IUlxGL+f8bvO7sby0x5DhfdfizAChJfHDSoR4UU0ORQ/onphqRi
C0YtsOPiQ1ecMUF53Imjp+xRSNXSVgF4H3lxVWVzdxg1tyKtPoa+nYUN7+24WhVF
GJ+/c/evHKGtH2p8kZzfDnFw2ybJsAqJ9Fsq0xXIw+hEiHVUJbucUhWW2GxvOOqA
8Oyt7cj1dLz/vyvF6H7XPI57v7d0bJBV7DtIaL3YEjhL9fTJ/Nfl2XAF5aOol71J
56zT2/3bjtoXYtiZhhGNT3Y9XJbLaPand62vkmdL/Q05NuIWk1jtWlFzt0ozWkbM
YEa6O8LpXl+qvWM4taYy8UdWGfuVNnsxOI9SoKrad9BCioCrKRNu2ouLLYQGzv03
ttpjWPCtLCane1VKIcFN6ExwXqOdjA5Iq1PR+iU+QGPVDeMceTAdBrAzSEnp9J9n
nCcVjZzqsescL9q2U6aGNHLoK6wvnVC/L8CYECWim4Ziw7lPmNDkWOc7RP7BgntC
lT5T1bDV/Udtg7VQHL/+ZpkZd2r6Ju80ONCpc+UiPCIeXtBXM9QcLBoPKv0qeuBx
qvzIAKk4x1OhWptvUhrZ1ugcN8lW5Z/StmpPGbu+vABEAB4dCIok2ExgrWuGGjvB
7B5uw23HjWkaPGUcYgMwisrr1Z1fJlGMOAF1CFbqSu6cxqQ3HTz8mVbNcNzrjp7C
eJyNYH02w9mgkIPoUzkC9wdWp+jOb0Fjn+Z7xSGQzC0MM8OTJTsNJ8csWgPLBNDe
WxIZ20Kl/oW3yWlYsKdrUU58mmoZspAKuoNfcH/zKqD8ou6mn0IaVApZhfAVQWza
cjwdHXw2tMnKYwkS18z5t66l6+w/fHK3j9WVOpJA3z2wpqjYLhTi/wakNGRc78Jd
7u/1KCXm5wYEdbIFqbtAiHMnRZp2R9bfYvlVxua2KqBXLn+4SjWkcRgckZN+pcxp
2KmZYuVsvAFBd8M6B1d5cLK2h0LUTYG1sMAjAXV3mygTEnNXIjRJpual2Mb9aDHG
NN9N2/s8sMrwPuhElkSqfzxntt5TR2SmYLnFWsf4YmP0TwocfYip7fYlkmrBNoLi
kd8zbD6GLX4SzUoJfYcyp/JJ3kZAz/O+fLFZK0VCMb0+eFRTotaX7MaA0k3+V/UD
/x/v+Rn3s8dhG2I4W1KM8DdNP31RHftvsTVUIRV5rnU+cYQjfoJF47zhv7wY/XKm
G1jdfWPZh5aLmkSJEa2zpKNdRSiQ41/01O97hGKCAivh08rBIT0ru3PRRq0Cms33
QkDWor/Hf70TTqvHxBhfdL7o0PU6DPcE9Y5Mj/PfuXivU+7VX07Samo2yZgDZB6W
Vo+VjIUB/Q0+WYzRrr0fnjUD8x3DdTE4HTXo5oo+VPAuGjYr54uwfJTzfD2Y+Qpq
WwvbVdcs0xw9cUQPhHM2Q22thn09d1tMSzvouY2SLR9QMMXa6mfUzwnhwBrVNV7B
rrKxRU6jKfyiDulqOtnqK386di2CEn3z82nSW5NPpDRO+a3m1hN75i9ir2xy7BcR
Yj5e86xIgTy/QF6aoQaqNK8c1vnN79D/xRrjHvV47gczO8tA7T8BEqGynLJpiQRX
UggnCp3iGexgbWDASX0CO3kyr/8wIe0bmrR10jWW2ju75m47U7/vamjgqkUt0jAE
T9heirapyoANg6ZrPD40oz3RIe4s7DpUlNJyyTgpFRXO1fL3OyqST7vOqRwhIIwf
KNa26MH/xFCo7ykY0HEC5YKQazsOu4uDfxGyTUiZoFqER8s5NkA4k7p3j2P3xr+/
E2wPGcWd8poWa8qXZj4JOTyFtbiIRFNRaxokWCWDf9WLV/tJQHNENvMYoZUNntrE
V/pCQss4ykpS2wJ9YldNYuQWezAx/anHHOBAjQ9elJ+lb9sDU4v0FCWyfOIjuYw7
PMJq9HEff9AwhiCB3vTc8djT/AXJ5COCiXg6Kmjl9QFcv2GTI4YpkRAfi5Z5nQ30
Whbzi4BEX1W1gCz0q+DLL6e6QchdFCnyoMNJ/x7VGbCsJijqMmWjthuW4Z0D5A4R
Seswxd3bZpu6gt/OZr1TiLuFt2VQvv2WSj0wcK/iDNuy2Zlv/iX4xseipM3kwxOr
np4YX55IDGNfVp3zxFvXxcYwnb3bl2shuS3NzCWXMMPopxlZcPbgBBdBPtDh7Dw3
0ZtZwHVdGVO6x634M7hRUVRCC5xTWOFd1LWGo8tjbKPCK5OKK+V43ATSHJDIqTbU
/kLcwpLd2b40Mtx67XjUAvI3sEcFjvf8Xz6mXoiY9C0P+roZy6vjkhuUI0U64i0P
JFJ1dU9ogiQ1U4Y+wX7qJmN/Kkq7J4w6Su3ODnZxQLoexXWWPIWLB+IDh3/iaasj
YmkK8wxsCwjb+RUKgbjpSuDJFj2Lx6MuujzC0YqhlMpaZGiXkOdKE3b4e1544j4W
NodbVaqclZE8tBLKAtQRlR9eK4EOjiYBRzGF9YT0ktPDRbFUDucpa33vwBKKrtbM
f4iVfn49vu2y7jpj3InHOrYcad4QMJWhV6NUc2stYI00bULOe/oSPcv4tlSGSOiX
hj2RkeqfI6jAsW/0hlSJTc5SHBp08upDfPgqggXFAt1Q5x5AzxJWlOBD+ueJ8ff8
mWJv/D5nRRYgnPWJ8aLIYMX8JIA3DqHmrLWsXKca8TmCyfpGI0WVvjh1/JC+BDJn
lNfsHdkI++9ClQHihVLGL4O6qnuujY8gvTicjDzwgOdRBPBimk6w/TZi8xREh1iv
B6nKvIo+cbGpJJDmvArVbglQlpKZEM3r2qdidkMZtpEto6XkymiRdCG9ym1c/y3x
mdT63yag+uoV+hk5Ru/h5eN12TJDpkzIms2k2w7q3AetkZX6MJreLis2XpA9Ubje
XHYEQBU0Dori1hbNjkwalEO7s5UXINtTzHrpFbfTj/1Smiua6PYen8MTV8yWwIrR
yG/PvJFYCndfnudhDpFaqjRlQd5U8xUE2UMY8+vCNtwtOdkUtkQvYcxGl+hWXAJw
I23QMC8mFY+UQVlOg83YqZEwEqU26B+Mq8EL8KeHtC/fQQXgCiaEnr6Ni8tZcgib
mhVF0N1/z0IiTWcp5ZKKSjVNrCBxlE8up/S9/0q+MJ/P/a724JkWV3AINWsFiMbB
IzeFsuHQMyy5qz0IbYDn1tyjjAxyMfZlDWI3mp7JGr1Pav8IZq+/kwurp8i1MQkv
rN2MwOREYSaI7DTfTOak3/BBU2V2iimKa08HCdKMo6T+SAMh6nqO3gV/0p5pklU6
M7XzqB8Zm4INIlgeKLHREFAqxxKjOrZ8dKytS2NqAaar93MiU0YplBkuxIBJkv9W
RgdT97OAdcozTRZzynRkjMuBHdhIjwdhhgSJxFXk/uhcOOP3GoKgI6O5UrPj7WHd
I1HCURUBQwOnLiC7QEQdqImO3QcS3qiT/zZ7dqal4F2N9dm69cVJvpcBYf3BV9Yt
UGIhrJWyplJ9x8ZbuJC/VYjIGXaX4o7VV+KScyQjwVtEu/a5tJyrJCFbl1VkMMoO
G7jSVV1gi1zEmOkgMfu3oZ0a3BET5UDDCpZ2mHUhobZzDdClFPwplHSYqtWIi6PA
zfxQvj//zfdChSLr0rQ7LruKUZfHdUMDZrnCJ6zVDycLm5Ciyk0Lown7k0585uA2
x7BzkiMzbY5tmBC6oBtZHlVcj9FUHFkiWnoDLSHtBxGO33b+ntSsMIor5AwS9AZd
pQXCEgFkb2ru1CVkQnqx9lSq1wBIMx4fb4Gqxb+xUd2B1N8UOAA9TjSEgRDnaZ30
KOTV5vt2A47TZp/VTtC2X/nY8UY/p98rj53d/EOSmPruP0yETu1GE6/+xxSSanjI
I2XL320XkiVwqhag8OZKHzr7Hsj2vdHJvGNkvHMdbaGq9yOtFUnzypEtGM7KzLKu
wmgo3TI95w/AbA/rFEAf3lfBIPTn8F4IIZI1CCndwnqOKVrS5zI6wnPpIcug6c70
GHoIyeGAGK90Pn2gRFJeo35CN/omINgtYm5P8ye86J65/mJ4SfMTZ1F8oD+jyodr
Fh9wnYO/0mM9WOg6ZqD8jQz/y5lvZQXfserydiHMM6tp5NEavjlxG0RdmMn+H4wh
WmMKxMsbsIm4kwbnYf/pLmOgPUEVoxbAVEMWZDX2brf/IphWBIED3Rhs6W8oM8GF
IpKUeHRwMxHZN89ySUhHlw1mpXd4zxEeRtbo0E3AKu5Mx7itoIKeI+vpjuBRw/Fd
vuhWqmIMzEKCxVvt6AKv226HvqmNRAmL7KtclncsJQJVaLraxUhSuUhbPPSo2M9B
fQ3KwSRu3hEXJRaDoj3UTtdrLJxZScTywPlNGTjyz8tAp1p1a4GgMku+GybUc/CJ
s2nG6xv+4xfdQLW9JtaUoYZxWHYFZ5FXn/BTXCWqohvhuyk1BfZVUwRtYrFMoSnZ
MhMckmWy9oW2hB6tXH9nU+FHIRnpBO+/ZA4A15F/vPcs+roWt2orKQOb7Cm4lEx4
SfnrH5rle6CpgHnFZGPqyFOl/a4u6nk5mgDFKlN1pjMEmqOQi9qam+lNwdhqzx8W
TTqFtD6W2Yhrs3O3hLsGPFQYOxeVmwag14s3BRvVwurOH6lo7ygM+BewiruPiUGO
CQPg2Gn4Se3vQw1W8QxJ3ZclkzTYQ368db0Ug6hzQRWgK116WAVxYQ6f0EKX6Cu5
n+QZlW1A8O6NOCcPZqOfu1Z/3snLycupeyskYdroVTiporzU+dEMlkKhb/fWAeYJ
ovB0XUSz3+lwV3vRz/0XhYs4FW03k09q7qEyKg2sujmVxAPjgnK8yKBsdGRGZ3p6
o4bR/n+JC9wuh7V9l2KwXAAyyeKp9xjXNRXnuaPji5Z4Jew7OtRg9E5Ct33UBUxp
4EbbS/rTecXGMFetPpxWve+hFTVWxPgNIOknLiUZ8oREgNbcdxVrRAa6541DC+mK
bC721Jn6usBHZaQ+9ZhtQdnYLje4UZtl1bDNV5RofVCuIxYxWb2E7+REhrZUNWQm
cCq6RJD7pcnbwzI5tdmUwkky9mzks2Rlgv7+GK88PWiWPza/rWq6jbN+6P5FOodm
XEX/ze1xoqTjZd/a5a4t5MfmaV7HjxtdaiaoFU4oooAdurtGrP1EwE6gQqpQe3SQ
FHS4rb2xTHjR3W+MrCJj0G8whIBOqZqFS54n3F3/UIFPmegu8DLcYYvhFRomg/t6
fVj9xzSIJEPdVaLCxZwsCtllsG2NMIfUQ9CWSOLYmFJ6LA2QnvEQiRDyUKIO/wCk
kX3x6Ii4Oq9H1+nOXxs06qWyfjum9N1QOT89L9wA9IliPu5AqB9qwCTT88L7ynCA
OexVtBtYOfr5Q9SKpaKyh1b6KGDT/bpVdLKc3P2lZaoRc6QX+KqvK1GCJ/Ey6jia
fomOX+/nJCZ5K4J2qVNM3Mg8OwBc5h8EOMDBmmDS67N1qC+42cbtzer+ttE2MI/G
QF2EfLvK531xJ2k+twxCwcwP3uDddFv5dJ7eZ51Sy20XxgaRO+3FTxATjXKBX4hr
AQhTr8QzcpuTBG1xOAdT2zd69w7fTe/TzY3I9Delu4SQ+hO+QAKtV2O/TcZ8v0Du
p8ZJmWZ86Z5Im5wxUKXQOuKK/7PGC6zh6qqGUQG9xDbHsGqhckiDHzsXRT4y16l9
/ASBWvR/XBliBWcnVGABkFoai12H2XPgBpNKCOIytGidzaWpb4K22r2Z1iaxhStY
2kZjIc+2erlbvPCvL1+y3GVj9mGDQTdtennwj9QshIbBX1bt3m8xvdY3Hhd3xRVa
hwGx+aoHcMhPNkFz9Z5frset/I31Iimzlr/fkCrzoxqlZNAL1F4a8FOYC7fosJBf
3chT6OIvIsZ4BalUyuKbXeC6XTBGO7Be+/AO86r0HTd6SAi0m0WTaBAHUAoDheUp
/0neqnxPrAi/aWdWGt8OoJ2DBPo/sRITcaWve9HvB/pYTPx0ctPfO7RLfimDlYIg
46729m/PSfqOX29YH/bXHm4sVqQQf7igLywtmUKNY+5Edr/idnCuF52cgi0jXXZY
5kNUyON1Qx3+1Ven0rKSjC323gSon0TEMBzQudPNOpMCUMoBjC9nNh3zrpls3LzB
74cZlVIPdW30RBnZszFM1b5FGu4gVQpvLs8yyM2uro6OugD9Qc75VbiagQF9Ij6z
YvTEwywELhMWVQ8CFLlIL6WCirAjWpp5JiisBfpE5zp0bazhI6XsWtWQaCa15Svc
cf7sMXz0sqmEI1mjmbWV+YDgVYrYQK++4E+zZkU5T40rvuWGKpayTuRIhYqi3XUG
aAMgNqz8lnVSPWc03uiedzlNBh/uolFlkbeJDI4PEFhi7CE8dfrRGnJkCCwrddgY
PWhjAxU9SOz69XrUuz6eiCyoaA88sI0QsG/MgkfCfql68BNW4mBgti6rekcuBBrA
5xriuYMciS+PTEQddrcV1ThJ9QYvqHCbL2XTUBE1fzHuJUooEAVAoxVY7pIDsudX
GnDfsECVDr9LJ8AfjGVymTVk2mKPB8zuZ7HTJ0swfVj7WARiDS+UZLc9cZo4LQg/
a/3z0A7Jsnh4SxDdIxkZWGrPw4gGyoh6mosMwiOSPk2rvPtmHkWbAgESf4Y9RQ0J
4LedIFGu5tqDcsYeFZugOcvf4minm7t5xwNsrNu6otQ26FPDaxmw8WJcdwSA/wo6
2FvDYelxcdOD33GCuZleSiRkPk5+gHJylKjnfgQJMP0YIgX9BKhFcQXhkZvJRNLa
04hGb6nV+mYmbzAAWJSMDdxjhphCc/cmbkuxiGY037gI58Siw1XrtUPYS5h+hDZz
2Ry6KM0M8AkjFJmxqJQPfhDC6+h0NwHwo+OX8eF7JwAkgkN4ylY9PO/mjqRsAEJR
58quyRd/4ctdvGbpxOxC71hJtmuxW25rGW43Fgu9fexBns1QiJPQt9DsK4Lmk/W4
dgl/ejC7eLYDnJNX0d0ozkVsaimM3ybu/rR4jRFpGj2EWJGsloepl0fh3p6Jia8K
EMvBx4pBp0MofJ010CVzxn4d8lv1b3GYiFPkZFW6K2RApsMberrsrMSmp2NgX/m5
L10I/OL6+sxH+i1BxSQVuumHaku8Rji5zksys2iyM7lZS2FpeFp4ZrgNSrZ6lCO+
nwcSOKQ6KUCXrr3WG732ppk3tAzGq13jua6En9E8A2quJ/Mdl6VKbkR8Dn2fCGCF
pf2dITHzvXAs/VJqSUNDI4JD4yaiujHTtFa760xBwt1obiwANDba0Rkpy/4LPwEX
lEH8Om1Ww/auxslAZ7PAhRuETivEJQfTPmre7V/xjGpZnKGpmGFGWbXZi95gOjRz
OqbxCrhQVh6TGSInwsLiJZ3ktYVcw3enEtQn6pkfflXP3JMvv6/i20/N9Sw297Kq
RaYjYkVeTLr+wempk8C13AuwpZjHu6WquNrOGTV3aVkvGsBgtQRp2EytPH6jEc94
DTvo0bi0bb808Xz25lOYH4NQqLxMYCdJoR+FrvtogE2qumSYY2s5Ux7ngJzt81oI
DCeDiLJVD+DDP8SoUqQSUIsH9e8j9iHkkJxuEhC6LslUapkNaheHNpiqZlS91IJS
VeX6+R0zwoLosfnTbMiQtZeVaxqfE1Ye/pecr8k6CFvXp5inwSUEetZbr+3LCk3+
jcCIOM7AvwTvCJWsE12Z2ADaUtJ2kwGAXf4Xuv8qIDiHc+FG27xfXWr34DLLnAE9
w54wAma/o6hZ+8R03+fiKQrjX1wQwFg/oK69gTS3Sflb19iIKhPfse8EBeL1o91N
FQ0JAaSmKedskJlUgQZGTJWM0FKx/wcE35jt2GpQ6naCq1gwIZjGqnwe85tYADzJ
uN0PCWn86GEc+bwkjtfZ9TzY/hzruYTb1FModJ280WRWnvRiyMVO+puNczvd4/Hj
4CiqMgm8gfS322KTwtRjOYAZY0yN+qlQ2Axe2FRyJQ2GByb7baqPu7SoeabaSnpA
Vf87pDM67XhKLBg1O/9RqWfsvLG2pHV46f1fZV/72F1PX78uJgkRL9GZ7P7bw0j4
/buZJVRQKo0B7PSjSl4nQ1Xpm6pX5ms4pHLDOzwiZT+AebQZtu/IUyQwid85Wvky
LydQbW2HbN0u/IM0FUR/DkAbArIZ4OgucWojtC6hqpo7e6hoC3xmBZhCfbvF2bRu
ONu970xT7ljKGQNIqhEc6rv5t+BaOHKXRjelpXqUUNf4K+JBfsZLeKLoz1v6Z48Z
ikdPFQ+lSypNMB2xcp+QX2m30ABGQ83Lm68+2vTEx0Kux3erTAoz+j29fX8x7Bry
r7ZPo0KfnioWr+5+g3vzN5dJLIjzS9HaaOOBTWI+MgF9JKhOu5A7j0Cy+nTaRIQI
AIr99u392I3arwfT2USF5mM9s973dqXgJUIyadnxB1h7XRzPjSIyBQ3UFCcAKMoH
DSTrCMtlTHmCY1r0IpfEpN+ZOz0QS1sIGjSh1Q2dCvtLa6NrYYj6q8QVU6pOkm/r
NjmQWTuSgRkcH9LgaUa0LmwxlQcUzHuKWEO4iVkEKolMaYz3Hg6aW63hHLz+TveP
uyi0qtDX+/qE1pGHYcUzrB0IzXO54bAaQSV2NQQOP+ovrDGMdHP179i/a2uxsaPy
fWx1UbB7Yc+KPfZWf/eJbPum1A2oqrSmO3sOvHuHeiHAECKUISbVxWmyDnrqlnRC
L/FsLqOVxXRI4t80EKl+1Sj6Jec3G/6YVHFgeFzkY1yve3ShgZGeNJrgyo0/vRt5
AyKLHs4BRlg0JEAfLZTttNUWeI74FKX3DIfs+Yq8QKDi+f27T4y/YBz/goADgMaJ
FgI479Qt1zXn3DAMC42ILLd7h9KIMCobuSckYgeOt4rQs5tQjaIRfC5lFzq8riSm
wbD+LCyK9K1rEdob/0cKZAsG8PPnUincBCp5IhYF9MOIVl1WDHp/AIDHL+CmDmdz
hdzqB/4PGoPLmUttfaED24WzRDQNZw4okM0LCQ1jBuZcy6Q2LX96l1yYS79bkJfa
SIE8ynlqAmu2hijCOSq4OnXGkuzJsb9boa5yEZEF6Dtx0N3eCFsEbhR3TJohbwIJ
gB/5BIzB4UOVUQ7tD+exBFlcv1eJx6jF7VrDveMY1wZ2d6eMvC9C1QQ9ZkD/nav6
l47SpiuaPdfGKjeOFol1bpud76kYT6Z/2Ug0NXOCK2QdmLrWh6uPjJYGiopgoUYZ
+PavtvGvNJhUQb5ZUcqIZZ95GKxLpfpsiEYd0VAguxQq7EFWcmByXx3/oPaAmAB/
g4PQSxhFR8RMptLZrOm2v/pIWozm5JiTc088N3x2xPPrAsN+YmIcHtZraTyqPAI1
oeCSAoMuwos6g9Sn4AR+OsBlEeZOYCBT120nLUvQcOgBhrIxP+Uf8TaSSoP1zee3
7pDmsKT/8htw/Kc6LVSXFiMUdCo9niVDyqnTYMOZAC3CSasrr9TBHhGBZ7+52096
aRF8WBrpfZUb5/HVHI6X3cKTYYh82o1gY8oaxQireKhlaArzufKzz2BGJxDRrtV2
17mEC3XrxlXHUsCzUXd+Mr/tkddkMVUqj1nkkC8tsK1XcOpcWq8yDtqOeXG8QyhI
/K65/3OWLJsKLomgpzzHNTFNKOGYjbVXGRXh/8BhBWQGYKl4jSVzTiUhyWFXHwu6
FI3KBCpxo5ZZ+nDPi7AuN3DUBKBaV1aVy2lb+DyPw/JZjI+QHmDXtKEZkaR2Poj7
B7aN9ixr5/KcI9bEw2J7rCgOIqEf+2s1zFved8JHcwHdvBHojNcZ6fCPsUMdPRwp
DxkpFyRlJz68eX2dpjJ5lzRbzx/eS3Zj21lrIQWA5ij/KYL/W4/dFwo+OUUHI0fN
OKkS+GyE6jyXyp8rvtAwlH4mPY7ir3nncEC+GoVpwTiTh/oQdK8wHmFsc/w3mY5z
tIoJzegut84myc1mF7f5XZJxDi3sGQOg29HGVNGR+jM8W3kx6A4O5fPrc0oKy26p
+t4eAy4U53NSVew4NRYz6J024JWfFY/OWBbPLA2vMmfw0Pjguod7W4u4d+lO3IPb
e9Rd0QuCcb2jyJEfZwNCK6dNIOYTDnPkW9DJN4s0vbT4u+F6WqQHdoP2XmN4N5tW
KrZLRmGDTPB4OamaHxWzIEDYfVTlp/835N1iR3Ep9utg64olcX1YN9Qc3QcYsk/o
2Veerw96NCqN5DDEKsZ5G7ip9rHHR/cgkUvGsXHcN7wTcPhg+TGkNJKNDFNdAnaa
D/f72+4Uh5kHJqTEuQT+PkjA2an0iLMYQNObokBZdgReJHrKKRr4n9jVm587Bf4a
mwFjRVBxTVnnKX13psShFeFV9vJBnGsnFDBVdTAihWzkKY4j6YCiZT91AiBA9pd5
VNt+AaetOW+OamTIPrJ6JfUp+T8RLJcXlGG5sUfXvfSlwOrNkZkpFHraWlwDSczJ
18brBzR8pswwY8GL3epQKnox0SRnaFfSk9rvMJk+89axG43J6OXHwT2I/KISJ9Vt
g4XsPx1ScBnEwbRPG/buzHI86Z+YixFV/fM+9EW5/1KAkQMHt3n0ca87TJYd0DXE
hsn7p7iUm+UIkcAG5RAnQq532zOmpICa0RESy0JKOi2IWUtdJFNIYPU4JvD2ad2c
yF2L53Wf3o3XWtsiL/m1iv0RMmLk5WpKegmgVG/b+3hQKjx+y2WI7SCidn6r9Qf4
TmMl1nN6BJpNUQqGfBe/kc2cEyR/2rG6lMyHbtSp/Rv+ynLwQ4i016nGRvhW67qI
eZx3Q62+ulaZX4i5B42/hQYYGICrOwU00kdjS20b2BixDIYwQC1ydp9nSdS98Z+u
02HzQ4R4fwrx0kC378Id2/7yT9qUfahYJOqBOC6UDSZq1UAh9MUVnDl327kPzkj6
7dMDS0zy09kYC1UFgWrhTCJCdwHhtr1Rd5fCXz0mVMZNZyJyn2WWtWc8o5XgQP31
7tNnwyUyGi4BRlc97FLJDGJBBjzQRqAssroeilwCA7ToD51U4/JZ8kQBEAt2FJaf
ZgcWBn6sjGzWU+zf4sqYM+nv5Z7iGsRneYbyI++P2fkDmmeNu2MF2Ew4/4qp40q4
FVh/8VwZAkctw0Qvt4+LSyiOi1oVDUaoC4Jp3TWc+gM9fHRJclA7TG8cH/FR4VYn
wlH0bD8mjHbHqNcky721YwEaKDLxN1wt+CVxRR7fvXzRlE8EQqH96M/3hL90/ItT
7ZjTkepzS0VoFJOBXdTTeFBmLP4cmKWSrvY5zjbQGg+NHtkJRicxOFmnV8aZJnge
zU0gTVsjTST6uWNm/TBovi7LVuTBs3A4QfJPUd9F+EoNF0fTWOIy3km7lVbwCoPO
a8gkQkkpKaaxy/Q5KRH9X3RMe1TyePGV+1tVa69v6L2ttNN2atD7aT20DHvYZm7O
G3biv+DINf4EoxU7PgSFb9+fbIdWioLcS6D/ueyLRUSi0HwhUcM2nGsxv/MsD0DX
FLTSHVt8q/wKSqz72md1qrmb8fXk9cUtEa6/4jvk/xRYzLkD0TB+RGssIVXSzomV
Q34msDJXcp/XEyzxocdRSoa81M5s+RGLTdrHV1YwrdbGNCqsOrMHtQm01VwBPR1U
fmJGn6kqASidz0LnRTAghRnTusGU1q31GWOJQO53quuLY45CkMU0u0TyiRyFBzNn
pMY3f46YIn7ItIPOF+gyhQaHiIPO5HuTs9sPHPkRszJB93eQFS7e4VwzmGeCEcIp
P1cjvwVQfoiihWn7olclTcMxE7b65JbBcdvxNXZQfRBaKQbKWAreyYZl0uMHEARC
sYWIl/fv3EkUDPxc0qO5Ou+6tWzcJbXA+sL9kZansIWZTv/lh8Ota/E8oGPSF4Iz
M3sQfwE5JOfdt4DCeGHRqPCiyEu9gJXnce04tb9bIaygWz3J2eglS29a7ZcTjzqN
d//5Mh9jTEgpf6eKjokH0bScFP0GVp9mT5tPbu6OSSbrecESkeN/QKPuZt1jbPvT
6RAlPCB5UqJk0Q2j0E0GV6/upvWBCU9T0OYQWXacZVbygP5/N0QO0ONYnVYbkfuI
WXiZyPeF99QrXnFoSmn8oAnub+qV6GNdZcUF61ibaOKzaQFx6JjzJPelbMGhrgxf
Eb7ydJlQOUmXD+s4ho2HRtLmzBeCrW+56aznRzzlEWCbsrdB73bcYNIzsNhVr7Up
dsKEXBZqf5eJlhW+IPom4jDl0lDShShBlWXnQn2RTwjXxDHJdbIRK/qEtm9QjHQP
5zS2CBDijtvFfaKe33u+HISfXnXEfpGR3a2haBhxxceH/QZQXO+u+udtzL1Ve3SX
YZzw9fqchlYqqbTEebtTFu4GDPzorQr2UuN6z/Mhrr5OLrXiweNjtpJB7NBFwF4A
oOwcd67h0DI7BfhrKajdEJuH14pyF8pFtIWp0HCe06SO28NAq/S3j3BK4qhsxRoh
KxWcukZRjBDaNf2BiLf175YmzTZcga5Zib1Ex18Vd9rWNFdYUpAO+xzccjbjKrBv
9IygOCLoORYdtLtClPtZ5AYdiZaUbJeAXvMmE2pbvdxC0OT2p4qHC5XlW+jRgKAL
2rHoDXyqayyxqoksGB5new87LUaCBt60vf3HdQVTsx6VEHfvz8GhK8W+Yskg82+3
CffWF8Q3d7fX5ycmJ3EdO9/pFeqYjg8axoaIBgDdlC7paHs0nS0NqM0CZiusBXFp
xG3dwUdyN6GRXg5mhX1DaAPH3nKNphSwqrY56gSE9Fx3pfAwc/a5KPXpGI0zgiSg
90S/tfTWURzTV+AFVj2xHQTtXy06s4niFReqL/Goxn83wbcKZ+LlwA074iIpctUh
bgeGIfmG2XI6WlCTtVMZjW5TIVLBwqGgLfHOi6Ck5Cq/+n+jV034XuUskWE2DCQE
98WxhP+j7Ma6ipGek43hbXC+3SnpUYC3t330gsZR/ne7zaWf1v7Ip9di/8cYkUAE
Z0ou6gRbwn5qo3W5J1esPocWOodVfu7KoORKNX3Op6eVOuZXTvqjs/e2tFClis2s
mixFRVworItxiVd6mNcJz/F9B6vZKpe99KT/LSKtWa3dmQZC5FEgLTv2jB4XcbqV
FtCCOTZiNo2XuNykczsnA5InEneveq6EgPZfS5tklCfmYxOXeruEdV2uaycgccZu
NyL/3J2ZmbJBZ0iHUxmYtq+66w3HwA+z4b7qpRfkoamFw/ytXeYV+WCmnPYqxABm
+w71AIomzoDmQDySkZHquKbogbPZ/ceD2pYKhp1ATN3EJBbE9f0PnVMnsMzcXXpf
5rBqxLnBIeQPAEREZ1Gmi+vwgZhYGkEnxCb+F3th0Nnq/bFd/MGfeKaxRTU0SHvO
GpCZ5cRXo4bmS2Go6CsJHwdFkoD8fXr3u80pEHIDNL87SfDTQBjYtackf9Ak6Tkz
I/aXAfGVTK9aP7emPWKL8ZBg2DHUyeBl/mNb/j/7SEWheCglHhH/sB1BjgJhEpY0
vv/dJNrnZJ997xof9uR+kuG8sC1aOC1ile14VGeFl4s70D2ueDoHJF1c1vs2FBgi
n/EmrQqlpCzS9AclniMhtCPm4XIuRvp0w+D6iFOD/e4tnvpWwiKaVsKnphFHHvcQ
GGRx20/zoyOHpWGajs9PvnMxXnKLMRHzf+QZPMC6M6SgmL8yWzUD27zj6Yzg8QIp
w2yW1JwpRPcBJ6GCGp7W2CynRj8Iy1ez6hogFey5xUVN9JYoan0TbW0BSTef3+cQ
YBIlKD1gvpDTI+/zalOPLLOkF0GTlGAlv11Pns95nDQu2I0Zqvhcwi7oaQcJp6Fj
CJneK3nZc/zXxsQGtmx+ksMtUO+a8tJnqMbPS0Hb/m8MHJC8s6uSmaIqfM2DkLxR
q6N/4BVA9irvekXJFEUx/PJCjMb7+LKyiyK32ISZJcrftI4u1NvJ9XVjhwembmCS
r6h6CHX4q2jxEXImEpyxNOpgAmFzNEfXoi2McFukfLih2W/lcC/knLRgPEeplBVv
YDkNtOTkOJdBpCUPQwJpO/FJ7YGoDl9afJe+JsCKaueAmWiM5WZfxpBhU/4rQWkx
A5piJDOO8xPI9YG3h/zAc70DUWnnrAdduGfBih4ajPo6O3q9Mcpr4wN9FetssKJu
La6uJypPmANyFjhGTOcVyJ34OqNKyIIpoZmwJyLJec1tzkxgtk0eftpSjwr2M5Z1
U/UP/0oCzNjocfSQtAroIF5XbrHzFoJsVnap+rIVTfnkeTFfoWo3TbzG7lH43jx5
xgSzrZqhqUXzIlXCXInHVz+g+sYh/iEL1J40o1YqKOwgYy3iXeIYDh52KANi5q8f
jcYBUAMHvlYcvmU+03yES3KprBkCutDG8oAwSthdbQf/1CbZRsZVlRADFyp92xo5
3Ccr0TtVywAzwrI33fAa48/yPG2POOP0TxxParbhaW3y6CFKi3gP6xmGLh2Y8LC5
W5H2npZlKF80rcW/1ggKOjHB1RsqCuFO7WbbcQ7X99MZdSMGlok32QBlPD2/Ubj8
8EZQkl3zBdWqume09gpulsc6BTh5bum0hveenZZzEmo2+yvdcsaZSdX0o4+P9AWW
+2KcCuS3c0Yyrvy60UeCutRTq60BNODaAGP9KfhAkmgCNHvsdgnFFZsT94iCzsNQ
Zy1aX3Ep8hc6aPtQA2NlXu6aeHzVDCswRTvDjte5mwvwCLRlYoaQezfhO8XEQlJf
TVfzNxHzqpY+lYiIMpjvgvlxXtmW1F53clb/pABGPvtkz6eBQuqRpFb3qkbaRiZM
BHy7ELFcYl98sXNvIEfTlVhEmMo8EStuBakrmaXH+cadRWa0ynK+zstGPXF+Y3uk
8ZIc7BlGkOBN02ytLOrDecm5SC2NGd71DEB34oVso0FG2wBRpZuPBtmq17UaUihQ
+LwUHXSfQwD7cGYTrC7VQSdeY2NfLT9vkcpcoFOz7xm5qmmQkGGYrd4wRFGJI0yU
GBntQUd50Z4C13MWWU1NvBbqjMwSon6buH+cMub0xRrSJkipWNVfYgHNeN4qGnFn
WhPQGDwG4zoIc/dU3sxmLBnH0V/Pz+a6Qzg2BY5JB7rrj/wM03EX0V4OMTmPgNsk
etuV3OsYH6bB3aNxAeZCgA02vbQH9Kr4+Q5xU0a2z5wy2FkPAj+MtI+CtWnKOf2K
vUH+glExu+hYxONP0fk3HCFpS1+O1Uvr8q7hO2nypymeV2gZzCvvXL0GN8feMrDB
revDvAMTvXzGXzTWsX+iUniRCoXnyh7LptVUmiXXY6b+ZrQ5VVmARtxiE45JdcZD
JC3VpdWvHrkAkh3lp38+BD13rezdBz1T1wY2UbjODbLNEjxjcP+RxgD2LdLVFazu
xmD1Ymf4m6wSj7i6kaf3uzk40IXJaXgpzo0/wfR+FDNtTjR6mfw8h8vP5wX66fMk
EP8buNOywDaWlizkrjE11Ec6fRHk3rwKNqrRKBaj1i0z2Uqj0AcqWlPh72mhKuBZ
qAOLUwA+qL+2c/BlifVyhOev3Qx7nZiyh37l0CjE7sFCToePkhggv27foEQ6UJUp
zdXaKw8FA/GKjwsNPGMaWSbadM0a1vAV7c/+hWKuHy++7fXuelCc4C6dl7sw9wnP
EswSSl17SX0h44RPNn/CZJJETEKPqSNZHlfulWvuvLOafu7t4Pty5yqe7cvDBBmg
PqrMaZ/Vn5v1ZZKEHc781APWbzgRzf13kwE+re6dLx57saabJSKjpIH87+LCX2Xj
uHTWzoEmCv0onCeRJRlHdgMdWaAYuHAW0uAY9Hc/7v4F5Y6oUZKIQ/SE/v+Fgdzr
VYK1+y26H+BnQFA0MOEWhmuEc4qAcIRq5Vk17LB7UBP9fQ5WdncA3TGwJy8ae61J
XQ0uCiXny/cxZXeoZktIET561mjX55yxma7KcSXP2VJHT7PZcE8G98oxz75Nd9L6
/W6ggmgkZs4XBnr7E5D0Wk32xhB+6DEYk+/c1gqTNzpk6JVoadjlkUtoSEHjdQYU
Evu/H1F5v+Bowsg5jolXTf8mZYcD2OyXx2p8q2iMuu6frKm2oOTKrNz/DrxfQw3A
SN5eXiyRh7JKCcCxntzT7QbNZjmMe6NGAyzujvtdl98W0sbvpDaSjKQ3gIzN3KQd
VxRV/9mIgIYklfikw0EwPIB/x9ax4SdWva/TucYp5rVe7xXjAjyj+0iLEz1Xdrhf
FFFvoy1BZufuMR7+G1JIXK0MToK3ArhaIOoBjItcm3UFZjWpwzRdTOhSTuGt867y
PfyNZb+uqYGi3y5pFqbIAs7Q4Ez6f9Utu89v1BdyszYShaIO0VXcOAHco9Ljpq/7
NcQF4tksJC57NKNAlVq2QCAY3XEEBp8rOK6G9JxXgnoY/eSzY91jBtiVbEKXbiHR
TEzr+IyXXAyEYBqPWu/Yv3HjX9X41CyIXfZLuDvUQSghhldmGu1An0zf5of8JNgX
4Y4Psglgt/6ptlIkQwVu9r+UNsA1WsmZ+oZ7jc5MivrERhep8NaVAdbf5wOvxPQi
wLb4L6dVktgDw+lsaa1AtJ+uWKWvePD2WzNoLqqBAd6yp/2fXYeQsz13Y1xGKw1Y
jsia0J0MKLlO3r0B1iWuJx2+67ISIz0OVNf7XBwHfh1xXWzzzLMz5QZXV6Dkf3Ld
4GQgZ8fZQm0AmaQhjxcP77n/I+ZxhvWCf9L224oXoCfMi5vWUJep1rRhdY0dv3bn
r70VRAUQjDU6wpFssD1XAF+3VpFPUZhBPentHLsBFMAJXLrnOsr8hmfZKi+Ttw6f
ZnigYhBiTl6MtWvLNML0/Z1Y17fzjCa5BKsn0o5+vi9s/yJVKWl3YIvkFbf1DVu6
PhBNGF4bJoT3uXRs2Xnm2cv451cGu5axO95XsoQ3b+x+TJ1fxYKO3fD4IMsjaNtT
5LYdxqf+t21dlwEg6Rd+BCY3tT9pBBhHZOPUB9LFmhhITs/AHfY6Uj6SKhp0SzPs
O3GbLwxTpNWoghrA8FCMAXJGHs/Ri/u+2vNul9TPeoWbPcsDF/YWQ0m8dXr2mi7n
V32AJl138FptSEodYPlWIlcpaUj04eeC94c5grMfdNHSNQlK+Z6LusYEWPrlpdKR
jyGql1Vym9pxlHGLBsTu3KuKi+xBo23HlluEbhjyv0VTk4a9nWsEilZ0PzH2BFVS
v4yxTkFPCrMATSg8uQJlg8sBQ/02U4fsgwr/76Z29J+MYqI2qJOwYmzc4s1Fj+nx
tnxUbtmkrN8vAtQar4c9hH23+kHgDrzrc/2thIbPjs0H78MuMc47p/z8uxWPcU9p
aG0zXFYckSttKtJ08FJG1CeF4DZwxQuYTH0glnBFhpptJ3X/WUYeCTTIxW6OP4Xj
Ucp4TDIzxKHZnHqNoscLQ5YU/Z/7xsowEpxW0CBbKwEBDRQ8c6Ug7d4Bc8Q/IlL4
08J25BXkoPW5Dv6lztLP/62QcKIyupvGMUS7/PokErDVnTVzzjjg28if4z4BKWO4
EKMbveWJhnbvskUfV1g+zScSFVR7gwnxBGdyzmnMeIS0snDPlbIS9Vx1G82CO4IR
G5A+lCdeVCIQVVm+UkTFwymjeXaEK7vpJdJsJwaK/45kDGrCbBXbS5FlPE1qSeVE
IfNWslww8MxY/2GuR4WBYN/XG9fB4KcVJgVs+qPNSLPqrtBqq54niN8JqOj5O9yN
0ElG7hBEjvFp93sJIBya8MvRu/UC2WyNMwIk44oLJpZW1wSbel5qooekXFpEYXEr
9v7e1qa2iLHojVNtRVdbcT5YxUFxlbNU3+xTFt40qr1Q+p+yAm+OSD2zF5RtxcWW
Y1h1ygB5yY++QrTQdyqhgVrJ1Kdw1oESmfPMh8Re2BcomGc4MZexKbF2XLy0+uI3
kMJAYW97yZCsGcvpxyKdguELoJfkDBcN7Ly2laByVHniIshV91QC8oci7P0I/Q+w
8+Q2AvemNM8wrF8dNuJFKwGnqPRQdN33nNTP1MkDtaBACpIp2I2Z9YitVHXKpeYW
i9WicAN9XUF+o58l3SFClJn1ej/H6NhFO4c2lkAVzKJNCkzHfOl1EB+97xS2aT7W
ZxQBaaTmb8sBFZ7g6bXSK6PQ/ajeuEb6r4HekrPAWzgpYV3j5tTnaCDeQxFZIZxt
xQlUrxP+czOHR8CLHwuE4Wk5vrSCWsUX6Vqx296XfAylQe+VqOKfSKYpTR8a6vdN
Nm2VR4V1Jn3xhwXc5hUsC29QJtLs5j0p0MUZzgUFWnyodx//lKVYHY/8fvl8hnIN
dZkqxCrtqBdyKJzTyTuYgAHuWdBI402675GcLYYtJviRey2h5uAPWKOtqecVEZ7z
cbhNKDe5pPRkor6JEIufMvfPV0R1g6MiU4kCHcEdieDvUkUsquK/aBhvVjy/rVuS
HRf0tK70c9i/4nWvc8u9qUtn+ui0mYr8Bm51yNEy59u2MVPeqWGXXheSE+a4N5/P
6yuGCofWaE3OmklpmZ76vn+8CJF4wrUi+1gC02LRK0TEustu4tfBENs3cJ8YHsKi
KqnY1+/aISZItBrbZT3YxCTt0TrD9kdugP0ECHwPZswlaMXNxfSljfxogYEBjunv
JT/lHhEaiRN/+bUxELt9hZvUTEVhiS8PtGbmxQTOksm3oc2vDTLyI/2iwU8Q2dP5
J2Ms8pmS2pFH0o6ZHaAOTIZn1/eL7Pm62uBDboiDD0OCQ1Wao73ca+CCYYvhQiad
Jzs93iOZrPczC+MF051dumcxICuHXJdPxYQRxZXPHfX+pWd0aWNVrxLKTugLs0+M
HVvmDKRjf2NqMPxiYj9ZzRxtHMi0e1mKOHWtLBitU15jwj+wxSHUSrgepFd6+fwe
4hAXONULqMWE+Wc5+XrDZwHBV+vwN1J7gF5+zKaniTAMuhRjGOSHtKBCgdV/v7k7
KOHM/k5S7bc1gcWvn0Wr+lQLYus2zpQKKTcOMv7IS6zU13sqT3V5jgCYm7jO/jaG
P86tJXRdjUtOs2Eyzc9oH4/t+UXTBkgitkn9xdsT3LuCqLglLeRnnCECw1mHp3ZN
Sur+B44T6jGqjl6z87tYkmf2p6cqZ0O7qSCvQjQq6MBSOfs6UAc5Ydn/faBJOl7Q
Qi90lJ/iUFUqhyTlQidaDsRlwRZdFVstwDXz7XshTNCFkk8SepOjnhrJHd7woBho
QwIvTcq9iXb14WEjsOiSnigL0GXtzKw37wVlMCACZTzBxpJcwFk2d66BbaLYFrme
ws/SBcbNG/7qmR+NanqHkvVh5x5GY0DiRmAm6AtgxD/L25Ec02/HwgBoUmO3oNEB
xEdbEnPW1LRfEeaO2UU2VkArbGfnE1ChnG7diKIwgzG/1S/J+7SYCxLnzvx9WuEg
TI+qtU3ZYQh9F4rNoz12N2uocaPDLWM5rCfeOAUxzskcT5eY9EmpxSJrPTSemoaP
dvFxdECpPMy4k6hgJLar0QO/FiFcUS5SRbLMa1z6hltUu9NfeBQkI3ny3MIj1Ejz
S4yvYQzUfSuJGyxIM8h7+qew5GlbPtxDX+otxAxChCtIeTJN7MCTUT64fETB9yXC
1U+aR2SGYq8Nvlt/jPU/Kx9T83P9ziiHwIC8QR3vQQ6iiDyFI45gIsNSg7NKwkY9
vMUnPGkeFB1A5gyomx3TG/vje5QqOn/dCk+v9DZu+fuDCDDqS65wu3twcP2+eY8Q
Xuuxmat2IWcuTqMiOIIE2o1jEMlyT0K90c0VibviRSmGfCOko0yQ4vKEimwUTriW
TGCxvs+houTExBq1FNCL+ELOpiUyV70YJnAu3LTQspBxkf76FXpasdX/wquWgTMw
rjs1zVC771WzEznPxcarGmUvmmjzJ9XdaHMoRcabtmcx2APaSAD+2PJLabuUO2x/
wPmNwjtA/kJyPHWdoi1wDFZbkmcUJC0gs2bSJxV2ifQo7B0HioV1y14Irw8PN9KW
Hr7U0vMqCSczwE2mz5yDzeNOBPDy1PDyjMdQDjjajh88lGDY38LdTHb3n7SDu00d
7cBR6V2e/UMg9ZIPOvH3lkf8woaXJdcxx2lqzJi8kAfo6XY0ArB7DCVQDmRKEP5W
ANNx5Wtj6BS1PbuHfkio4SgpFTboHmVNiXuljdTB2qJ3oqAz06OmgiRuEQy2k8wu
RR/562n849M3JZ5j3PaCCK4kHsIkw0kxei22u+lgA5FBQADAP2YNG6ZqC4RhLsAd
W4r9y3UaqFxpt1sgXg5HMlW5ccPzfzzrTU042nY0jJ9k62UpP1gBQRQbyyqY6UAF
RjpbiReQLyo6UGPFuopDUJBtKIRIFWGNrPYrV+deZ6hfjtQlHNY+0HKTR+twdF0T
TXdaqEIvOSWQoVVG0MssL/vjcasJc+FMXUKWZc4UGKPBmoGHWcodRlx3a1YLHUdf
V7OK2NJriqcky1EzEjCwDgg8V3E8ubIKI3LU+fXIdcoXBmSlfqstqbOjUjhlYCqC
18wjUQXjd6J34odoueE1sd4X7UqnX/AOoFGP4k4u8+8thVl5bGwgSvWY4cUVi7EQ
cMHufIdAueo+lVQ0zn9y/aprXbGKd0w2eQ8T6CQouxJPwEkMANu6nxnFmLkZ84aJ
UWhIWkI2trNnyKVwHz2NiInJuVEFiLM4xABs4/P9AiXcoQSmBjVb+E4pWBksIaN/
kevNTRy7fsE+YWLY/X31Kg6JXkHRTm51YAi1bmloHSY86f+x0QuqOIFdjA8ctiYJ
eILtfwth88K0rdn8GQSWR872rkDT0d4FgmMUFSvnSRe+B4TwsNZU/O9lwQlAGoS7
GIlStPmsOu0zWRl9vn7u33rdxTOvyacQjUtDoJQ/sVWOY5hyaFHb41QEBgJFFb6G
umWR3xT95eISs55GoX9J6YY7mONYOFzQ+ZYZtha1Ij8jWwSRFedVFIs1xOkS/7lR
aNkxQlSJGOa+pIpJiyHw2D6jstV+uIcOISRwcDnM3FpiWxYTHWbgnjFvJu7c1DNb
Mhp5p5VBUE5ATzFpHVN0yBHNCqZzEsVYjv5pou779Q69TYb0H92HTQWe0VQwalod
U6e6sD0yUEGNT5FDPQPosItzAdBx6+a+czZaTtB4vZYAdYJy+S4XsLikNVrv5tZn
keG5kN/s6pRL/nA+oKP7BRJzaQulGy1Jiblvtcr3qXCMS+vg+Ya5IH4BV9DlaxwY
gPQeGJcQS/AbAzEX116coCeisHvYoTt3Atd3LYjHpeXV1eKBiUtRUBw3ppVuYxPA
0/Xs0krvsCKLLJuWw6Ee7IoqAf2mpOl5/dQh+tDWMbVEqp4cBk+DJM3YDBdEzzil
VSR7xiq1S0rUTIeoRcMpDhdfkbh2bVzLDNylM97FkCl8Yzwpgob2fdTB4V9NNif0
rZYWogdJTHl+tTNRws37ZaAH+fqUdFdkR5MS3eXwp2xmWFKJXtEolG8vfuNFEX1a
5xWR4nhFfPQ6EN4YBF7w/zCNnfzYF/R2yWi6GeZ+pTLmlHQKNMzuCMxtKnol3VPf
40xy4XjPQQThDyNlAxJPnVH6zkJWuCl2R58cz/0sdazhN0FGAi3zDBlU5dx7usL6
K0Ym58SXHU4KxeIci/fdqAXVln39SV0eXx2nyC/94UYDQfu9VJv6CzuEjZYkL7QR
t9pDs8pPJikfsaeGwSrzY/746CdsuagikIHh0xaeaTbD8WDx9CRLBS5LjPwNyoXb
OG/DRpUlQZpiL1jsdjCtPzwA3co+JQ5Ru+JWxUPE17Si+SK5Q3wIAyNk2I2LwkyO
8x5GQsfW5IY7+E0AiVBCX4/UBasSXKM+eFJS843Z8zhVi7Y3NYwXrj3ipxM248EN
qm52sDKxmxxfiGwGogPuYvOKdXLVZLvIl21cvAamfi2NzQ2vL7ghF1CacQuxSmt+
ENzrsH9V527vv0ilfcyYbomGwqkyT292Qj4LSFTb0wAFyf5/v7hpBH+nVTKnKMk1
JeCCQjz7eMhfeuyszY/QCaS+auvVOm9rmnteEXp/GYaiqpr5admPbRFVK6E2S0D8
J059D81AaFyZzPN6XRgOQBG48A3kD3nwKqi3zZtZ0w4lNSqBNo+IrG/azUc9swC3
KAMX6Y1BIqyjpGZ+wIFrWiusao5xKvXW/o4a4V6GyvvInsbDeNLhT7aLIGrax1JW
jSmWkizJvMb3xwa796RPEe2i4Owmtv6wHXIAdBJvPDIuisLQ9PqceB6CLUwStmLp
Dqh2RL7Mhflt2aIK2H96dRLUJl9xoqUgPxvxcrLj9g/+R1J9unf9WsNYDXwjQOIU
NwSIznWGn/jUFvU8Q+BRCuTUQ/BXIAH0pjJDi0SwMJg0xFwqPJ3wXhxm9rZIIIuD
K9ISi29AxIsb7fibF771dm7IaF4SgJ8YvN2fCCo0LOTN/gxzcem+3hWZ0balouSN
nsWYiz5zqaa+k/y9LzzxukRfHk+LwFuaVRs/Slr1LuzSh8J5zHL+gQMkElGldi7I
lr/tQiW9WEymI46ngyDpKlRzAiCkz4e7DYVTeQ3FGYtfedyT/P/W/5sAyzigt+gf
sAw85Ne13oKieshVmGo7VuwgcruqD7crtFOwMxTTkNnBbyJxz87bA9haThQlPPgZ
KWELPxjydAFj41ppKj8uhQdiJySzMGND+5b4434Nb+H2yzjh2uwSwEvMEHTcImgS
4zohN6ZePUAzzNuKRPuX78QUxft4PObwKcgORmtUk4Vsg7Dg6nA2ZR7MFd+DXFsT
Q/x3qJQuFMkBCw45+OhRMWlEPPcJsgSDB/j6HCKJiPZIJvpvsphRLHNGisOhoZut
iQyLcyfI2UTH6HTKE+QOLEb3L5Pk/jgVppA/5DKJDYRwWmqgX66BtUVMDFJtR+zg
izE29dXfs2m3jr5uhtg3lwgR1rCAr73WdiKX+XoXpGm2cIOj3TULRikO8jb93p8u
z8HPVldqUlDsOhU/6fNXonpNisoh2lrV0ROGSUm6bIxEBbiso7uaOyy7xnDXf6pg
/THYBDEuS+vSI/KhvgkoqzuQQC6yWkSgC8N3Y4IckTYnjmRiSUPU3Mc5iDTQm9J+
Vv96YRCXmZm/LBr3U7k2IEtx7XM/FaE7nPwu/I/sb2r+2aQXMKl6bPa/9gMN6kVk
pu4yWw5HiJXPI/C9I1g2c7VQa3ytJdg4KVPaSEngLT/RDOqYHRsTEKSpc3nZLcSo
27tQd89Kcgwa21bRdlMqfO21PqfRjKeHcd+t+ASJ4CAGK2iU84DX+66O23MmMn3A
HiduONWK2fuy0ZIxdM1tBQROCzYLv++ysjAxz4KcseukRb4zWnhDmLLsfWpICf0G
rXHELZunpCnLZ2lwWCVHeVssuf6tulmWqCxjfTrw10QaOEwwJ2dD50UZq0A++Zu0
MnTpPlwIr/BwTpPHjxokrJhetH4/P5quyNGA/91Bf4nGRdRoUW8Bhw9IQPSdOoXz
crRERAIhOeMBeXvUUd/yqAjFaiiZO5x8g7YjempWaBbN3tkd3YweDUhuXyzUPMQB
2DML2ofH4G+tlWDTqTpwuI9FQGDtuNRTNy98fwuo6f9lDVk9p8ju3vF5w+ECXoNo
3E7M3wyYhDhli8rK4boDRCM40YOFyCxSIaczLRxdb2KgW9D9wnP5Kw9/yCRWj9Kd
14MGSCGURyT5cWxK108EH43J2DNZnamGFhsLeNKgcXjKgzNePnt4MiHt9VlUxwrv
YNK/fU3D1o3H1A5D+8is60LwrqwyPK9SPNgSNKzad6FKOUXkAbnyOQfeKQFCkMY7
Tf7w8hugFKOHp+gt0M1iOLc3PgYRqDrUsqXmJVzQux4qRwiAKlb6lA6IIF3teAWy
7mEhb3py7iF3KSvv5dmGez9+c3p+IB9wDbBKjDNWf9WTRkgsBe6l/ONP6qAyx/kR
bNnyeFNK4rDYvMxM0ainueER0jP1TBsispQDdzy4YxroExerIifI/74Zd+y4DCoa
oZjmkWiBFFZa6chrLKbaS9SChxbCzgwxr2DuOeAGJSGlS6V4syGRe6NXlR9R5cS6
1r3cmCvr0snY2f7j9ODc6SSQ5g+dMQQI3qetMhvU8xM6y9k+Glv1zdT5gZl1CDuX
cP7rRFQd+yXMK2b9ItboWHCrhNo/VJxPrJ+uVKWfMAxQpUURlq+PGzIA2g9z3q+F
SfA1i80Dfa6Tz2Ynuct2HKpyOSVTCM3MIWXYcbQtHGK/Ne4w0rEGosEBLmb16mUS
uwzrZOb4Wpkbjo5/uDVP3mDdEV/Wip/1Nd4fLrTVf8MjNGNntENHpPqDxz9iLRMF
ixcrpgiMRjDRW6fy6YYck4hqWUKaRVgY7xRvmtyZDFdD+RNYIlUCqQpHW3RpC3L0
rMWcfbuGNx8VJN7tf0KJmOJugPIRibiDy0yoGmPnijU7eqV/As6+NKo2y1CJVX1O
BDksRrovxwswJECZjgdHpu5m6BT/VlQlmCXzvJPjTK+aVI69nd0mzgL5zEuCr14L
EaQSiuNxRvozor8UvxMqezLNYt7e+Qlp0IP5n2i4wUTY6IXRbUjnRvznt4lB4BYq
U9PJtet8uONVShgqn42MpLs7AzyhRrX0BrErItjQzeTvfdmQteGtcaanIzq4y8Ng
FljZtZenO2gUO7asSRI4aTz+LoCTYR9mvMuPnWBuEUqYKV4PJS0hQSbwrXZouOKb
dpMCZyfoWSuN9jDhTyI2APaMEBRo+2HEXeO96ID6KWWO0RxmjiXU+TQS0UloWXcU
zMtcOOykPw+TUMC/WqgpJE0r5iT7L0MVcS0D2wBa+NZumxdq3gCFrq3pZm0Wq9xY
ppxskSA5rKWDnAcrJj0rZJCJO/2f6uE11FuCHmXlvHvOT9eo0g2Twny5aClw4aL/
LcSmV19w12twWTZDlV8KLfMp60JZTdMaxPdaIkk6BlfnV2fAoCy7NciAMQr0fjuX
XLguPTRZdaa7vCvVBNRVN/WMLLwkx5at1Cwl5ZDalruGcuPAfEwrOYDL9yfIJ7og
GZuV+ovmzECC9+Tb55H0EJDEGzUNhQYocz7nuYAWa8JPD4sT0ocGDBlFUgQSKg/r
FOVKbcWHxVWwgYhke3eVxjlDei/ckaxaPg9hygUaS8bKm9Ghvyl01FDDFnz1bIjH
MzSbc3ATsPR5iWxrUF5ZzWH994ORxzhWJwegO4rabn5yhv1qH4NLDh4/7b93pb/W
5Zl93WWebAL3mnN1QtY9jLFAux8Twr5zZeHIX3b6C7vsDxyOjShcH3PQu7f4kvJ8
WUKVMfr6otd+jVrJmGwJqJ2nzSjo3C8xI+wSaYa4hkGSXU83o90BzR8BtqaiqYCX
nD2gjIcLo9ojGxXcaUZ1DxQa0jVZcgfCTc5J3f8nB2Y8Iu7UeamFLyzD51olc6A5
92aNjeMer/XF9JWfinIJoRlRRV5SafubuI0bxHbfn7nfGxjhLAnXhy/+DhlPjOOt
x/Nc/eQd+Hcde93bA8fkXutfpQw04yTHgF+lL6JkFc4cBm6mLFRIxDiZALm6Zw3M
+V9moGxbuhVcaagKWck9+Ow/mlvip6Uxb2B7IGiJ/f+Ah1ohCVxIy3vErTUQXVZB
qJxNCvRXJACrpj+sTXH+1Q==
`pragma protect end_protected
